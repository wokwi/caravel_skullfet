magic
tech sky130A
timestamp 1641006614
<< locali >>
rect 44080 325330 44170 325340
rect 44080 325310 44090 325330
rect 44160 325310 44170 325330
rect 44080 325220 44170 325310
<< viali >>
rect 275750 337500 275780 337560
rect 276370 337280 276400 337320
rect 45110 326150 45140 326180
rect 45010 326030 45040 326060
rect 44090 325310 44160 325330
rect 242300 295600 242600 296200
rect 248400 295900 248700 296200
<< metal1 >>
rect 275270 338070 284400 338140
rect 284570 338070 284630 338140
rect 275270 338040 284630 338070
rect 275270 337580 275370 338040
rect 275270 337560 275790 337580
rect 275270 337500 275750 337560
rect 275780 337500 275790 337560
rect 275270 337480 275790 337500
rect 276360 337320 289100 337330
rect 276360 337280 276370 337320
rect 276400 337280 289100 337320
rect 276360 337230 289100 337280
rect 43290 326550 43510 326570
rect 43290 326460 43310 326550
rect 43470 326490 43510 326550
rect 43470 326460 45050 326490
rect 43290 326450 43510 326460
rect 45000 326060 45050 326460
rect 45100 326410 45150 326420
rect 45100 326340 45110 326410
rect 45140 326340 45150 326410
rect 45100 326180 45150 326340
rect 45100 326150 45110 326180
rect 45140 326150 45150 326180
rect 45100 326140 45150 326150
rect 45000 326030 45010 326060
rect 45040 326030 45050 326060
rect 45000 326020 45050 326030
rect 43700 325310 43710 325340
rect 43770 325330 44170 325340
rect 43770 325310 44090 325330
rect 44160 325310 44170 325330
rect 43700 325300 44170 325310
rect 248200 300400 249500 300500
rect 248200 300200 248300 300400
rect 248700 300200 249500 300400
rect 248200 300100 249500 300200
rect 249000 296300 249500 300100
rect 241400 296200 242700 296300
rect 241400 295600 241500 296200
rect 241900 295600 242300 296200
rect 242600 295600 242700 296200
rect 248300 296200 249500 296300
rect 248300 295900 248400 296200
rect 248700 295900 249500 296200
rect 248300 295800 249500 295900
rect 241400 295500 242700 295600
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< via1 >>
rect 284400 338070 284570 338140
rect 275520 337910 275590 337940
rect 275510 336500 275580 336530
rect 43310 326460 43470 326550
rect 45110 326340 45140 326410
rect 43710 325310 43770 325340
rect 45330 325120 45360 325180
rect 43910 325060 43940 325110
rect 249300 302500 250300 302700
rect 248300 300200 248700 300400
rect 241500 295600 241900 296200
rect 249200 288500 249800 288700
<< metal2 >>
rect 9350 351530 9750 351610
rect 207600 351600 208400 351700
rect 9350 351280 9450 351530
rect 9680 351280 9750 351530
rect 9350 329210 9750 351280
rect 35450 351550 35810 351600
rect 35450 351190 35490 351550
rect 35760 351190 35810 351550
rect 35450 335700 35810 351190
rect 61480 351460 61700 351500
rect 61480 351190 61500 351460
rect 61660 351190 61700 351460
rect 35430 335660 37330 335700
rect 35430 335530 43780 335660
rect 35430 335510 37330 335530
rect 9310 326570 9760 329210
rect 43680 329020 43780 335530
rect 9310 326550 43510 326570
rect 9310 326460 43310 326550
rect 43470 326460 43510 326550
rect 9310 326450 43510 326460
rect 43700 325340 43770 329020
rect 61480 326420 61700 351190
rect 45100 326410 61700 326420
rect 45100 326340 45110 326410
rect 45140 326340 61700 326410
rect 45100 326320 61700 326340
rect 207600 351300 207700 351600
rect 208300 351300 208400 351600
rect 43700 325310 43710 325340
rect 43700 325300 43770 325310
rect 45320 325180 45510 325190
rect 45320 325120 45330 325180
rect 45360 325120 45510 325180
rect 43600 325110 43950 325120
rect 43600 325060 43620 325110
rect 43730 325060 43910 325110
rect 43940 325060 43950 325110
rect 43600 325050 43950 325060
rect 45320 324240 45510 325120
rect 45320 324140 45360 324240
rect 45490 324140 45510 324240
rect 45320 323870 45510 324140
rect 207600 296300 208400 351300
rect 233500 351400 234200 351500
rect 233500 351200 233600 351400
rect 234100 351200 234200 351400
rect 233500 314400 234200 351200
rect 284360 349440 284630 349490
rect 284360 349220 284420 349440
rect 284560 349220 284630 349440
rect 284360 338140 284630 349220
rect 284360 338070 284400 338140
rect 284570 338070 284630 338140
rect 284360 338040 284630 338070
rect 288710 340370 289070 340420
rect 288710 340130 288760 340370
rect 289030 340130 289070 340370
rect 275500 338000 275600 338010
rect 275500 337950 275520 338000
rect 275580 337950 275600 338000
rect 275500 337940 275600 337950
rect 275500 337910 275520 337940
rect 275590 337910 275600 337940
rect 275500 337900 275600 337910
rect 288710 337220 289070 340130
rect 275500 336530 275590 336540
rect 275500 336500 275510 336530
rect 275580 336500 275590 336530
rect 275500 336490 275590 336500
rect 275500 336450 275520 336490
rect 275570 336450 275590 336490
rect 275500 336400 275590 336450
rect 248200 314400 248800 314500
rect 233500 313800 248800 314400
rect 248200 300400 248800 313800
rect 249200 303200 250400 303300
rect 249200 302900 249300 303200
rect 250300 302900 250400 303200
rect 249200 302700 250400 302900
rect 249200 302500 249300 302700
rect 250300 302500 250400 302700
rect 249200 302400 250400 302500
rect 248200 300200 248300 300400
rect 248700 300200 248800 300400
rect 248200 300100 248800 300200
rect 207600 296200 242000 296300
rect 207600 295600 241500 296200
rect 241900 295600 242000 296200
rect 207600 295500 242000 295600
rect 249000 288700 250000 288800
rect 249000 288500 249200 288700
rect 249800 288500 250000 288700
rect 249000 277000 250000 288500
rect 278000 277000 281000 278000
rect 249000 276000 279000 277000
rect 280000 276000 281000 277000
rect 278000 275003 281000 276000
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< via2 >>
rect 9450 351280 9680 351530
rect 35490 351190 35760 351550
rect 61500 351190 61660 351460
rect 207700 351300 208300 351600
rect 43620 325060 43730 325110
rect 45360 324140 45490 324240
rect 233600 351200 234100 351400
rect 284420 349220 284560 349440
rect 288760 340130 289030 340370
rect 275520 337950 275580 338000
rect 275520 336450 275570 336490
rect 249300 302900 250300 303200
rect 279000 276000 280000 277000
<< metal3 >>
rect 8097 351530 10597 352400
rect 8097 351280 9450 351530
rect 9680 351280 10597 351530
rect 8097 351150 10597 351280
rect 34097 351550 36597 352400
rect 34097 351190 35490 351550
rect 35760 351190 36597 351550
rect 34097 351150 36597 351190
rect 60097 351460 62597 352400
rect 60097 351190 61500 351460
rect 61660 351190 62597 351460
rect 60097 351150 62597 351190
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351600 209197 352400
rect 206697 351300 207700 351600
rect 208300 351300 209197 351600
rect 206697 351150 209197 351300
rect 232697 351400 235197 352400
rect 232697 351200 233600 351400
rect 234100 351200 235197 351400
rect 232697 351150 235197 351200
rect 255297 351500 257697 352400
rect 260297 351500 262697 352400
rect 255297 351170 257700 351500
rect 260297 351170 262700 351500
rect 255300 350407 257700 351170
rect 255275 349200 257700 350407
rect 260300 349200 262700 351170
rect 283297 351150 285797 352400
rect 255275 348040 262700 349200
rect 284300 349440 284700 351150
rect 284300 349220 284420 349440
rect 284560 349220 284700 349440
rect 284300 348800 284700 349220
rect 274710 348040 275610 348050
rect 255275 347500 275610 348040
rect -400 340121 850 342621
rect 43480 331950 43760 331960
rect 255275 331950 256842 347500
rect 260660 347490 275610 347500
rect 275460 338000 275610 347490
rect 291150 340400 292400 341492
rect 288600 340370 292400 340400
rect 288600 340130 288760 340370
rect 289030 340130 292400 340370
rect 288600 340100 292400 340130
rect 291150 338992 292400 340100
rect 275460 337950 275520 338000
rect 275580 337950 275610 338000
rect 275460 337930 275610 337950
rect 275300 336490 275900 336500
rect 275300 336450 275520 336490
rect 275570 336450 275900 336490
rect 43480 330700 256860 331950
rect 43480 330340 43760 330700
rect 43490 325110 43750 330340
rect 43490 325060 43620 325110
rect 43730 325060 43750 325110
rect 43490 325050 43750 325060
rect -400 321921 830 324321
rect 45300 324240 45970 324260
rect 45300 324140 45360 324240
rect 45490 324140 45970 324240
rect -400 316921 830 319321
rect 45300 284100 45970 324140
rect 255275 307400 256842 330700
rect 255300 307300 256842 307400
rect 249200 305900 256842 307300
rect 249200 303200 250400 305900
rect 249200 302900 249300 303200
rect 250300 302900 250400 303200
rect 249200 302600 250400 302900
rect 45260 284050 66400 284100
rect 275300 284050 275900 336450
rect 291170 319892 292400 322292
rect 291170 314892 292400 317292
rect 291760 294736 292400 294792
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 291760 292372 292400 292428
rect 291760 291781 292400 291837
rect 45260 282800 276000 284050
rect 45260 282780 66400 282800
rect -400 279721 830 282121
rect 275300 277800 275900 282800
rect 275300 277700 290300 277800
rect 275300 277681 291800 277700
rect -400 274721 830 277121
rect 275300 277000 292400 277681
rect 275300 276000 279000 277000
rect 280000 276000 292400 277000
rect 275300 275300 292400 276000
rect 275300 275200 290300 275300
rect 291170 275281 292400 275300
rect 287300 272700 288370 275200
rect 287300 272681 291800 272700
rect 287300 270300 292400 272681
rect 287300 270290 288370 270300
rect 291170 270281 292400 270300
rect -400 255765 240 255821
rect 111182 255271 192182 260671
rect -400 255174 240 255230
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect -400 234154 240 234210
rect -400 233563 240 233619
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect -400 212543 240 212599
rect -400 211952 240 212008
rect -400 211361 240 211417
rect -400 210770 240 210826
rect -400 210179 240 210235
rect -400 209588 240 209644
rect -400 190932 240 190988
rect -400 190341 240 190397
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect -400 169321 240 169377
rect -400 168730 240 168786
rect -400 168139 240 168195
rect -400 167548 240 167604
rect -400 166957 240 167013
rect -400 166366 240 166422
rect -400 147710 240 147766
rect -400 147119 240 147175
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect -400 126199 240 126255
rect -400 125608 240 125664
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect 111182 120271 116582 255271
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
rect 186782 120271 192182 255271
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect 291760 227814 292400 227870
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 291760 202648 292400 202704
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 291760 179437 292400 179493
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect 291760 137570 292400 137626
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect 111182 114871 192182 120271
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect -400 107444 830 109844
rect -400 102444 830 104844
rect 291170 95715 292400 98115
rect 291170 90715 292400 93115
rect -400 86444 830 88844
rect -400 81444 830 83844
rect 291170 73415 292400 75815
rect 291170 68415 292400 70815
rect -400 62388 240 62444
rect -400 61797 240 61853
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect -400 40777 240 40833
rect -400 40186 240 40242
rect -400 39595 240 39651
rect -400 39004 240 39060
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect -400 19166 240 19222
rect -400 18575 240 18631
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect -400 8455 240 8511
rect 291760 8455 292400 8511
rect -400 7864 240 7920
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< metal4 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
rect 86280 48800 86440 48960
rect 86440 47680 86600 47840
rect 86440 47840 86600 48000
rect 86440 48000 86600 48160
rect 86440 48160 86600 48320
rect 86440 48320 86600 48480
rect 86440 48480 86600 48640
rect 86440 48640 86600 48800
rect 86440 48800 86600 48960
rect 86440 48960 86600 49120
rect 86440 49120 86600 49280
rect 86440 49280 86600 49440
rect 86440 49440 86600 49600
rect 86440 49600 86600 49760
rect 86600 47200 86760 47360
rect 86600 47360 86760 47520
rect 86600 47520 86760 47680
rect 86600 47680 86760 47840
rect 86600 47840 86760 48000
rect 86600 48000 86760 48160
rect 86600 48160 86760 48320
rect 86600 48320 86760 48480
rect 86600 48480 86760 48640
rect 86600 48640 86760 48800
rect 86600 48800 86760 48960
rect 86600 48960 86760 49120
rect 86600 49120 86760 49280
rect 86600 49280 86760 49440
rect 86600 49440 86760 49600
rect 86600 49600 86760 49760
rect 86600 49760 86760 49920
rect 86600 49920 86760 50080
rect 86600 50080 86760 50240
rect 86760 46880 86920 47040
rect 86760 47040 86920 47200
rect 86760 47200 86920 47360
rect 86760 47360 86920 47520
rect 86760 47520 86920 47680
rect 86760 47680 86920 47840
rect 86760 47840 86920 48000
rect 86760 48000 86920 48160
rect 86760 48160 86920 48320
rect 86760 48320 86920 48480
rect 86760 48480 86920 48640
rect 86760 48640 86920 48800
rect 86760 48800 86920 48960
rect 86760 48960 86920 49120
rect 86760 49120 86920 49280
rect 86760 49280 86920 49440
rect 86760 49440 86920 49600
rect 86760 49600 86920 49760
rect 86760 49760 86920 49920
rect 86760 49920 86920 50080
rect 86760 50080 86920 50240
rect 86760 50240 86920 50400
rect 86760 50400 86920 50560
rect 86920 46560 87080 46720
rect 86920 46720 87080 46880
rect 86920 46880 87080 47040
rect 86920 47040 87080 47200
rect 86920 47200 87080 47360
rect 86920 47360 87080 47520
rect 86920 47520 87080 47680
rect 86920 47680 87080 47840
rect 86920 47840 87080 48000
rect 86920 48000 87080 48160
rect 86920 48160 87080 48320
rect 86920 48320 87080 48480
rect 86920 48480 87080 48640
rect 86920 48640 87080 48800
rect 86920 48800 87080 48960
rect 86920 48960 87080 49120
rect 86920 49120 87080 49280
rect 86920 49280 87080 49440
rect 86920 49440 87080 49600
rect 86920 49600 87080 49760
rect 86920 49760 87080 49920
rect 86920 49920 87080 50080
rect 86920 50080 87080 50240
rect 86920 50240 87080 50400
rect 86920 50400 87080 50560
rect 86920 50560 87080 50720
rect 87080 46400 87240 46560
rect 87080 46560 87240 46720
rect 87080 46720 87240 46880
rect 87080 46880 87240 47040
rect 87080 47040 87240 47200
rect 87080 47200 87240 47360
rect 87080 47360 87240 47520
rect 87080 47520 87240 47680
rect 87080 47680 87240 47840
rect 87080 47840 87240 48000
rect 87080 48000 87240 48160
rect 87080 48160 87240 48320
rect 87080 48320 87240 48480
rect 87080 48480 87240 48640
rect 87080 48640 87240 48800
rect 87080 48800 87240 48960
rect 87080 48960 87240 49120
rect 87080 49120 87240 49280
rect 87080 49280 87240 49440
rect 87080 49440 87240 49600
rect 87080 49600 87240 49760
rect 87080 49760 87240 49920
rect 87080 49920 87240 50080
rect 87080 50080 87240 50240
rect 87080 50240 87240 50400
rect 87080 50400 87240 50560
rect 87080 50560 87240 50720
rect 87080 50720 87240 50880
rect 87080 50880 87240 51040
rect 87240 46240 87400 46400
rect 87240 46400 87400 46560
rect 87240 46560 87400 46720
rect 87240 46720 87400 46880
rect 87240 46880 87400 47040
rect 87240 47040 87400 47200
rect 87240 47200 87400 47360
rect 87240 47360 87400 47520
rect 87240 47520 87400 47680
rect 87240 47680 87400 47840
rect 87240 47840 87400 48000
rect 87240 48000 87400 48160
rect 87240 48160 87400 48320
rect 87240 48320 87400 48480
rect 87240 48480 87400 48640
rect 87240 48640 87400 48800
rect 87240 48800 87400 48960
rect 87240 48960 87400 49120
rect 87240 49120 87400 49280
rect 87240 49280 87400 49440
rect 87240 49440 87400 49600
rect 87240 49600 87400 49760
rect 87240 49760 87400 49920
rect 87240 49920 87400 50080
rect 87240 50080 87400 50240
rect 87240 50240 87400 50400
rect 87240 50400 87400 50560
rect 87240 50560 87400 50720
rect 87240 50720 87400 50880
rect 87240 50880 87400 51040
rect 87240 51040 87400 51200
rect 87400 46080 87560 46240
rect 87400 46240 87560 46400
rect 87400 46400 87560 46560
rect 87400 46560 87560 46720
rect 87400 46720 87560 46880
rect 87400 46880 87560 47040
rect 87400 47040 87560 47200
rect 87400 47200 87560 47360
rect 87400 47360 87560 47520
rect 87400 47520 87560 47680
rect 87400 47680 87560 47840
rect 87400 47840 87560 48000
rect 87400 48000 87560 48160
rect 87400 48160 87560 48320
rect 87400 48320 87560 48480
rect 87400 48480 87560 48640
rect 87400 48640 87560 48800
rect 87400 48800 87560 48960
rect 87400 48960 87560 49120
rect 87400 49120 87560 49280
rect 87400 49280 87560 49440
rect 87400 49440 87560 49600
rect 87400 49600 87560 49760
rect 87400 49760 87560 49920
rect 87400 49920 87560 50080
rect 87400 50080 87560 50240
rect 87400 50240 87560 50400
rect 87400 50400 87560 50560
rect 87400 50560 87560 50720
rect 87400 50720 87560 50880
rect 87400 50880 87560 51040
rect 87400 51040 87560 51200
rect 87400 51200 87560 51360
rect 87560 45760 87720 45920
rect 87560 45920 87720 46080
rect 87560 46080 87720 46240
rect 87560 46240 87720 46400
rect 87560 46400 87720 46560
rect 87560 46560 87720 46720
rect 87560 46720 87720 46880
rect 87560 46880 87720 47040
rect 87560 47040 87720 47200
rect 87560 47200 87720 47360
rect 87560 47360 87720 47520
rect 87560 47520 87720 47680
rect 87560 47680 87720 47840
rect 87560 47840 87720 48000
rect 87560 48000 87720 48160
rect 87560 48160 87720 48320
rect 87560 48320 87720 48480
rect 87560 48480 87720 48640
rect 87560 48640 87720 48800
rect 87560 48800 87720 48960
rect 87560 48960 87720 49120
rect 87560 49120 87720 49280
rect 87560 49280 87720 49440
rect 87560 49440 87720 49600
rect 87560 49600 87720 49760
rect 87560 49760 87720 49920
rect 87560 49920 87720 50080
rect 87560 50080 87720 50240
rect 87560 50240 87720 50400
rect 87560 50400 87720 50560
rect 87560 50560 87720 50720
rect 87560 50720 87720 50880
rect 87560 50880 87720 51040
rect 87560 51040 87720 51200
rect 87560 51200 87720 51360
rect 87560 51360 87720 51520
rect 87720 45760 87880 45920
rect 87720 45920 87880 46080
rect 87720 46080 87880 46240
rect 87720 46240 87880 46400
rect 87720 46400 87880 46560
rect 87720 46560 87880 46720
rect 87720 46720 87880 46880
rect 87720 46880 87880 47040
rect 87720 47040 87880 47200
rect 87720 47200 87880 47360
rect 87720 47360 87880 47520
rect 87720 47520 87880 47680
rect 87720 47680 87880 47840
rect 87720 47840 87880 48000
rect 87720 48000 87880 48160
rect 87720 48160 87880 48320
rect 87720 48320 87880 48480
rect 87720 48480 87880 48640
rect 87720 48640 87880 48800
rect 87720 48800 87880 48960
rect 87720 48960 87880 49120
rect 87720 49120 87880 49280
rect 87720 49280 87880 49440
rect 87720 49440 87880 49600
rect 87720 49600 87880 49760
rect 87720 49760 87880 49920
rect 87720 49920 87880 50080
rect 87720 50080 87880 50240
rect 87720 50240 87880 50400
rect 87720 50400 87880 50560
rect 87720 50560 87880 50720
rect 87720 50720 87880 50880
rect 87720 50880 87880 51040
rect 87720 51040 87880 51200
rect 87720 51200 87880 51360
rect 87720 51360 87880 51520
rect 87720 51520 87880 51680
rect 87880 45600 88040 45760
rect 87880 45760 88040 45920
rect 87880 45920 88040 46080
rect 87880 46080 88040 46240
rect 87880 46240 88040 46400
rect 87880 46400 88040 46560
rect 87880 46560 88040 46720
rect 87880 46720 88040 46880
rect 87880 46880 88040 47040
rect 87880 47040 88040 47200
rect 87880 47200 88040 47360
rect 87880 47360 88040 47520
rect 87880 47520 88040 47680
rect 87880 47680 88040 47840
rect 87880 47840 88040 48000
rect 87880 48000 88040 48160
rect 87880 48160 88040 48320
rect 87880 48320 88040 48480
rect 87880 48480 88040 48640
rect 87880 48640 88040 48800
rect 87880 48800 88040 48960
rect 87880 48960 88040 49120
rect 87880 49120 88040 49280
rect 87880 49280 88040 49440
rect 87880 49440 88040 49600
rect 87880 49600 88040 49760
rect 87880 49760 88040 49920
rect 87880 49920 88040 50080
rect 87880 50080 88040 50240
rect 87880 50240 88040 50400
rect 87880 50400 88040 50560
rect 87880 50560 88040 50720
rect 87880 50720 88040 50880
rect 87880 50880 88040 51040
rect 87880 51040 88040 51200
rect 87880 51200 88040 51360
rect 87880 51360 88040 51520
rect 87880 51520 88040 51680
rect 88040 45440 88200 45600
rect 88040 45600 88200 45760
rect 88040 45760 88200 45920
rect 88040 45920 88200 46080
rect 88040 46080 88200 46240
rect 88040 46240 88200 46400
rect 88040 46400 88200 46560
rect 88040 46560 88200 46720
rect 88040 46720 88200 46880
rect 88040 46880 88200 47040
rect 88040 47040 88200 47200
rect 88040 47200 88200 47360
rect 88040 47360 88200 47520
rect 88040 47520 88200 47680
rect 88040 47680 88200 47840
rect 88040 47840 88200 48000
rect 88040 48000 88200 48160
rect 88040 48160 88200 48320
rect 88040 48320 88200 48480
rect 88040 48480 88200 48640
rect 88040 48640 88200 48800
rect 88040 48800 88200 48960
rect 88040 48960 88200 49120
rect 88040 49120 88200 49280
rect 88040 49280 88200 49440
rect 88040 49440 88200 49600
rect 88040 49600 88200 49760
rect 88040 49760 88200 49920
rect 88040 49920 88200 50080
rect 88040 50080 88200 50240
rect 88040 50240 88200 50400
rect 88040 50400 88200 50560
rect 88040 50560 88200 50720
rect 88040 50720 88200 50880
rect 88040 50880 88200 51040
rect 88040 51040 88200 51200
rect 88040 51200 88200 51360
rect 88040 51360 88200 51520
rect 88040 51520 88200 51680
rect 88040 51680 88200 51840
rect 88200 45280 88360 45440
rect 88200 45440 88360 45600
rect 88200 45600 88360 45760
rect 88200 45760 88360 45920
rect 88200 45920 88360 46080
rect 88200 46080 88360 46240
rect 88200 46240 88360 46400
rect 88200 46400 88360 46560
rect 88200 46560 88360 46720
rect 88200 46720 88360 46880
rect 88200 46880 88360 47040
rect 88200 47040 88360 47200
rect 88200 47200 88360 47360
rect 88200 47360 88360 47520
rect 88200 47520 88360 47680
rect 88200 47680 88360 47840
rect 88200 47840 88360 48000
rect 88200 48000 88360 48160
rect 88200 48160 88360 48320
rect 88200 48320 88360 48480
rect 88200 48480 88360 48640
rect 88200 48640 88360 48800
rect 88200 48800 88360 48960
rect 88200 48960 88360 49120
rect 88200 49120 88360 49280
rect 88200 49280 88360 49440
rect 88200 49440 88360 49600
rect 88200 49600 88360 49760
rect 88200 49760 88360 49920
rect 88200 49920 88360 50080
rect 88200 50080 88360 50240
rect 88200 50240 88360 50400
rect 88200 50400 88360 50560
rect 88200 50560 88360 50720
rect 88200 50720 88360 50880
rect 88200 50880 88360 51040
rect 88200 51040 88360 51200
rect 88200 51200 88360 51360
rect 88200 51360 88360 51520
rect 88200 51520 88360 51680
rect 88200 51680 88360 51840
rect 88200 51840 88360 52000
rect 88360 45280 88520 45440
rect 88360 45440 88520 45600
rect 88360 45600 88520 45760
rect 88360 45760 88520 45920
rect 88360 45920 88520 46080
rect 88360 46080 88520 46240
rect 88360 46240 88520 46400
rect 88360 46400 88520 46560
rect 88360 46560 88520 46720
rect 88360 46720 88520 46880
rect 88360 46880 88520 47040
rect 88360 47040 88520 47200
rect 88360 47200 88520 47360
rect 88360 47360 88520 47520
rect 88360 47520 88520 47680
rect 88360 47680 88520 47840
rect 88360 47840 88520 48000
rect 88360 48000 88520 48160
rect 88360 48160 88520 48320
rect 88360 48320 88520 48480
rect 88360 48480 88520 48640
rect 88360 48640 88520 48800
rect 88360 48800 88520 48960
rect 88360 48960 88520 49120
rect 88360 49120 88520 49280
rect 88360 49280 88520 49440
rect 88360 49440 88520 49600
rect 88360 49600 88520 49760
rect 88360 49760 88520 49920
rect 88360 49920 88520 50080
rect 88360 50080 88520 50240
rect 88360 50240 88520 50400
rect 88360 50400 88520 50560
rect 88360 50560 88520 50720
rect 88360 50720 88520 50880
rect 88360 50880 88520 51040
rect 88360 51040 88520 51200
rect 88360 51200 88520 51360
rect 88360 51360 88520 51520
rect 88360 51520 88520 51680
rect 88360 51680 88520 51840
rect 88360 51840 88520 52000
rect 88520 45120 88680 45280
rect 88520 45280 88680 45440
rect 88520 45440 88680 45600
rect 88520 45600 88680 45760
rect 88520 45760 88680 45920
rect 88520 45920 88680 46080
rect 88520 46080 88680 46240
rect 88520 46240 88680 46400
rect 88520 46400 88680 46560
rect 88520 46560 88680 46720
rect 88520 46720 88680 46880
rect 88520 46880 88680 47040
rect 88520 47040 88680 47200
rect 88520 47200 88680 47360
rect 88520 47360 88680 47520
rect 88520 47520 88680 47680
rect 88520 47680 88680 47840
rect 88520 47840 88680 48000
rect 88520 48000 88680 48160
rect 88520 48160 88680 48320
rect 88520 48320 88680 48480
rect 88520 48480 88680 48640
rect 88520 48640 88680 48800
rect 88520 48800 88680 48960
rect 88520 48960 88680 49120
rect 88520 49120 88680 49280
rect 88520 49280 88680 49440
rect 88520 49440 88680 49600
rect 88520 49600 88680 49760
rect 88520 49760 88680 49920
rect 88520 49920 88680 50080
rect 88520 50080 88680 50240
rect 88520 50240 88680 50400
rect 88520 50400 88680 50560
rect 88520 50560 88680 50720
rect 88520 50720 88680 50880
rect 88520 50880 88680 51040
rect 88520 51040 88680 51200
rect 88520 51200 88680 51360
rect 88520 51360 88680 51520
rect 88520 51520 88680 51680
rect 88520 51680 88680 51840
rect 88520 51840 88680 52000
rect 88520 52000 88680 52160
rect 88680 45120 88840 45280
rect 88680 45280 88840 45440
rect 88680 45440 88840 45600
rect 88680 45600 88840 45760
rect 88680 45760 88840 45920
rect 88680 45920 88840 46080
rect 88680 46080 88840 46240
rect 88680 46240 88840 46400
rect 88680 46400 88840 46560
rect 88680 46560 88840 46720
rect 88680 46720 88840 46880
rect 88680 46880 88840 47040
rect 88680 47040 88840 47200
rect 88680 47200 88840 47360
rect 88680 47360 88840 47520
rect 88680 47520 88840 47680
rect 88680 47680 88840 47840
rect 88680 47840 88840 48000
rect 88680 48000 88840 48160
rect 88680 48160 88840 48320
rect 88680 48320 88840 48480
rect 88680 48480 88840 48640
rect 88680 48640 88840 48800
rect 88680 48800 88840 48960
rect 88680 48960 88840 49120
rect 88680 49120 88840 49280
rect 88680 49280 88840 49440
rect 88680 49440 88840 49600
rect 88680 49600 88840 49760
rect 88680 49760 88840 49920
rect 88680 49920 88840 50080
rect 88680 50080 88840 50240
rect 88680 50240 88840 50400
rect 88680 50400 88840 50560
rect 88680 50560 88840 50720
rect 88680 50720 88840 50880
rect 88680 50880 88840 51040
rect 88680 51040 88840 51200
rect 88680 51200 88840 51360
rect 88680 51360 88840 51520
rect 88680 51520 88840 51680
rect 88680 51680 88840 51840
rect 88680 51840 88840 52000
rect 88680 52000 88840 52160
rect 88840 44960 89000 45120
rect 88840 45120 89000 45280
rect 88840 45280 89000 45440
rect 88840 45440 89000 45600
rect 88840 45600 89000 45760
rect 88840 45760 89000 45920
rect 88840 45920 89000 46080
rect 88840 46080 89000 46240
rect 88840 46240 89000 46400
rect 88840 46400 89000 46560
rect 88840 46560 89000 46720
rect 88840 46720 89000 46880
rect 88840 46880 89000 47040
rect 88840 47040 89000 47200
rect 88840 47200 89000 47360
rect 88840 47360 89000 47520
rect 88840 47520 89000 47680
rect 88840 47680 89000 47840
rect 88840 47840 89000 48000
rect 88840 48000 89000 48160
rect 88840 48160 89000 48320
rect 88840 48320 89000 48480
rect 88840 48480 89000 48640
rect 88840 48640 89000 48800
rect 88840 48800 89000 48960
rect 88840 48960 89000 49120
rect 88840 49120 89000 49280
rect 88840 49280 89000 49440
rect 88840 49440 89000 49600
rect 88840 49600 89000 49760
rect 88840 49760 89000 49920
rect 88840 49920 89000 50080
rect 88840 50080 89000 50240
rect 88840 50240 89000 50400
rect 88840 50400 89000 50560
rect 88840 50560 89000 50720
rect 88840 50720 89000 50880
rect 88840 50880 89000 51040
rect 88840 51040 89000 51200
rect 88840 51200 89000 51360
rect 88840 51360 89000 51520
rect 88840 51520 89000 51680
rect 88840 51680 89000 51840
rect 88840 51840 89000 52000
rect 88840 52000 89000 52160
rect 89000 44800 89160 44960
rect 89000 44960 89160 45120
rect 89000 45120 89160 45280
rect 89000 45280 89160 45440
rect 89000 45440 89160 45600
rect 89000 45600 89160 45760
rect 89000 45760 89160 45920
rect 89000 45920 89160 46080
rect 89000 46080 89160 46240
rect 89000 46240 89160 46400
rect 89000 46400 89160 46560
rect 89000 46560 89160 46720
rect 89000 46720 89160 46880
rect 89000 46880 89160 47040
rect 89000 47040 89160 47200
rect 89000 47200 89160 47360
rect 89000 47360 89160 47520
rect 89000 47520 89160 47680
rect 89000 47680 89160 47840
rect 89000 47840 89160 48000
rect 89000 48000 89160 48160
rect 89000 48160 89160 48320
rect 89000 48320 89160 48480
rect 89000 48960 89160 49120
rect 89000 49120 89160 49280
rect 89000 49280 89160 49440
rect 89000 49440 89160 49600
rect 89000 49600 89160 49760
rect 89000 49760 89160 49920
rect 89000 49920 89160 50080
rect 89000 50080 89160 50240
rect 89000 50240 89160 50400
rect 89000 50400 89160 50560
rect 89000 50560 89160 50720
rect 89000 50720 89160 50880
rect 89000 50880 89160 51040
rect 89000 51040 89160 51200
rect 89000 51200 89160 51360
rect 89000 51360 89160 51520
rect 89000 51520 89160 51680
rect 89000 51680 89160 51840
rect 89000 51840 89160 52000
rect 89000 52000 89160 52160
rect 89000 52160 89160 52320
rect 89160 44800 89320 44960
rect 89160 44960 89320 45120
rect 89160 45120 89320 45280
rect 89160 45280 89320 45440
rect 89160 45440 89320 45600
rect 89160 45600 89320 45760
rect 89160 45760 89320 45920
rect 89160 45920 89320 46080
rect 89160 46080 89320 46240
rect 89160 46240 89320 46400
rect 89160 46400 89320 46560
rect 89160 46560 89320 46720
rect 89160 46720 89320 46880
rect 89160 46880 89320 47040
rect 89160 47040 89320 47200
rect 89160 47200 89320 47360
rect 89160 47360 89320 47520
rect 89160 47520 89320 47680
rect 89160 47680 89320 47840
rect 89160 47840 89320 48000
rect 89160 48000 89320 48160
rect 89160 49280 89320 49440
rect 89160 49440 89320 49600
rect 89160 49600 89320 49760
rect 89160 49760 89320 49920
rect 89160 49920 89320 50080
rect 89160 50080 89320 50240
rect 89160 50240 89320 50400
rect 89160 50400 89320 50560
rect 89160 50560 89320 50720
rect 89160 50720 89320 50880
rect 89160 50880 89320 51040
rect 89160 51040 89320 51200
rect 89160 51200 89320 51360
rect 89160 51360 89320 51520
rect 89160 51520 89320 51680
rect 89160 51680 89320 51840
rect 89160 51840 89320 52000
rect 89160 52000 89320 52160
rect 89160 52160 89320 52320
rect 89320 44640 89480 44800
rect 89320 44800 89480 44960
rect 89320 44960 89480 45120
rect 89320 45120 89480 45280
rect 89320 45280 89480 45440
rect 89320 45440 89480 45600
rect 89320 45600 89480 45760
rect 89320 45760 89480 45920
rect 89320 45920 89480 46080
rect 89320 46080 89480 46240
rect 89320 46240 89480 46400
rect 89320 46400 89480 46560
rect 89320 46560 89480 46720
rect 89320 46720 89480 46880
rect 89320 46880 89480 47040
rect 89320 47040 89480 47200
rect 89320 47200 89480 47360
rect 89320 47360 89480 47520
rect 89320 47520 89480 47680
rect 89320 47680 89480 47840
rect 89320 47840 89480 48000
rect 89320 49440 89480 49600
rect 89320 49600 89480 49760
rect 89320 49760 89480 49920
rect 89320 49920 89480 50080
rect 89320 50080 89480 50240
rect 89320 50240 89480 50400
rect 89320 50400 89480 50560
rect 89320 50560 89480 50720
rect 89320 50720 89480 50880
rect 89320 50880 89480 51040
rect 89320 51040 89480 51200
rect 89320 51200 89480 51360
rect 89320 51360 89480 51520
rect 89320 51520 89480 51680
rect 89320 51680 89480 51840
rect 89320 51840 89480 52000
rect 89320 52000 89480 52160
rect 89320 52160 89480 52320
rect 89480 44640 89640 44800
rect 89480 44800 89640 44960
rect 89480 44960 89640 45120
rect 89480 45120 89640 45280
rect 89480 45280 89640 45440
rect 89480 45440 89640 45600
rect 89480 45600 89640 45760
rect 89480 45760 89640 45920
rect 89480 45920 89640 46080
rect 89480 46080 89640 46240
rect 89480 46240 89640 46400
rect 89480 46400 89640 46560
rect 89480 46560 89640 46720
rect 89480 46720 89640 46880
rect 89480 46880 89640 47040
rect 89480 47040 89640 47200
rect 89480 47200 89640 47360
rect 89480 47360 89640 47520
rect 89480 47520 89640 47680
rect 89480 47680 89640 47840
rect 89480 49600 89640 49760
rect 89480 49760 89640 49920
rect 89480 49920 89640 50080
rect 89480 50080 89640 50240
rect 89480 50240 89640 50400
rect 89480 50400 89640 50560
rect 89480 50560 89640 50720
rect 89480 50720 89640 50880
rect 89480 50880 89640 51040
rect 89480 51040 89640 51200
rect 89480 51200 89640 51360
rect 89480 51360 89640 51520
rect 89480 51520 89640 51680
rect 89480 51680 89640 51840
rect 89480 51840 89640 52000
rect 89480 52000 89640 52160
rect 89480 52160 89640 52320
rect 89640 44480 89800 44640
rect 89640 44640 89800 44800
rect 89640 44800 89800 44960
rect 89640 44960 89800 45120
rect 89640 45120 89800 45280
rect 89640 45280 89800 45440
rect 89640 45440 89800 45600
rect 89640 45600 89800 45760
rect 89640 45760 89800 45920
rect 89640 45920 89800 46080
rect 89640 46080 89800 46240
rect 89640 46240 89800 46400
rect 89640 46400 89800 46560
rect 89640 46560 89800 46720
rect 89640 46720 89800 46880
rect 89640 46880 89800 47040
rect 89640 47040 89800 47200
rect 89640 47200 89800 47360
rect 89640 47360 89800 47520
rect 89640 47520 89800 47680
rect 89640 47680 89800 47840
rect 89640 49760 89800 49920
rect 89640 49920 89800 50080
rect 89640 50080 89800 50240
rect 89640 50240 89800 50400
rect 89640 50400 89800 50560
rect 89640 50560 89800 50720
rect 89640 50720 89800 50880
rect 89640 50880 89800 51040
rect 89640 51040 89800 51200
rect 89640 51200 89800 51360
rect 89640 51360 89800 51520
rect 89640 51520 89800 51680
rect 89640 51680 89800 51840
rect 89640 51840 89800 52000
rect 89640 52000 89800 52160
rect 89640 52160 89800 52320
rect 89640 52320 89800 52480
rect 89800 44320 89960 44480
rect 89800 44480 89960 44640
rect 89800 44640 89960 44800
rect 89800 44800 89960 44960
rect 89800 44960 89960 45120
rect 89800 45120 89960 45280
rect 89800 45280 89960 45440
rect 89800 45440 89960 45600
rect 89800 45600 89960 45760
rect 89800 45760 89960 45920
rect 89800 45920 89960 46080
rect 89800 46080 89960 46240
rect 89800 46240 89960 46400
rect 89800 46400 89960 46560
rect 89800 46560 89960 46720
rect 89800 46720 89960 46880
rect 89800 46880 89960 47040
rect 89800 47040 89960 47200
rect 89800 47200 89960 47360
rect 89800 47360 89960 47520
rect 89800 47520 89960 47680
rect 89800 49760 89960 49920
rect 89800 49920 89960 50080
rect 89800 50080 89960 50240
rect 89800 50240 89960 50400
rect 89800 50400 89960 50560
rect 89800 50560 89960 50720
rect 89800 50720 89960 50880
rect 89800 50880 89960 51040
rect 89800 51040 89960 51200
rect 89800 51200 89960 51360
rect 89800 51360 89960 51520
rect 89800 51520 89960 51680
rect 89800 51680 89960 51840
rect 89800 51840 89960 52000
rect 89800 52000 89960 52160
rect 89800 52160 89960 52320
rect 89800 52320 89960 52480
rect 89960 44160 90120 44320
rect 89960 44320 90120 44480
rect 89960 44480 90120 44640
rect 89960 44640 90120 44800
rect 89960 44800 90120 44960
rect 89960 44960 90120 45120
rect 89960 45120 90120 45280
rect 89960 45280 90120 45440
rect 89960 45440 90120 45600
rect 89960 45600 90120 45760
rect 89960 45760 90120 45920
rect 89960 45920 90120 46080
rect 89960 46080 90120 46240
rect 89960 46240 90120 46400
rect 89960 46400 90120 46560
rect 89960 46560 90120 46720
rect 89960 46720 90120 46880
rect 89960 46880 90120 47040
rect 89960 47040 90120 47200
rect 89960 47200 90120 47360
rect 89960 47360 90120 47520
rect 89960 47520 90120 47680
rect 89960 49920 90120 50080
rect 89960 50080 90120 50240
rect 89960 50240 90120 50400
rect 89960 50400 90120 50560
rect 89960 50560 90120 50720
rect 89960 50720 90120 50880
rect 89960 50880 90120 51040
rect 89960 51040 90120 51200
rect 89960 51200 90120 51360
rect 89960 51360 90120 51520
rect 89960 51520 90120 51680
rect 89960 51680 90120 51840
rect 89960 51840 90120 52000
rect 89960 52000 90120 52160
rect 89960 52160 90120 52320
rect 89960 52320 90120 52480
rect 90120 44000 90280 44160
rect 90120 44160 90280 44320
rect 90120 44320 90280 44480
rect 90120 44480 90280 44640
rect 90120 44640 90280 44800
rect 90120 44800 90280 44960
rect 90120 44960 90280 45120
rect 90120 45120 90280 45280
rect 90120 45280 90280 45440
rect 90120 45440 90280 45600
rect 90120 45600 90280 45760
rect 90120 45760 90280 45920
rect 90120 45920 90280 46080
rect 90120 46080 90280 46240
rect 90120 46240 90280 46400
rect 90120 46400 90280 46560
rect 90120 46560 90280 46720
rect 90120 46720 90280 46880
rect 90120 46880 90280 47040
rect 90120 47040 90280 47200
rect 90120 47200 90280 47360
rect 90120 47360 90280 47520
rect 90120 49920 90280 50080
rect 90120 50080 90280 50240
rect 90120 50240 90280 50400
rect 90120 50400 90280 50560
rect 90120 50560 90280 50720
rect 90120 50720 90280 50880
rect 90120 50880 90280 51040
rect 90120 51040 90280 51200
rect 90120 51200 90280 51360
rect 90120 51360 90280 51520
rect 90120 51520 90280 51680
rect 90120 51680 90280 51840
rect 90120 51840 90280 52000
rect 90120 52000 90280 52160
rect 90120 52160 90280 52320
rect 90120 52320 90280 52480
rect 90280 43680 90440 43840
rect 90280 43840 90440 44000
rect 90280 44000 90440 44160
rect 90280 44160 90440 44320
rect 90280 44320 90440 44480
rect 90280 44480 90440 44640
rect 90280 44640 90440 44800
rect 90280 44800 90440 44960
rect 90280 44960 90440 45120
rect 90280 45120 90440 45280
rect 90280 45280 90440 45440
rect 90280 45440 90440 45600
rect 90280 45600 90440 45760
rect 90280 45760 90440 45920
rect 90280 45920 90440 46080
rect 90280 46080 90440 46240
rect 90280 46240 90440 46400
rect 90280 46400 90440 46560
rect 90280 46560 90440 46720
rect 90280 46720 90440 46880
rect 90280 46880 90440 47040
rect 90280 47040 90440 47200
rect 90280 47200 90440 47360
rect 90280 47360 90440 47520
rect 90280 49920 90440 50080
rect 90280 50080 90440 50240
rect 90280 50240 90440 50400
rect 90280 50400 90440 50560
rect 90280 50560 90440 50720
rect 90280 50720 90440 50880
rect 90280 50880 90440 51040
rect 90280 51040 90440 51200
rect 90280 51200 90440 51360
rect 90280 51360 90440 51520
rect 90280 51520 90440 51680
rect 90280 51680 90440 51840
rect 90280 51840 90440 52000
rect 90280 52000 90440 52160
rect 90280 52160 90440 52320
rect 90280 52320 90440 52480
rect 90440 43360 90600 43520
rect 90440 43520 90600 43680
rect 90440 43680 90600 43840
rect 90440 43840 90600 44000
rect 90440 44000 90600 44160
rect 90440 44160 90600 44320
rect 90440 44320 90600 44480
rect 90440 44480 90600 44640
rect 90440 44640 90600 44800
rect 90440 44800 90600 44960
rect 90440 44960 90600 45120
rect 90440 45120 90600 45280
rect 90440 45280 90600 45440
rect 90440 45440 90600 45600
rect 90440 45600 90600 45760
rect 90440 45760 90600 45920
rect 90440 45920 90600 46080
rect 90440 46080 90600 46240
rect 90440 46240 90600 46400
rect 90440 46400 90600 46560
rect 90440 46560 90600 46720
rect 90440 46720 90600 46880
rect 90440 46880 90600 47040
rect 90440 47040 90600 47200
rect 90440 47200 90600 47360
rect 90440 47360 90600 47520
rect 90440 49920 90600 50080
rect 90440 50080 90600 50240
rect 90440 50240 90600 50400
rect 90440 50400 90600 50560
rect 90440 50560 90600 50720
rect 90440 50720 90600 50880
rect 90440 50880 90600 51040
rect 90440 51040 90600 51200
rect 90440 51200 90600 51360
rect 90440 51360 90600 51520
rect 90440 51520 90600 51680
rect 90440 51680 90600 51840
rect 90440 51840 90600 52000
rect 90440 52000 90600 52160
rect 90440 52160 90600 52320
rect 90440 52320 90600 52480
rect 90600 43200 90760 43360
rect 90600 43360 90760 43520
rect 90600 43520 90760 43680
rect 90600 43680 90760 43840
rect 90600 43840 90760 44000
rect 90600 44000 90760 44160
rect 90600 44160 90760 44320
rect 90600 44320 90760 44480
rect 90600 44480 90760 44640
rect 90600 44640 90760 44800
rect 90600 44800 90760 44960
rect 90600 44960 90760 45120
rect 90600 45120 90760 45280
rect 90600 45280 90760 45440
rect 90600 45440 90760 45600
rect 90600 45600 90760 45760
rect 90600 45760 90760 45920
rect 90600 45920 90760 46080
rect 90600 46080 90760 46240
rect 90600 46240 90760 46400
rect 90600 46400 90760 46560
rect 90600 46560 90760 46720
rect 90600 46720 90760 46880
rect 90600 46880 90760 47040
rect 90600 47040 90760 47200
rect 90600 47200 90760 47360
rect 90600 47360 90760 47520
rect 90600 49920 90760 50080
rect 90600 50080 90760 50240
rect 90600 50240 90760 50400
rect 90600 50400 90760 50560
rect 90600 50560 90760 50720
rect 90600 50720 90760 50880
rect 90600 50880 90760 51040
rect 90600 51040 90760 51200
rect 90600 51200 90760 51360
rect 90600 51360 90760 51520
rect 90600 51520 90760 51680
rect 90600 51680 90760 51840
rect 90600 51840 90760 52000
rect 90600 52000 90760 52160
rect 90600 52160 90760 52320
rect 90600 52320 90760 52480
rect 90760 42720 90920 42880
rect 90760 42880 90920 43040
rect 90760 43040 90920 43200
rect 90760 43200 90920 43360
rect 90760 43360 90920 43520
rect 90760 43520 90920 43680
rect 90760 43680 90920 43840
rect 90760 43840 90920 44000
rect 90760 44000 90920 44160
rect 90760 44160 90920 44320
rect 90760 44320 90920 44480
rect 90760 44480 90920 44640
rect 90760 44640 90920 44800
rect 90760 44800 90920 44960
rect 90760 44960 90920 45120
rect 90760 45120 90920 45280
rect 90760 45280 90920 45440
rect 90760 45440 90920 45600
rect 90760 45600 90920 45760
rect 90760 45760 90920 45920
rect 90760 45920 90920 46080
rect 90760 46080 90920 46240
rect 90760 46240 90920 46400
rect 90760 46400 90920 46560
rect 90760 46560 90920 46720
rect 90760 46720 90920 46880
rect 90760 46880 90920 47040
rect 90760 47040 90920 47200
rect 90760 47200 90920 47360
rect 90760 47360 90920 47520
rect 90760 49920 90920 50080
rect 90760 50080 90920 50240
rect 90760 50240 90920 50400
rect 90760 50400 90920 50560
rect 90760 50560 90920 50720
rect 90760 50720 90920 50880
rect 90760 50880 90920 51040
rect 90760 51040 90920 51200
rect 90760 51200 90920 51360
rect 90760 51360 90920 51520
rect 90760 51520 90920 51680
rect 90760 51680 90920 51840
rect 90760 51840 90920 52000
rect 90760 52000 90920 52160
rect 90760 52160 90920 52320
rect 90760 52320 90920 52480
rect 90920 42400 91080 42560
rect 90920 42560 91080 42720
rect 90920 42720 91080 42880
rect 90920 42880 91080 43040
rect 90920 43040 91080 43200
rect 90920 43200 91080 43360
rect 90920 43360 91080 43520
rect 90920 43520 91080 43680
rect 90920 43680 91080 43840
rect 90920 43840 91080 44000
rect 90920 44000 91080 44160
rect 90920 44160 91080 44320
rect 90920 44320 91080 44480
rect 90920 44480 91080 44640
rect 90920 44640 91080 44800
rect 90920 44800 91080 44960
rect 90920 44960 91080 45120
rect 90920 45120 91080 45280
rect 90920 45280 91080 45440
rect 90920 45440 91080 45600
rect 90920 45600 91080 45760
rect 90920 45760 91080 45920
rect 90920 45920 91080 46080
rect 90920 46080 91080 46240
rect 90920 46240 91080 46400
rect 90920 46400 91080 46560
rect 90920 46560 91080 46720
rect 90920 46720 91080 46880
rect 90920 46880 91080 47040
rect 90920 47040 91080 47200
rect 90920 47200 91080 47360
rect 90920 47360 91080 47520
rect 90920 49760 91080 49920
rect 90920 49920 91080 50080
rect 90920 50080 91080 50240
rect 90920 50240 91080 50400
rect 90920 50400 91080 50560
rect 90920 50560 91080 50720
rect 90920 50720 91080 50880
rect 90920 50880 91080 51040
rect 90920 51040 91080 51200
rect 90920 51200 91080 51360
rect 90920 51360 91080 51520
rect 90920 51520 91080 51680
rect 90920 51680 91080 51840
rect 90920 51840 91080 52000
rect 90920 52000 91080 52160
rect 90920 52160 91080 52320
rect 90920 52320 91080 52480
rect 91080 42080 91240 42240
rect 91080 42240 91240 42400
rect 91080 42400 91240 42560
rect 91080 42560 91240 42720
rect 91080 42720 91240 42880
rect 91080 42880 91240 43040
rect 91080 43040 91240 43200
rect 91080 43200 91240 43360
rect 91080 43360 91240 43520
rect 91080 43520 91240 43680
rect 91080 43680 91240 43840
rect 91080 43840 91240 44000
rect 91080 44000 91240 44160
rect 91080 44160 91240 44320
rect 91080 44320 91240 44480
rect 91080 44480 91240 44640
rect 91080 44640 91240 44800
rect 91080 44800 91240 44960
rect 91080 44960 91240 45120
rect 91080 45120 91240 45280
rect 91080 45280 91240 45440
rect 91080 45440 91240 45600
rect 91080 45600 91240 45760
rect 91080 45760 91240 45920
rect 91080 45920 91240 46080
rect 91080 46080 91240 46240
rect 91080 46240 91240 46400
rect 91080 46400 91240 46560
rect 91080 46560 91240 46720
rect 91080 46720 91240 46880
rect 91080 46880 91240 47040
rect 91080 47040 91240 47200
rect 91080 47200 91240 47360
rect 91080 47360 91240 47520
rect 91080 49600 91240 49760
rect 91080 49760 91240 49920
rect 91080 49920 91240 50080
rect 91080 50080 91240 50240
rect 91080 50240 91240 50400
rect 91080 50400 91240 50560
rect 91080 50560 91240 50720
rect 91080 50720 91240 50880
rect 91080 50880 91240 51040
rect 91080 51040 91240 51200
rect 91080 51200 91240 51360
rect 91080 51360 91240 51520
rect 91080 51520 91240 51680
rect 91080 51680 91240 51840
rect 91080 51840 91240 52000
rect 91080 52000 91240 52160
rect 91080 52160 91240 52320
rect 91080 52320 91240 52480
rect 91240 41600 91400 41760
rect 91240 41760 91400 41920
rect 91240 41920 91400 42080
rect 91240 42080 91400 42240
rect 91240 42240 91400 42400
rect 91240 42400 91400 42560
rect 91240 42560 91400 42720
rect 91240 42720 91400 42880
rect 91240 42880 91400 43040
rect 91240 43040 91400 43200
rect 91240 43200 91400 43360
rect 91240 43360 91400 43520
rect 91240 43520 91400 43680
rect 91240 43680 91400 43840
rect 91240 43840 91400 44000
rect 91240 44000 91400 44160
rect 91240 44160 91400 44320
rect 91240 44320 91400 44480
rect 91240 44480 91400 44640
rect 91240 44640 91400 44800
rect 91240 44800 91400 44960
rect 91240 44960 91400 45120
rect 91240 45120 91400 45280
rect 91240 45280 91400 45440
rect 91240 45440 91400 45600
rect 91240 45600 91400 45760
rect 91240 45760 91400 45920
rect 91240 45920 91400 46080
rect 91240 46080 91400 46240
rect 91240 46240 91400 46400
rect 91240 46400 91400 46560
rect 91240 46560 91400 46720
rect 91240 46720 91400 46880
rect 91240 46880 91400 47040
rect 91240 47040 91400 47200
rect 91240 47200 91400 47360
rect 91240 47360 91400 47520
rect 91240 47520 91400 47680
rect 91240 49280 91400 49440
rect 91240 49440 91400 49600
rect 91240 49600 91400 49760
rect 91240 49760 91400 49920
rect 91240 49920 91400 50080
rect 91240 50080 91400 50240
rect 91240 50240 91400 50400
rect 91240 50400 91400 50560
rect 91240 50560 91400 50720
rect 91240 50720 91400 50880
rect 91240 50880 91400 51040
rect 91240 51040 91400 51200
rect 91240 51200 91400 51360
rect 91240 51360 91400 51520
rect 91240 51520 91400 51680
rect 91240 51680 91400 51840
rect 91240 51840 91400 52000
rect 91240 52000 91400 52160
rect 91240 52160 91400 52320
rect 91400 41280 91560 41440
rect 91400 41440 91560 41600
rect 91400 41600 91560 41760
rect 91400 41760 91560 41920
rect 91400 41920 91560 42080
rect 91400 42080 91560 42240
rect 91400 42240 91560 42400
rect 91400 42400 91560 42560
rect 91400 42560 91560 42720
rect 91400 42720 91560 42880
rect 91400 42880 91560 43040
rect 91400 43040 91560 43200
rect 91400 43200 91560 43360
rect 91400 43360 91560 43520
rect 91400 43520 91560 43680
rect 91400 43680 91560 43840
rect 91400 43840 91560 44000
rect 91400 44000 91560 44160
rect 91400 44160 91560 44320
rect 91400 44320 91560 44480
rect 91400 44480 91560 44640
rect 91400 44640 91560 44800
rect 91400 44800 91560 44960
rect 91400 44960 91560 45120
rect 91400 45120 91560 45280
rect 91400 45280 91560 45440
rect 91400 45440 91560 45600
rect 91400 45600 91560 45760
rect 91400 45760 91560 45920
rect 91400 45920 91560 46080
rect 91400 46080 91560 46240
rect 91400 46240 91560 46400
rect 91400 46400 91560 46560
rect 91400 46560 91560 46720
rect 91400 46720 91560 46880
rect 91400 46880 91560 47040
rect 91400 47040 91560 47200
rect 91400 47200 91560 47360
rect 91400 47360 91560 47520
rect 91400 47520 91560 47680
rect 91400 47680 91560 47840
rect 91400 47840 91560 48000
rect 91400 48000 91560 48160
rect 91400 48480 91560 48640
rect 91400 48800 91560 48960
rect 91400 48960 91560 49120
rect 91400 49120 91560 49280
rect 91400 49280 91560 49440
rect 91400 49440 91560 49600
rect 91400 49600 91560 49760
rect 91400 49760 91560 49920
rect 91400 49920 91560 50080
rect 91400 50080 91560 50240
rect 91400 50240 91560 50400
rect 91400 50400 91560 50560
rect 91400 50560 91560 50720
rect 91400 50720 91560 50880
rect 91400 50880 91560 51040
rect 91400 51040 91560 51200
rect 91400 51200 91560 51360
rect 91400 51360 91560 51520
rect 91400 51520 91560 51680
rect 91400 51680 91560 51840
rect 91400 51840 91560 52000
rect 91400 52000 91560 52160
rect 91400 52160 91560 52320
rect 91560 40800 91720 40960
rect 91560 40960 91720 41120
rect 91560 41120 91720 41280
rect 91560 41280 91720 41440
rect 91560 41440 91720 41600
rect 91560 41600 91720 41760
rect 91560 41760 91720 41920
rect 91560 41920 91720 42080
rect 91560 42080 91720 42240
rect 91560 42240 91720 42400
rect 91560 42400 91720 42560
rect 91560 42560 91720 42720
rect 91560 42720 91720 42880
rect 91560 42880 91720 43040
rect 91560 43040 91720 43200
rect 91560 43200 91720 43360
rect 91560 43360 91720 43520
rect 91560 43520 91720 43680
rect 91560 43680 91720 43840
rect 91560 43840 91720 44000
rect 91560 44000 91720 44160
rect 91560 44160 91720 44320
rect 91560 44320 91720 44480
rect 91560 44480 91720 44640
rect 91560 44640 91720 44800
rect 91560 44800 91720 44960
rect 91560 44960 91720 45120
rect 91560 45120 91720 45280
rect 91560 45280 91720 45440
rect 91560 45440 91720 45600
rect 91560 45600 91720 45760
rect 91560 45760 91720 45920
rect 91560 45920 91720 46080
rect 91560 46080 91720 46240
rect 91560 46240 91720 46400
rect 91560 46400 91720 46560
rect 91560 46560 91720 46720
rect 91560 46720 91720 46880
rect 91560 46880 91720 47040
rect 91560 47040 91720 47200
rect 91560 47200 91720 47360
rect 91560 47360 91720 47520
rect 91560 47520 91720 47680
rect 91560 47680 91720 47840
rect 91560 47840 91720 48000
rect 91560 48000 91720 48160
rect 91560 48160 91720 48320
rect 91560 48320 91720 48480
rect 91560 48480 91720 48640
rect 91560 48640 91720 48800
rect 91560 48800 91720 48960
rect 91560 48960 91720 49120
rect 91560 49120 91720 49280
rect 91560 49280 91720 49440
rect 91560 49440 91720 49600
rect 91560 49600 91720 49760
rect 91560 49760 91720 49920
rect 91560 49920 91720 50080
rect 91560 50080 91720 50240
rect 91560 50240 91720 50400
rect 91560 50400 91720 50560
rect 91560 50560 91720 50720
rect 91560 50720 91720 50880
rect 91560 50880 91720 51040
rect 91560 51040 91720 51200
rect 91560 51200 91720 51360
rect 91560 51360 91720 51520
rect 91560 51520 91720 51680
rect 91560 51680 91720 51840
rect 91560 51840 91720 52000
rect 91560 52000 91720 52160
rect 91560 52160 91720 52320
rect 91720 40320 91880 40480
rect 91720 40480 91880 40640
rect 91720 40640 91880 40800
rect 91720 40800 91880 40960
rect 91720 40960 91880 41120
rect 91720 41120 91880 41280
rect 91720 41280 91880 41440
rect 91720 41440 91880 41600
rect 91720 41600 91880 41760
rect 91720 41760 91880 41920
rect 91720 41920 91880 42080
rect 91720 42080 91880 42240
rect 91720 42240 91880 42400
rect 91720 42400 91880 42560
rect 91720 42560 91880 42720
rect 91720 42720 91880 42880
rect 91720 42880 91880 43040
rect 91720 43040 91880 43200
rect 91720 43200 91880 43360
rect 91720 43360 91880 43520
rect 91720 43520 91880 43680
rect 91720 43680 91880 43840
rect 91720 43840 91880 44000
rect 91720 44000 91880 44160
rect 91720 44160 91880 44320
rect 91720 44320 91880 44480
rect 91720 44480 91880 44640
rect 91720 44640 91880 44800
rect 91720 44800 91880 44960
rect 91720 44960 91880 45120
rect 91720 45120 91880 45280
rect 91720 45280 91880 45440
rect 91720 45440 91880 45600
rect 91720 45600 91880 45760
rect 91720 45760 91880 45920
rect 91720 45920 91880 46080
rect 91720 46080 91880 46240
rect 91720 46240 91880 46400
rect 91720 46400 91880 46560
rect 91720 46560 91880 46720
rect 91720 46720 91880 46880
rect 91720 46880 91880 47040
rect 91720 47040 91880 47200
rect 91720 47200 91880 47360
rect 91720 47360 91880 47520
rect 91720 47520 91880 47680
rect 91720 47680 91880 47840
rect 91720 47840 91880 48000
rect 91720 48000 91880 48160
rect 91720 48160 91880 48320
rect 91720 48320 91880 48480
rect 91720 48480 91880 48640
rect 91720 48640 91880 48800
rect 91720 48800 91880 48960
rect 91720 48960 91880 49120
rect 91720 49120 91880 49280
rect 91720 49280 91880 49440
rect 91720 49440 91880 49600
rect 91720 49600 91880 49760
rect 91720 49760 91880 49920
rect 91720 49920 91880 50080
rect 91720 50080 91880 50240
rect 91720 50240 91880 50400
rect 91720 50400 91880 50560
rect 91720 50560 91880 50720
rect 91720 50720 91880 50880
rect 91720 50880 91880 51040
rect 91720 51040 91880 51200
rect 91720 51200 91880 51360
rect 91720 51360 91880 51520
rect 91720 51520 91880 51680
rect 91720 51680 91880 51840
rect 91720 51840 91880 52000
rect 91720 52000 91880 52160
rect 91880 39840 92040 40000
rect 91880 40000 92040 40160
rect 91880 40160 92040 40320
rect 91880 40320 92040 40480
rect 91880 40480 92040 40640
rect 91880 40640 92040 40800
rect 91880 40800 92040 40960
rect 91880 40960 92040 41120
rect 91880 41120 92040 41280
rect 91880 41280 92040 41440
rect 91880 41440 92040 41600
rect 91880 41600 92040 41760
rect 91880 41760 92040 41920
rect 91880 41920 92040 42080
rect 91880 42080 92040 42240
rect 91880 42240 92040 42400
rect 91880 42400 92040 42560
rect 91880 42560 92040 42720
rect 91880 42720 92040 42880
rect 91880 42880 92040 43040
rect 91880 43040 92040 43200
rect 91880 43200 92040 43360
rect 91880 43360 92040 43520
rect 91880 43520 92040 43680
rect 91880 43680 92040 43840
rect 91880 43840 92040 44000
rect 91880 44000 92040 44160
rect 91880 44160 92040 44320
rect 91880 44320 92040 44480
rect 91880 44480 92040 44640
rect 91880 44640 92040 44800
rect 91880 44800 92040 44960
rect 91880 44960 92040 45120
rect 91880 45120 92040 45280
rect 91880 45280 92040 45440
rect 91880 45440 92040 45600
rect 91880 45600 92040 45760
rect 91880 45760 92040 45920
rect 91880 45920 92040 46080
rect 91880 46080 92040 46240
rect 91880 46240 92040 46400
rect 91880 46400 92040 46560
rect 91880 46560 92040 46720
rect 91880 46720 92040 46880
rect 91880 46880 92040 47040
rect 91880 47040 92040 47200
rect 91880 47200 92040 47360
rect 91880 47360 92040 47520
rect 91880 47520 92040 47680
rect 91880 47680 92040 47840
rect 91880 47840 92040 48000
rect 91880 48000 92040 48160
rect 91880 48160 92040 48320
rect 91880 48320 92040 48480
rect 91880 48480 92040 48640
rect 91880 48640 92040 48800
rect 91880 48800 92040 48960
rect 91880 48960 92040 49120
rect 91880 49120 92040 49280
rect 91880 49280 92040 49440
rect 91880 49440 92040 49600
rect 91880 49600 92040 49760
rect 91880 49760 92040 49920
rect 91880 49920 92040 50080
rect 91880 50080 92040 50240
rect 91880 50240 92040 50400
rect 91880 50400 92040 50560
rect 91880 50560 92040 50720
rect 91880 50720 92040 50880
rect 91880 50880 92040 51040
rect 91880 51040 92040 51200
rect 91880 51200 92040 51360
rect 91880 51360 92040 51520
rect 91880 51520 92040 51680
rect 91880 51680 92040 51840
rect 91880 51840 92040 52000
rect 91880 52000 92040 52160
rect 92040 39360 92200 39520
rect 92040 39520 92200 39680
rect 92040 39680 92200 39840
rect 92040 39840 92200 40000
rect 92040 40000 92200 40160
rect 92040 40160 92200 40320
rect 92040 40320 92200 40480
rect 92040 40480 92200 40640
rect 92040 40640 92200 40800
rect 92040 40800 92200 40960
rect 92040 40960 92200 41120
rect 92040 41120 92200 41280
rect 92040 41280 92200 41440
rect 92040 41440 92200 41600
rect 92040 41600 92200 41760
rect 92040 41760 92200 41920
rect 92040 41920 92200 42080
rect 92040 42080 92200 42240
rect 92040 42240 92200 42400
rect 92040 42400 92200 42560
rect 92040 42560 92200 42720
rect 92040 42720 92200 42880
rect 92040 42880 92200 43040
rect 92040 43040 92200 43200
rect 92040 43200 92200 43360
rect 92040 43360 92200 43520
rect 92040 43520 92200 43680
rect 92040 43680 92200 43840
rect 92040 43840 92200 44000
rect 92040 44000 92200 44160
rect 92040 44160 92200 44320
rect 92040 44320 92200 44480
rect 92040 44480 92200 44640
rect 92040 44640 92200 44800
rect 92040 44800 92200 44960
rect 92040 44960 92200 45120
rect 92040 45120 92200 45280
rect 92040 45280 92200 45440
rect 92040 45440 92200 45600
rect 92040 45600 92200 45760
rect 92040 45760 92200 45920
rect 92040 45920 92200 46080
rect 92040 46080 92200 46240
rect 92040 46240 92200 46400
rect 92040 46400 92200 46560
rect 92040 46560 92200 46720
rect 92040 46720 92200 46880
rect 92040 46880 92200 47040
rect 92040 47040 92200 47200
rect 92040 47200 92200 47360
rect 92040 47360 92200 47520
rect 92040 47520 92200 47680
rect 92040 47680 92200 47840
rect 92040 47840 92200 48000
rect 92040 48000 92200 48160
rect 92040 48160 92200 48320
rect 92040 48320 92200 48480
rect 92040 48480 92200 48640
rect 92040 48640 92200 48800
rect 92040 48800 92200 48960
rect 92040 48960 92200 49120
rect 92040 49120 92200 49280
rect 92040 49280 92200 49440
rect 92040 49440 92200 49600
rect 92040 49600 92200 49760
rect 92040 49760 92200 49920
rect 92040 49920 92200 50080
rect 92040 50080 92200 50240
rect 92040 50240 92200 50400
rect 92040 50400 92200 50560
rect 92040 50560 92200 50720
rect 92040 50720 92200 50880
rect 92040 50880 92200 51040
rect 92040 51040 92200 51200
rect 92040 51200 92200 51360
rect 92040 51360 92200 51520
rect 92040 51520 92200 51680
rect 92040 51680 92200 51840
rect 92040 51840 92200 52000
rect 92040 52000 92200 52160
rect 92200 38880 92360 39040
rect 92200 39040 92360 39200
rect 92200 39200 92360 39360
rect 92200 39360 92360 39520
rect 92200 39520 92360 39680
rect 92200 39680 92360 39840
rect 92200 39840 92360 40000
rect 92200 40000 92360 40160
rect 92200 40160 92360 40320
rect 92200 40320 92360 40480
rect 92200 40480 92360 40640
rect 92200 40640 92360 40800
rect 92200 40800 92360 40960
rect 92200 40960 92360 41120
rect 92200 41120 92360 41280
rect 92200 41280 92360 41440
rect 92200 41440 92360 41600
rect 92200 41600 92360 41760
rect 92200 41760 92360 41920
rect 92200 41920 92360 42080
rect 92200 42080 92360 42240
rect 92200 42240 92360 42400
rect 92200 42400 92360 42560
rect 92200 42560 92360 42720
rect 92200 42720 92360 42880
rect 92200 42880 92360 43040
rect 92200 43040 92360 43200
rect 92200 43200 92360 43360
rect 92200 43360 92360 43520
rect 92200 43520 92360 43680
rect 92200 43680 92360 43840
rect 92200 43840 92360 44000
rect 92200 44000 92360 44160
rect 92200 44160 92360 44320
rect 92200 44320 92360 44480
rect 92200 44480 92360 44640
rect 92200 44640 92360 44800
rect 92200 44800 92360 44960
rect 92200 44960 92360 45120
rect 92200 45120 92360 45280
rect 92200 45280 92360 45440
rect 92200 45440 92360 45600
rect 92200 45600 92360 45760
rect 92200 45760 92360 45920
rect 92200 45920 92360 46080
rect 92200 46080 92360 46240
rect 92200 46240 92360 46400
rect 92200 46400 92360 46560
rect 92200 46560 92360 46720
rect 92200 46720 92360 46880
rect 92200 46880 92360 47040
rect 92200 47040 92360 47200
rect 92200 47200 92360 47360
rect 92200 47360 92360 47520
rect 92200 47520 92360 47680
rect 92200 47680 92360 47840
rect 92200 47840 92360 48000
rect 92200 48000 92360 48160
rect 92200 48160 92360 48320
rect 92200 48320 92360 48480
rect 92200 48480 92360 48640
rect 92200 48640 92360 48800
rect 92200 48800 92360 48960
rect 92200 48960 92360 49120
rect 92200 49120 92360 49280
rect 92200 49280 92360 49440
rect 92200 49440 92360 49600
rect 92200 49600 92360 49760
rect 92200 49760 92360 49920
rect 92200 49920 92360 50080
rect 92200 50080 92360 50240
rect 92200 50240 92360 50400
rect 92200 50400 92360 50560
rect 92200 50560 92360 50720
rect 92200 50720 92360 50880
rect 92200 50880 92360 51040
rect 92200 51040 92360 51200
rect 92200 51200 92360 51360
rect 92200 51360 92360 51520
rect 92200 51520 92360 51680
rect 92200 51680 92360 51840
rect 92200 51840 92360 52000
rect 92360 38560 92520 38720
rect 92360 38720 92520 38880
rect 92360 38880 92520 39040
rect 92360 39040 92520 39200
rect 92360 39200 92520 39360
rect 92360 39360 92520 39520
rect 92360 39520 92520 39680
rect 92360 39680 92520 39840
rect 92360 39840 92520 40000
rect 92360 40000 92520 40160
rect 92360 40160 92520 40320
rect 92360 40320 92520 40480
rect 92360 40480 92520 40640
rect 92360 40640 92520 40800
rect 92360 40800 92520 40960
rect 92360 40960 92520 41120
rect 92360 41120 92520 41280
rect 92360 41280 92520 41440
rect 92360 41440 92520 41600
rect 92360 41600 92520 41760
rect 92360 41760 92520 41920
rect 92360 41920 92520 42080
rect 92360 42080 92520 42240
rect 92360 42240 92520 42400
rect 92360 42400 92520 42560
rect 92360 42560 92520 42720
rect 92360 42720 92520 42880
rect 92360 42880 92520 43040
rect 92360 43040 92520 43200
rect 92360 43200 92520 43360
rect 92360 43360 92520 43520
rect 92360 43520 92520 43680
rect 92360 43680 92520 43840
rect 92360 43840 92520 44000
rect 92360 44000 92520 44160
rect 92360 44160 92520 44320
rect 92360 44320 92520 44480
rect 92360 44480 92520 44640
rect 92360 44640 92520 44800
rect 92360 44800 92520 44960
rect 92360 44960 92520 45120
rect 92360 45120 92520 45280
rect 92360 45280 92520 45440
rect 92360 45440 92520 45600
rect 92360 45600 92520 45760
rect 92360 45760 92520 45920
rect 92360 45920 92520 46080
rect 92360 46080 92520 46240
rect 92360 46240 92520 46400
rect 92360 46400 92520 46560
rect 92360 46560 92520 46720
rect 92360 46720 92520 46880
rect 92360 46880 92520 47040
rect 92360 47040 92520 47200
rect 92360 47200 92520 47360
rect 92360 47360 92520 47520
rect 92360 47520 92520 47680
rect 92360 47680 92520 47840
rect 92360 47840 92520 48000
rect 92360 48000 92520 48160
rect 92360 48160 92520 48320
rect 92360 48320 92520 48480
rect 92360 48480 92520 48640
rect 92360 48640 92520 48800
rect 92360 48800 92520 48960
rect 92360 48960 92520 49120
rect 92360 49120 92520 49280
rect 92360 49280 92520 49440
rect 92360 49440 92520 49600
rect 92360 49600 92520 49760
rect 92360 49760 92520 49920
rect 92360 49920 92520 50080
rect 92360 50080 92520 50240
rect 92360 50240 92520 50400
rect 92360 50400 92520 50560
rect 92360 50560 92520 50720
rect 92360 50720 92520 50880
rect 92360 50880 92520 51040
rect 92360 51040 92520 51200
rect 92360 51200 92520 51360
rect 92360 51360 92520 51520
rect 92360 51520 92520 51680
rect 92360 51680 92520 51840
rect 92520 28320 92680 28480
rect 92520 28480 92680 28640
rect 92520 28640 92680 28800
rect 92520 28800 92680 28960
rect 92520 28960 92680 29120
rect 92520 29120 92680 29280
rect 92520 29280 92680 29440
rect 92520 29440 92680 29600
rect 92520 29600 92680 29760
rect 92520 29760 92680 29920
rect 92520 29920 92680 30080
rect 92520 38080 92680 38240
rect 92520 38240 92680 38400
rect 92520 38400 92680 38560
rect 92520 38560 92680 38720
rect 92520 38720 92680 38880
rect 92520 38880 92680 39040
rect 92520 39040 92680 39200
rect 92520 39200 92680 39360
rect 92520 39360 92680 39520
rect 92520 39520 92680 39680
rect 92520 39680 92680 39840
rect 92520 39840 92680 40000
rect 92520 40000 92680 40160
rect 92520 40160 92680 40320
rect 92520 40320 92680 40480
rect 92520 40480 92680 40640
rect 92520 40640 92680 40800
rect 92520 40800 92680 40960
rect 92520 40960 92680 41120
rect 92520 41120 92680 41280
rect 92520 41280 92680 41440
rect 92520 41440 92680 41600
rect 92520 41600 92680 41760
rect 92520 41760 92680 41920
rect 92520 41920 92680 42080
rect 92520 42080 92680 42240
rect 92520 42240 92680 42400
rect 92520 42400 92680 42560
rect 92520 42560 92680 42720
rect 92520 42720 92680 42880
rect 92520 42880 92680 43040
rect 92520 43040 92680 43200
rect 92520 43200 92680 43360
rect 92520 43360 92680 43520
rect 92520 43520 92680 43680
rect 92520 43680 92680 43840
rect 92520 43840 92680 44000
rect 92520 44000 92680 44160
rect 92520 44160 92680 44320
rect 92520 44320 92680 44480
rect 92520 44480 92680 44640
rect 92520 44640 92680 44800
rect 92520 44800 92680 44960
rect 92520 44960 92680 45120
rect 92520 45120 92680 45280
rect 92520 45280 92680 45440
rect 92520 45440 92680 45600
rect 92520 45600 92680 45760
rect 92520 45760 92680 45920
rect 92520 45920 92680 46080
rect 92520 46080 92680 46240
rect 92520 46240 92680 46400
rect 92520 46400 92680 46560
rect 92520 46560 92680 46720
rect 92520 46720 92680 46880
rect 92520 46880 92680 47040
rect 92520 47040 92680 47200
rect 92520 47200 92680 47360
rect 92520 47360 92680 47520
rect 92520 47520 92680 47680
rect 92520 47680 92680 47840
rect 92520 47840 92680 48000
rect 92520 48000 92680 48160
rect 92520 48160 92680 48320
rect 92520 48320 92680 48480
rect 92520 48480 92680 48640
rect 92520 48640 92680 48800
rect 92520 48800 92680 48960
rect 92520 48960 92680 49120
rect 92520 49120 92680 49280
rect 92520 49280 92680 49440
rect 92520 49440 92680 49600
rect 92520 49600 92680 49760
rect 92520 49760 92680 49920
rect 92520 49920 92680 50080
rect 92520 50080 92680 50240
rect 92520 50240 92680 50400
rect 92520 50400 92680 50560
rect 92520 50560 92680 50720
rect 92520 50720 92680 50880
rect 92520 50880 92680 51040
rect 92520 51040 92680 51200
rect 92520 51200 92680 51360
rect 92520 51360 92680 51520
rect 92520 51520 92680 51680
rect 92520 51680 92680 51840
rect 92680 27680 92840 27840
rect 92680 27840 92840 28000
rect 92680 28000 92840 28160
rect 92680 28160 92840 28320
rect 92680 28320 92840 28480
rect 92680 28480 92840 28640
rect 92680 28640 92840 28800
rect 92680 28800 92840 28960
rect 92680 28960 92840 29120
rect 92680 29120 92840 29280
rect 92680 29280 92840 29440
rect 92680 29440 92840 29600
rect 92680 29600 92840 29760
rect 92680 29760 92840 29920
rect 92680 29920 92840 30080
rect 92680 30080 92840 30240
rect 92680 30240 92840 30400
rect 92680 30400 92840 30560
rect 92680 37600 92840 37760
rect 92680 37760 92840 37920
rect 92680 37920 92840 38080
rect 92680 38080 92840 38240
rect 92680 38240 92840 38400
rect 92680 38400 92840 38560
rect 92680 38560 92840 38720
rect 92680 38720 92840 38880
rect 92680 38880 92840 39040
rect 92680 39040 92840 39200
rect 92680 39200 92840 39360
rect 92680 39360 92840 39520
rect 92680 39520 92840 39680
rect 92680 39680 92840 39840
rect 92680 39840 92840 40000
rect 92680 40000 92840 40160
rect 92680 40160 92840 40320
rect 92680 40320 92840 40480
rect 92680 40480 92840 40640
rect 92680 40640 92840 40800
rect 92680 40800 92840 40960
rect 92680 40960 92840 41120
rect 92680 41120 92840 41280
rect 92680 41280 92840 41440
rect 92680 41440 92840 41600
rect 92680 41600 92840 41760
rect 92680 41760 92840 41920
rect 92680 41920 92840 42080
rect 92680 42080 92840 42240
rect 92680 42240 92840 42400
rect 92680 42400 92840 42560
rect 92680 42560 92840 42720
rect 92680 42720 92840 42880
rect 92680 42880 92840 43040
rect 92680 43040 92840 43200
rect 92680 43200 92840 43360
rect 92680 43360 92840 43520
rect 92680 43520 92840 43680
rect 92680 43680 92840 43840
rect 92680 43840 92840 44000
rect 92680 44000 92840 44160
rect 92680 44160 92840 44320
rect 92680 44320 92840 44480
rect 92680 44480 92840 44640
rect 92680 44640 92840 44800
rect 92680 44800 92840 44960
rect 92680 44960 92840 45120
rect 92680 45120 92840 45280
rect 92680 45280 92840 45440
rect 92680 45440 92840 45600
rect 92680 45600 92840 45760
rect 92680 45760 92840 45920
rect 92680 45920 92840 46080
rect 92680 46080 92840 46240
rect 92680 46240 92840 46400
rect 92680 46400 92840 46560
rect 92680 46560 92840 46720
rect 92680 46720 92840 46880
rect 92680 46880 92840 47040
rect 92680 47040 92840 47200
rect 92680 47200 92840 47360
rect 92680 47360 92840 47520
rect 92680 47520 92840 47680
rect 92680 47680 92840 47840
rect 92680 47840 92840 48000
rect 92680 48000 92840 48160
rect 92680 48160 92840 48320
rect 92680 48320 92840 48480
rect 92680 48480 92840 48640
rect 92680 48640 92840 48800
rect 92680 48800 92840 48960
rect 92680 48960 92840 49120
rect 92680 49120 92840 49280
rect 92680 49280 92840 49440
rect 92680 49440 92840 49600
rect 92680 49600 92840 49760
rect 92680 49760 92840 49920
rect 92680 49920 92840 50080
rect 92680 50080 92840 50240
rect 92680 50240 92840 50400
rect 92680 50400 92840 50560
rect 92680 50560 92840 50720
rect 92680 50720 92840 50880
rect 92680 50880 92840 51040
rect 92680 51040 92840 51200
rect 92680 51200 92840 51360
rect 92680 51360 92840 51520
rect 92680 51520 92840 51680
rect 92840 27360 93000 27520
rect 92840 27520 93000 27680
rect 92840 27680 93000 27840
rect 92840 27840 93000 28000
rect 92840 28000 93000 28160
rect 92840 28160 93000 28320
rect 92840 28320 93000 28480
rect 92840 28480 93000 28640
rect 92840 28640 93000 28800
rect 92840 28800 93000 28960
rect 92840 28960 93000 29120
rect 92840 29120 93000 29280
rect 92840 29280 93000 29440
rect 92840 29440 93000 29600
rect 92840 29600 93000 29760
rect 92840 29760 93000 29920
rect 92840 29920 93000 30080
rect 92840 30080 93000 30240
rect 92840 30240 93000 30400
rect 92840 30400 93000 30560
rect 92840 30560 93000 30720
rect 92840 30720 93000 30880
rect 92840 30880 93000 31040
rect 92840 37120 93000 37280
rect 92840 37280 93000 37440
rect 92840 37440 93000 37600
rect 92840 37600 93000 37760
rect 92840 37760 93000 37920
rect 92840 37920 93000 38080
rect 92840 38080 93000 38240
rect 92840 38240 93000 38400
rect 92840 38400 93000 38560
rect 92840 38560 93000 38720
rect 92840 38720 93000 38880
rect 92840 38880 93000 39040
rect 92840 39040 93000 39200
rect 92840 39200 93000 39360
rect 92840 39360 93000 39520
rect 92840 39520 93000 39680
rect 92840 39680 93000 39840
rect 92840 39840 93000 40000
rect 92840 40000 93000 40160
rect 92840 40160 93000 40320
rect 92840 40320 93000 40480
rect 92840 40480 93000 40640
rect 92840 40640 93000 40800
rect 92840 40800 93000 40960
rect 92840 40960 93000 41120
rect 92840 41120 93000 41280
rect 92840 41280 93000 41440
rect 92840 41440 93000 41600
rect 92840 41600 93000 41760
rect 92840 41760 93000 41920
rect 92840 41920 93000 42080
rect 92840 42080 93000 42240
rect 92840 42240 93000 42400
rect 92840 42400 93000 42560
rect 92840 42560 93000 42720
rect 92840 42720 93000 42880
rect 92840 42880 93000 43040
rect 92840 43040 93000 43200
rect 92840 43200 93000 43360
rect 92840 43360 93000 43520
rect 92840 43520 93000 43680
rect 92840 43680 93000 43840
rect 92840 43840 93000 44000
rect 92840 44000 93000 44160
rect 92840 44160 93000 44320
rect 92840 44320 93000 44480
rect 92840 44480 93000 44640
rect 92840 44640 93000 44800
rect 92840 44800 93000 44960
rect 92840 44960 93000 45120
rect 92840 45120 93000 45280
rect 92840 45280 93000 45440
rect 92840 45440 93000 45600
rect 92840 45600 93000 45760
rect 92840 45760 93000 45920
rect 92840 45920 93000 46080
rect 92840 46080 93000 46240
rect 92840 46240 93000 46400
rect 92840 46400 93000 46560
rect 92840 46560 93000 46720
rect 92840 46720 93000 46880
rect 92840 46880 93000 47040
rect 92840 47040 93000 47200
rect 92840 47200 93000 47360
rect 92840 47360 93000 47520
rect 92840 47520 93000 47680
rect 92840 47680 93000 47840
rect 92840 47840 93000 48000
rect 92840 48000 93000 48160
rect 92840 48160 93000 48320
rect 92840 48320 93000 48480
rect 92840 48480 93000 48640
rect 92840 48640 93000 48800
rect 92840 48800 93000 48960
rect 92840 48960 93000 49120
rect 92840 49120 93000 49280
rect 92840 49280 93000 49440
rect 92840 49440 93000 49600
rect 92840 49600 93000 49760
rect 92840 49760 93000 49920
rect 92840 49920 93000 50080
rect 92840 50080 93000 50240
rect 92840 50240 93000 50400
rect 92840 50400 93000 50560
rect 92840 50560 93000 50720
rect 92840 50720 93000 50880
rect 92840 50880 93000 51040
rect 92840 51040 93000 51200
rect 92840 51200 93000 51360
rect 92840 51360 93000 51520
rect 93000 27040 93160 27200
rect 93000 27200 93160 27360
rect 93000 27360 93160 27520
rect 93000 27520 93160 27680
rect 93000 27680 93160 27840
rect 93000 27840 93160 28000
rect 93000 28000 93160 28160
rect 93000 28160 93160 28320
rect 93000 28320 93160 28480
rect 93000 28480 93160 28640
rect 93000 28640 93160 28800
rect 93000 28800 93160 28960
rect 93000 28960 93160 29120
rect 93000 29120 93160 29280
rect 93000 29280 93160 29440
rect 93000 29440 93160 29600
rect 93000 29600 93160 29760
rect 93000 29760 93160 29920
rect 93000 29920 93160 30080
rect 93000 30080 93160 30240
rect 93000 30240 93160 30400
rect 93000 30400 93160 30560
rect 93000 30560 93160 30720
rect 93000 30720 93160 30880
rect 93000 30880 93160 31040
rect 93000 31040 93160 31200
rect 93000 31200 93160 31360
rect 93000 36640 93160 36800
rect 93000 36800 93160 36960
rect 93000 36960 93160 37120
rect 93000 37120 93160 37280
rect 93000 37280 93160 37440
rect 93000 37440 93160 37600
rect 93000 37600 93160 37760
rect 93000 37760 93160 37920
rect 93000 37920 93160 38080
rect 93000 38080 93160 38240
rect 93000 38240 93160 38400
rect 93000 38400 93160 38560
rect 93000 38560 93160 38720
rect 93000 38720 93160 38880
rect 93000 38880 93160 39040
rect 93000 39040 93160 39200
rect 93000 39200 93160 39360
rect 93000 39360 93160 39520
rect 93000 39520 93160 39680
rect 93000 39680 93160 39840
rect 93000 39840 93160 40000
rect 93000 40000 93160 40160
rect 93000 40160 93160 40320
rect 93000 40320 93160 40480
rect 93000 40480 93160 40640
rect 93000 40640 93160 40800
rect 93000 40800 93160 40960
rect 93000 40960 93160 41120
rect 93000 41120 93160 41280
rect 93000 41280 93160 41440
rect 93000 41440 93160 41600
rect 93000 41600 93160 41760
rect 93000 41760 93160 41920
rect 93000 41920 93160 42080
rect 93000 42080 93160 42240
rect 93000 42240 93160 42400
rect 93000 42400 93160 42560
rect 93000 42560 93160 42720
rect 93000 42720 93160 42880
rect 93000 42880 93160 43040
rect 93000 43040 93160 43200
rect 93000 43200 93160 43360
rect 93000 43360 93160 43520
rect 93000 43520 93160 43680
rect 93000 43680 93160 43840
rect 93000 43840 93160 44000
rect 93000 44000 93160 44160
rect 93000 44160 93160 44320
rect 93000 44320 93160 44480
rect 93000 44480 93160 44640
rect 93000 44640 93160 44800
rect 93000 44800 93160 44960
rect 93000 44960 93160 45120
rect 93000 45120 93160 45280
rect 93000 45280 93160 45440
rect 93000 45440 93160 45600
rect 93000 45600 93160 45760
rect 93000 45760 93160 45920
rect 93000 45920 93160 46080
rect 93000 46080 93160 46240
rect 93000 46240 93160 46400
rect 93000 46400 93160 46560
rect 93000 46560 93160 46720
rect 93000 46720 93160 46880
rect 93000 46880 93160 47040
rect 93000 47040 93160 47200
rect 93000 47200 93160 47360
rect 93000 47360 93160 47520
rect 93000 47520 93160 47680
rect 93000 47680 93160 47840
rect 93000 47840 93160 48000
rect 93000 48000 93160 48160
rect 93000 48160 93160 48320
rect 93000 48320 93160 48480
rect 93000 48480 93160 48640
rect 93000 48640 93160 48800
rect 93000 48800 93160 48960
rect 93000 48960 93160 49120
rect 93000 49120 93160 49280
rect 93000 49280 93160 49440
rect 93000 49440 93160 49600
rect 93000 49600 93160 49760
rect 93000 49760 93160 49920
rect 93000 49920 93160 50080
rect 93000 50080 93160 50240
rect 93000 50240 93160 50400
rect 93000 50400 93160 50560
rect 93000 50560 93160 50720
rect 93000 50720 93160 50880
rect 93000 50880 93160 51040
rect 93000 51040 93160 51200
rect 93000 51200 93160 51360
rect 93160 26880 93320 27040
rect 93160 27040 93320 27200
rect 93160 27200 93320 27360
rect 93160 27360 93320 27520
rect 93160 27520 93320 27680
rect 93160 27680 93320 27840
rect 93160 27840 93320 28000
rect 93160 28000 93320 28160
rect 93160 28160 93320 28320
rect 93160 28320 93320 28480
rect 93160 28480 93320 28640
rect 93160 28640 93320 28800
rect 93160 28800 93320 28960
rect 93160 28960 93320 29120
rect 93160 29120 93320 29280
rect 93160 29280 93320 29440
rect 93160 29440 93320 29600
rect 93160 29600 93320 29760
rect 93160 29760 93320 29920
rect 93160 29920 93320 30080
rect 93160 30080 93320 30240
rect 93160 30240 93320 30400
rect 93160 30400 93320 30560
rect 93160 30560 93320 30720
rect 93160 30720 93320 30880
rect 93160 30880 93320 31040
rect 93160 31040 93320 31200
rect 93160 31200 93320 31360
rect 93160 31360 93320 31520
rect 93160 36000 93320 36160
rect 93160 36160 93320 36320
rect 93160 36320 93320 36480
rect 93160 36480 93320 36640
rect 93160 36640 93320 36800
rect 93160 36800 93320 36960
rect 93160 36960 93320 37120
rect 93160 37120 93320 37280
rect 93160 37280 93320 37440
rect 93160 37440 93320 37600
rect 93160 37600 93320 37760
rect 93160 37760 93320 37920
rect 93160 37920 93320 38080
rect 93160 38080 93320 38240
rect 93160 38240 93320 38400
rect 93160 38400 93320 38560
rect 93160 38560 93320 38720
rect 93160 38720 93320 38880
rect 93160 38880 93320 39040
rect 93160 39040 93320 39200
rect 93160 39200 93320 39360
rect 93160 39360 93320 39520
rect 93160 39520 93320 39680
rect 93160 39680 93320 39840
rect 93160 39840 93320 40000
rect 93160 40000 93320 40160
rect 93160 40160 93320 40320
rect 93160 40320 93320 40480
rect 93160 40480 93320 40640
rect 93160 40640 93320 40800
rect 93160 40800 93320 40960
rect 93160 40960 93320 41120
rect 93160 41120 93320 41280
rect 93160 41280 93320 41440
rect 93160 41440 93320 41600
rect 93160 41600 93320 41760
rect 93160 41760 93320 41920
rect 93160 41920 93320 42080
rect 93160 42080 93320 42240
rect 93160 42240 93320 42400
rect 93160 42400 93320 42560
rect 93160 42560 93320 42720
rect 93160 42720 93320 42880
rect 93160 42880 93320 43040
rect 93160 43040 93320 43200
rect 93160 43200 93320 43360
rect 93160 43360 93320 43520
rect 93160 43520 93320 43680
rect 93160 43680 93320 43840
rect 93160 43840 93320 44000
rect 93160 44000 93320 44160
rect 93160 44160 93320 44320
rect 93160 44320 93320 44480
rect 93160 44480 93320 44640
rect 93160 44640 93320 44800
rect 93160 44800 93320 44960
rect 93160 44960 93320 45120
rect 93160 45120 93320 45280
rect 93160 45280 93320 45440
rect 93160 45440 93320 45600
rect 93160 45600 93320 45760
rect 93160 45760 93320 45920
rect 93160 45920 93320 46080
rect 93160 46080 93320 46240
rect 93160 46240 93320 46400
rect 93160 46400 93320 46560
rect 93160 46560 93320 46720
rect 93160 46720 93320 46880
rect 93160 46880 93320 47040
rect 93160 47040 93320 47200
rect 93160 47200 93320 47360
rect 93160 47360 93320 47520
rect 93160 47520 93320 47680
rect 93160 47680 93320 47840
rect 93160 47840 93320 48000
rect 93160 48000 93320 48160
rect 93160 48160 93320 48320
rect 93160 48320 93320 48480
rect 93160 48480 93320 48640
rect 93160 48640 93320 48800
rect 93160 48800 93320 48960
rect 93160 48960 93320 49120
rect 93160 49120 93320 49280
rect 93160 49280 93320 49440
rect 93160 49440 93320 49600
rect 93160 49600 93320 49760
rect 93160 49760 93320 49920
rect 93160 49920 93320 50080
rect 93160 50080 93320 50240
rect 93160 50240 93320 50400
rect 93160 50400 93320 50560
rect 93160 50560 93320 50720
rect 93160 50720 93320 50880
rect 93160 50880 93320 51040
rect 93160 51040 93320 51200
rect 93320 26560 93480 26720
rect 93320 26720 93480 26880
rect 93320 26880 93480 27040
rect 93320 27040 93480 27200
rect 93320 27200 93480 27360
rect 93320 27360 93480 27520
rect 93320 27520 93480 27680
rect 93320 27680 93480 27840
rect 93320 27840 93480 28000
rect 93320 28000 93480 28160
rect 93320 28160 93480 28320
rect 93320 28320 93480 28480
rect 93320 28480 93480 28640
rect 93320 28640 93480 28800
rect 93320 28800 93480 28960
rect 93320 28960 93480 29120
rect 93320 29120 93480 29280
rect 93320 29280 93480 29440
rect 93320 29440 93480 29600
rect 93320 29600 93480 29760
rect 93320 29760 93480 29920
rect 93320 29920 93480 30080
rect 93320 30080 93480 30240
rect 93320 30240 93480 30400
rect 93320 30400 93480 30560
rect 93320 30560 93480 30720
rect 93320 30720 93480 30880
rect 93320 30880 93480 31040
rect 93320 31040 93480 31200
rect 93320 31200 93480 31360
rect 93320 31360 93480 31520
rect 93320 31520 93480 31680
rect 93320 35520 93480 35680
rect 93320 35680 93480 35840
rect 93320 35840 93480 36000
rect 93320 36000 93480 36160
rect 93320 36160 93480 36320
rect 93320 36320 93480 36480
rect 93320 36480 93480 36640
rect 93320 36640 93480 36800
rect 93320 36800 93480 36960
rect 93320 36960 93480 37120
rect 93320 37120 93480 37280
rect 93320 37280 93480 37440
rect 93320 37440 93480 37600
rect 93320 37600 93480 37760
rect 93320 37760 93480 37920
rect 93320 37920 93480 38080
rect 93320 38080 93480 38240
rect 93320 38240 93480 38400
rect 93320 38400 93480 38560
rect 93320 38560 93480 38720
rect 93320 38720 93480 38880
rect 93320 38880 93480 39040
rect 93320 39040 93480 39200
rect 93320 39200 93480 39360
rect 93320 39360 93480 39520
rect 93320 39520 93480 39680
rect 93320 39680 93480 39840
rect 93320 39840 93480 40000
rect 93320 40000 93480 40160
rect 93320 40160 93480 40320
rect 93320 40320 93480 40480
rect 93320 40480 93480 40640
rect 93320 40640 93480 40800
rect 93320 40800 93480 40960
rect 93320 40960 93480 41120
rect 93320 41120 93480 41280
rect 93320 41280 93480 41440
rect 93320 41440 93480 41600
rect 93320 41600 93480 41760
rect 93320 41760 93480 41920
rect 93320 41920 93480 42080
rect 93320 42080 93480 42240
rect 93320 42240 93480 42400
rect 93320 42400 93480 42560
rect 93320 42560 93480 42720
rect 93320 42720 93480 42880
rect 93320 42880 93480 43040
rect 93320 43040 93480 43200
rect 93320 43200 93480 43360
rect 93320 43360 93480 43520
rect 93320 43520 93480 43680
rect 93320 43680 93480 43840
rect 93320 43840 93480 44000
rect 93320 45920 93480 46080
rect 93320 46080 93480 46240
rect 93320 46240 93480 46400
rect 93320 46400 93480 46560
rect 93320 46560 93480 46720
rect 93320 46720 93480 46880
rect 93320 46880 93480 47040
rect 93320 47040 93480 47200
rect 93320 47200 93480 47360
rect 93320 47360 93480 47520
rect 93320 47520 93480 47680
rect 93320 47680 93480 47840
rect 93320 47840 93480 48000
rect 93320 48000 93480 48160
rect 93320 48160 93480 48320
rect 93320 48320 93480 48480
rect 93320 48480 93480 48640
rect 93320 48640 93480 48800
rect 93320 48800 93480 48960
rect 93320 48960 93480 49120
rect 93320 49120 93480 49280
rect 93320 49280 93480 49440
rect 93320 49440 93480 49600
rect 93320 49600 93480 49760
rect 93320 49760 93480 49920
rect 93320 49920 93480 50080
rect 93320 50080 93480 50240
rect 93320 50240 93480 50400
rect 93320 50400 93480 50560
rect 93320 50560 93480 50720
rect 93320 50720 93480 50880
rect 93320 50880 93480 51040
rect 93480 26400 93640 26560
rect 93480 26560 93640 26720
rect 93480 26720 93640 26880
rect 93480 26880 93640 27040
rect 93480 27040 93640 27200
rect 93480 27200 93640 27360
rect 93480 27360 93640 27520
rect 93480 27520 93640 27680
rect 93480 27680 93640 27840
rect 93480 27840 93640 28000
rect 93480 28000 93640 28160
rect 93480 28160 93640 28320
rect 93480 28320 93640 28480
rect 93480 28480 93640 28640
rect 93480 28640 93640 28800
rect 93480 28800 93640 28960
rect 93480 28960 93640 29120
rect 93480 29120 93640 29280
rect 93480 29280 93640 29440
rect 93480 29440 93640 29600
rect 93480 29600 93640 29760
rect 93480 29760 93640 29920
rect 93480 29920 93640 30080
rect 93480 30080 93640 30240
rect 93480 30240 93640 30400
rect 93480 30400 93640 30560
rect 93480 30560 93640 30720
rect 93480 30720 93640 30880
rect 93480 30880 93640 31040
rect 93480 31040 93640 31200
rect 93480 31200 93640 31360
rect 93480 31360 93640 31520
rect 93480 31520 93640 31680
rect 93480 31680 93640 31840
rect 93480 31840 93640 32000
rect 93480 35040 93640 35200
rect 93480 35200 93640 35360
rect 93480 35360 93640 35520
rect 93480 35520 93640 35680
rect 93480 35680 93640 35840
rect 93480 35840 93640 36000
rect 93480 36000 93640 36160
rect 93480 36160 93640 36320
rect 93480 36320 93640 36480
rect 93480 36480 93640 36640
rect 93480 36640 93640 36800
rect 93480 36800 93640 36960
rect 93480 36960 93640 37120
rect 93480 37120 93640 37280
rect 93480 37280 93640 37440
rect 93480 37440 93640 37600
rect 93480 37600 93640 37760
rect 93480 37760 93640 37920
rect 93480 37920 93640 38080
rect 93480 38080 93640 38240
rect 93480 38240 93640 38400
rect 93480 38400 93640 38560
rect 93480 38560 93640 38720
rect 93480 38720 93640 38880
rect 93480 38880 93640 39040
rect 93480 39040 93640 39200
rect 93480 39200 93640 39360
rect 93480 39360 93640 39520
rect 93480 39520 93640 39680
rect 93480 39680 93640 39840
rect 93480 39840 93640 40000
rect 93480 40000 93640 40160
rect 93480 40160 93640 40320
rect 93480 40320 93640 40480
rect 93480 40480 93640 40640
rect 93480 40640 93640 40800
rect 93480 40800 93640 40960
rect 93480 40960 93640 41120
rect 93480 41120 93640 41280
rect 93480 41280 93640 41440
rect 93480 41440 93640 41600
rect 93480 41600 93640 41760
rect 93480 41760 93640 41920
rect 93480 41920 93640 42080
rect 93480 42080 93640 42240
rect 93480 42240 93640 42400
rect 93480 42400 93640 42560
rect 93480 42560 93640 42720
rect 93480 42720 93640 42880
rect 93480 42880 93640 43040
rect 93480 43040 93640 43200
rect 93480 43200 93640 43360
rect 93480 46400 93640 46560
rect 93480 46560 93640 46720
rect 93480 46720 93640 46880
rect 93480 46880 93640 47040
rect 93480 47040 93640 47200
rect 93480 47200 93640 47360
rect 93480 47360 93640 47520
rect 93480 47520 93640 47680
rect 93480 47680 93640 47840
rect 93480 47840 93640 48000
rect 93480 48000 93640 48160
rect 93480 48160 93640 48320
rect 93480 48320 93640 48480
rect 93480 48480 93640 48640
rect 93480 48640 93640 48800
rect 93480 48800 93640 48960
rect 93480 48960 93640 49120
rect 93480 49120 93640 49280
rect 93480 49280 93640 49440
rect 93480 49440 93640 49600
rect 93480 49600 93640 49760
rect 93480 49760 93640 49920
rect 93480 49920 93640 50080
rect 93480 50080 93640 50240
rect 93480 50240 93640 50400
rect 93480 50400 93640 50560
rect 93480 50560 93640 50720
rect 93480 50720 93640 50880
rect 93640 26240 93800 26400
rect 93640 26400 93800 26560
rect 93640 26560 93800 26720
rect 93640 26720 93800 26880
rect 93640 26880 93800 27040
rect 93640 27040 93800 27200
rect 93640 27200 93800 27360
rect 93640 27360 93800 27520
rect 93640 27520 93800 27680
rect 93640 27680 93800 27840
rect 93640 27840 93800 28000
rect 93640 28000 93800 28160
rect 93640 28160 93800 28320
rect 93640 28320 93800 28480
rect 93640 28480 93800 28640
rect 93640 28640 93800 28800
rect 93640 28800 93800 28960
rect 93640 28960 93800 29120
rect 93640 29120 93800 29280
rect 93640 29280 93800 29440
rect 93640 29440 93800 29600
rect 93640 29600 93800 29760
rect 93640 29760 93800 29920
rect 93640 29920 93800 30080
rect 93640 30080 93800 30240
rect 93640 30240 93800 30400
rect 93640 30400 93800 30560
rect 93640 30560 93800 30720
rect 93640 30720 93800 30880
rect 93640 30880 93800 31040
rect 93640 31040 93800 31200
rect 93640 31200 93800 31360
rect 93640 31360 93800 31520
rect 93640 31520 93800 31680
rect 93640 31680 93800 31840
rect 93640 31840 93800 32000
rect 93640 32000 93800 32160
rect 93640 32160 93800 32320
rect 93640 34240 93800 34400
rect 93640 34400 93800 34560
rect 93640 34560 93800 34720
rect 93640 34720 93800 34880
rect 93640 34880 93800 35040
rect 93640 35040 93800 35200
rect 93640 35200 93800 35360
rect 93640 35360 93800 35520
rect 93640 35520 93800 35680
rect 93640 35680 93800 35840
rect 93640 35840 93800 36000
rect 93640 36000 93800 36160
rect 93640 36160 93800 36320
rect 93640 36320 93800 36480
rect 93640 36480 93800 36640
rect 93640 36640 93800 36800
rect 93640 36800 93800 36960
rect 93640 36960 93800 37120
rect 93640 37120 93800 37280
rect 93640 37280 93800 37440
rect 93640 37440 93800 37600
rect 93640 37600 93800 37760
rect 93640 37760 93800 37920
rect 93640 37920 93800 38080
rect 93640 38080 93800 38240
rect 93640 38240 93800 38400
rect 93640 38400 93800 38560
rect 93640 38560 93800 38720
rect 93640 38720 93800 38880
rect 93640 38880 93800 39040
rect 93640 39040 93800 39200
rect 93640 39200 93800 39360
rect 93640 39360 93800 39520
rect 93640 39520 93800 39680
rect 93640 39680 93800 39840
rect 93640 39840 93800 40000
rect 93640 40000 93800 40160
rect 93640 40160 93800 40320
rect 93640 40320 93800 40480
rect 93640 40480 93800 40640
rect 93640 40640 93800 40800
rect 93640 40800 93800 40960
rect 93640 40960 93800 41120
rect 93640 41120 93800 41280
rect 93640 41280 93800 41440
rect 93640 41440 93800 41600
rect 93640 41600 93800 41760
rect 93640 41760 93800 41920
rect 93640 41920 93800 42080
rect 93640 42080 93800 42240
rect 93640 42240 93800 42400
rect 93640 42400 93800 42560
rect 93640 42560 93800 42720
rect 93640 42720 93800 42880
rect 93640 46720 93800 46880
rect 93640 46880 93800 47040
rect 93640 47040 93800 47200
rect 93640 47200 93800 47360
rect 93640 47360 93800 47520
rect 93640 47520 93800 47680
rect 93640 47680 93800 47840
rect 93640 47840 93800 48000
rect 93640 48000 93800 48160
rect 93640 48160 93800 48320
rect 93640 48320 93800 48480
rect 93640 48480 93800 48640
rect 93640 48640 93800 48800
rect 93640 48800 93800 48960
rect 93640 48960 93800 49120
rect 93640 49120 93800 49280
rect 93640 49280 93800 49440
rect 93640 49440 93800 49600
rect 93640 49600 93800 49760
rect 93640 49760 93800 49920
rect 93640 49920 93800 50080
rect 93640 50080 93800 50240
rect 93640 50240 93800 50400
rect 93640 50400 93800 50560
rect 93800 26080 93960 26240
rect 93800 26240 93960 26400
rect 93800 26400 93960 26560
rect 93800 26560 93960 26720
rect 93800 26720 93960 26880
rect 93800 26880 93960 27040
rect 93800 27040 93960 27200
rect 93800 27200 93960 27360
rect 93800 27360 93960 27520
rect 93800 27520 93960 27680
rect 93800 27680 93960 27840
rect 93800 27840 93960 28000
rect 93800 28000 93960 28160
rect 93800 28160 93960 28320
rect 93800 28320 93960 28480
rect 93800 28480 93960 28640
rect 93800 28640 93960 28800
rect 93800 28800 93960 28960
rect 93800 28960 93960 29120
rect 93800 29120 93960 29280
rect 93800 29280 93960 29440
rect 93800 29440 93960 29600
rect 93800 29600 93960 29760
rect 93800 29760 93960 29920
rect 93800 29920 93960 30080
rect 93800 30080 93960 30240
rect 93800 30240 93960 30400
rect 93800 30400 93960 30560
rect 93800 30560 93960 30720
rect 93800 30720 93960 30880
rect 93800 30880 93960 31040
rect 93800 31040 93960 31200
rect 93800 31200 93960 31360
rect 93800 31360 93960 31520
rect 93800 31520 93960 31680
rect 93800 31680 93960 31840
rect 93800 31840 93960 32000
rect 93800 32000 93960 32160
rect 93800 32160 93960 32320
rect 93800 32320 93960 32480
rect 93800 32480 93960 32640
rect 93800 32640 93960 32800
rect 93800 32800 93960 32960
rect 93800 32960 93960 33120
rect 93800 33120 93960 33280
rect 93800 33280 93960 33440
rect 93800 33440 93960 33600
rect 93800 33600 93960 33760
rect 93800 33760 93960 33920
rect 93800 33920 93960 34080
rect 93800 34080 93960 34240
rect 93800 34240 93960 34400
rect 93800 34400 93960 34560
rect 93800 34560 93960 34720
rect 93800 34720 93960 34880
rect 93800 34880 93960 35040
rect 93800 35040 93960 35200
rect 93800 35200 93960 35360
rect 93800 35360 93960 35520
rect 93800 35520 93960 35680
rect 93800 35680 93960 35840
rect 93800 35840 93960 36000
rect 93800 36000 93960 36160
rect 93800 36160 93960 36320
rect 93800 36320 93960 36480
rect 93800 36480 93960 36640
rect 93800 36640 93960 36800
rect 93800 36800 93960 36960
rect 93800 36960 93960 37120
rect 93800 37120 93960 37280
rect 93800 37280 93960 37440
rect 93800 37440 93960 37600
rect 93800 37600 93960 37760
rect 93800 37760 93960 37920
rect 93800 37920 93960 38080
rect 93800 38080 93960 38240
rect 93800 38240 93960 38400
rect 93800 38400 93960 38560
rect 93800 38560 93960 38720
rect 93800 38720 93960 38880
rect 93800 38880 93960 39040
rect 93800 39040 93960 39200
rect 93800 39200 93960 39360
rect 93800 39360 93960 39520
rect 93800 39520 93960 39680
rect 93800 39680 93960 39840
rect 93800 39840 93960 40000
rect 93800 40000 93960 40160
rect 93800 40160 93960 40320
rect 93800 40320 93960 40480
rect 93800 40480 93960 40640
rect 93800 40640 93960 40800
rect 93800 40800 93960 40960
rect 93800 40960 93960 41120
rect 93800 41120 93960 41280
rect 93800 41280 93960 41440
rect 93800 41440 93960 41600
rect 93800 41600 93960 41760
rect 93800 41760 93960 41920
rect 93800 41920 93960 42080
rect 93800 42080 93960 42240
rect 93800 47040 93960 47200
rect 93800 47200 93960 47360
rect 93800 47360 93960 47520
rect 93800 47520 93960 47680
rect 93800 47680 93960 47840
rect 93800 47840 93960 48000
rect 93800 48000 93960 48160
rect 93800 48160 93960 48320
rect 93800 48320 93960 48480
rect 93800 48480 93960 48640
rect 93800 48640 93960 48800
rect 93800 48800 93960 48960
rect 93800 48960 93960 49120
rect 93800 49120 93960 49280
rect 93800 49280 93960 49440
rect 93800 49440 93960 49600
rect 93800 49600 93960 49760
rect 93800 49760 93960 49920
rect 93800 49920 93960 50080
rect 93800 50080 93960 50240
rect 93960 25920 94120 26080
rect 93960 26080 94120 26240
rect 93960 26240 94120 26400
rect 93960 26400 94120 26560
rect 93960 26560 94120 26720
rect 93960 26720 94120 26880
rect 93960 26880 94120 27040
rect 93960 27040 94120 27200
rect 93960 27200 94120 27360
rect 93960 27360 94120 27520
rect 93960 27520 94120 27680
rect 93960 27680 94120 27840
rect 93960 27840 94120 28000
rect 93960 28000 94120 28160
rect 93960 28160 94120 28320
rect 93960 28320 94120 28480
rect 93960 28480 94120 28640
rect 93960 28640 94120 28800
rect 93960 28800 94120 28960
rect 93960 28960 94120 29120
rect 93960 29120 94120 29280
rect 93960 29280 94120 29440
rect 93960 29440 94120 29600
rect 93960 29600 94120 29760
rect 93960 29760 94120 29920
rect 93960 29920 94120 30080
rect 93960 30080 94120 30240
rect 93960 30240 94120 30400
rect 93960 30400 94120 30560
rect 93960 30560 94120 30720
rect 93960 30720 94120 30880
rect 93960 30880 94120 31040
rect 93960 31040 94120 31200
rect 93960 31200 94120 31360
rect 93960 31360 94120 31520
rect 93960 31520 94120 31680
rect 93960 31680 94120 31840
rect 93960 31840 94120 32000
rect 93960 32000 94120 32160
rect 93960 32160 94120 32320
rect 93960 32320 94120 32480
rect 93960 32480 94120 32640
rect 93960 32640 94120 32800
rect 93960 32800 94120 32960
rect 93960 32960 94120 33120
rect 93960 33120 94120 33280
rect 93960 33280 94120 33440
rect 93960 33440 94120 33600
rect 93960 33600 94120 33760
rect 93960 33760 94120 33920
rect 93960 33920 94120 34080
rect 93960 34080 94120 34240
rect 93960 34240 94120 34400
rect 93960 34400 94120 34560
rect 93960 34560 94120 34720
rect 93960 34720 94120 34880
rect 93960 34880 94120 35040
rect 93960 35040 94120 35200
rect 93960 35200 94120 35360
rect 93960 35360 94120 35520
rect 93960 35520 94120 35680
rect 93960 35680 94120 35840
rect 93960 35840 94120 36000
rect 93960 36000 94120 36160
rect 93960 36160 94120 36320
rect 93960 36320 94120 36480
rect 93960 36480 94120 36640
rect 93960 36640 94120 36800
rect 93960 36800 94120 36960
rect 93960 36960 94120 37120
rect 93960 37120 94120 37280
rect 93960 37280 94120 37440
rect 93960 37440 94120 37600
rect 93960 37600 94120 37760
rect 93960 37760 94120 37920
rect 93960 37920 94120 38080
rect 93960 38080 94120 38240
rect 93960 38240 94120 38400
rect 93960 38400 94120 38560
rect 93960 38560 94120 38720
rect 93960 38720 94120 38880
rect 93960 38880 94120 39040
rect 93960 39040 94120 39200
rect 93960 39200 94120 39360
rect 93960 39360 94120 39520
rect 93960 39520 94120 39680
rect 93960 39680 94120 39840
rect 93960 39840 94120 40000
rect 93960 40000 94120 40160
rect 93960 40160 94120 40320
rect 93960 40320 94120 40480
rect 93960 40480 94120 40640
rect 93960 40640 94120 40800
rect 93960 40800 94120 40960
rect 93960 40960 94120 41120
rect 93960 41120 94120 41280
rect 93960 41280 94120 41440
rect 93960 41440 94120 41600
rect 93960 41600 94120 41760
rect 93960 47360 94120 47520
rect 93960 47520 94120 47680
rect 93960 47680 94120 47840
rect 93960 47840 94120 48000
rect 93960 48000 94120 48160
rect 93960 48160 94120 48320
rect 93960 48320 94120 48480
rect 93960 48480 94120 48640
rect 93960 48640 94120 48800
rect 93960 48800 94120 48960
rect 93960 48960 94120 49120
rect 93960 49120 94120 49280
rect 93960 49280 94120 49440
rect 93960 49440 94120 49600
rect 93960 49600 94120 49760
rect 93960 49760 94120 49920
rect 94120 25760 94280 25920
rect 94120 25920 94280 26080
rect 94120 26080 94280 26240
rect 94120 26240 94280 26400
rect 94120 26400 94280 26560
rect 94120 26560 94280 26720
rect 94120 26720 94280 26880
rect 94120 26880 94280 27040
rect 94120 27040 94280 27200
rect 94120 27200 94280 27360
rect 94120 27360 94280 27520
rect 94120 27520 94280 27680
rect 94120 27680 94280 27840
rect 94120 27840 94280 28000
rect 94120 28000 94280 28160
rect 94120 28160 94280 28320
rect 94120 28320 94280 28480
rect 94120 28480 94280 28640
rect 94120 28640 94280 28800
rect 94120 28800 94280 28960
rect 94120 28960 94280 29120
rect 94120 29120 94280 29280
rect 94120 29280 94280 29440
rect 94120 29440 94280 29600
rect 94120 29600 94280 29760
rect 94120 29760 94280 29920
rect 94120 29920 94280 30080
rect 94120 30080 94280 30240
rect 94120 30240 94280 30400
rect 94120 30400 94280 30560
rect 94120 30560 94280 30720
rect 94120 30720 94280 30880
rect 94120 30880 94280 31040
rect 94120 31040 94280 31200
rect 94120 31200 94280 31360
rect 94120 31360 94280 31520
rect 94120 31520 94280 31680
rect 94120 31680 94280 31840
rect 94120 31840 94280 32000
rect 94120 32000 94280 32160
rect 94120 32160 94280 32320
rect 94120 32320 94280 32480
rect 94120 32480 94280 32640
rect 94120 32640 94280 32800
rect 94120 32800 94280 32960
rect 94120 32960 94280 33120
rect 94120 33120 94280 33280
rect 94120 33280 94280 33440
rect 94120 33440 94280 33600
rect 94120 33600 94280 33760
rect 94120 33760 94280 33920
rect 94120 33920 94280 34080
rect 94120 34080 94280 34240
rect 94120 34240 94280 34400
rect 94120 34400 94280 34560
rect 94120 34560 94280 34720
rect 94120 34720 94280 34880
rect 94120 34880 94280 35040
rect 94120 35040 94280 35200
rect 94120 35200 94280 35360
rect 94120 35360 94280 35520
rect 94120 35520 94280 35680
rect 94120 35680 94280 35840
rect 94120 35840 94280 36000
rect 94120 36000 94280 36160
rect 94120 36160 94280 36320
rect 94120 36320 94280 36480
rect 94120 36480 94280 36640
rect 94120 36640 94280 36800
rect 94120 36800 94280 36960
rect 94120 36960 94280 37120
rect 94120 37120 94280 37280
rect 94120 37280 94280 37440
rect 94120 37440 94280 37600
rect 94120 37600 94280 37760
rect 94120 37760 94280 37920
rect 94120 37920 94280 38080
rect 94120 38080 94280 38240
rect 94120 38240 94280 38400
rect 94120 38400 94280 38560
rect 94120 38560 94280 38720
rect 94120 38720 94280 38880
rect 94120 38880 94280 39040
rect 94120 39040 94280 39200
rect 94120 39200 94280 39360
rect 94120 39360 94280 39520
rect 94120 39520 94280 39680
rect 94120 39680 94280 39840
rect 94120 39840 94280 40000
rect 94120 40000 94280 40160
rect 94120 40160 94280 40320
rect 94120 40320 94280 40480
rect 94120 40480 94280 40640
rect 94120 40640 94280 40800
rect 94120 40800 94280 40960
rect 94120 40960 94280 41120
rect 94120 41120 94280 41280
rect 94120 48160 94280 48320
rect 94120 48320 94280 48480
rect 94120 48480 94280 48640
rect 94120 48640 94280 48800
rect 94120 48800 94280 48960
rect 94120 48960 94280 49120
rect 94120 49120 94280 49280
rect 94280 25760 94440 25920
rect 94280 25920 94440 26080
rect 94280 26080 94440 26240
rect 94280 26240 94440 26400
rect 94280 26400 94440 26560
rect 94280 26560 94440 26720
rect 94280 26720 94440 26880
rect 94280 26880 94440 27040
rect 94280 27040 94440 27200
rect 94280 27200 94440 27360
rect 94280 27360 94440 27520
rect 94280 27520 94440 27680
rect 94280 27680 94440 27840
rect 94280 27840 94440 28000
rect 94280 28000 94440 28160
rect 94280 28160 94440 28320
rect 94280 28320 94440 28480
rect 94280 28480 94440 28640
rect 94280 28640 94440 28800
rect 94280 28800 94440 28960
rect 94280 28960 94440 29120
rect 94280 29120 94440 29280
rect 94280 29280 94440 29440
rect 94280 29440 94440 29600
rect 94280 29600 94440 29760
rect 94280 29760 94440 29920
rect 94280 29920 94440 30080
rect 94280 30080 94440 30240
rect 94280 30240 94440 30400
rect 94280 30400 94440 30560
rect 94280 30560 94440 30720
rect 94280 30720 94440 30880
rect 94280 30880 94440 31040
rect 94280 31040 94440 31200
rect 94280 31200 94440 31360
rect 94280 31360 94440 31520
rect 94280 31520 94440 31680
rect 94280 31680 94440 31840
rect 94280 31840 94440 32000
rect 94280 32000 94440 32160
rect 94280 32160 94440 32320
rect 94280 32320 94440 32480
rect 94280 32480 94440 32640
rect 94280 32640 94440 32800
rect 94280 32800 94440 32960
rect 94280 32960 94440 33120
rect 94280 33120 94440 33280
rect 94280 33280 94440 33440
rect 94280 33440 94440 33600
rect 94280 33600 94440 33760
rect 94280 33760 94440 33920
rect 94280 33920 94440 34080
rect 94280 34080 94440 34240
rect 94280 34240 94440 34400
rect 94280 34400 94440 34560
rect 94280 34560 94440 34720
rect 94280 34720 94440 34880
rect 94280 34880 94440 35040
rect 94280 35040 94440 35200
rect 94280 35200 94440 35360
rect 94280 35360 94440 35520
rect 94280 35520 94440 35680
rect 94280 35680 94440 35840
rect 94280 35840 94440 36000
rect 94280 36000 94440 36160
rect 94280 36160 94440 36320
rect 94280 36320 94440 36480
rect 94280 36480 94440 36640
rect 94280 36640 94440 36800
rect 94280 36800 94440 36960
rect 94280 36960 94440 37120
rect 94280 37120 94440 37280
rect 94280 37280 94440 37440
rect 94280 37440 94440 37600
rect 94280 37600 94440 37760
rect 94280 37760 94440 37920
rect 94280 37920 94440 38080
rect 94280 38080 94440 38240
rect 94280 38240 94440 38400
rect 94280 38400 94440 38560
rect 94280 38560 94440 38720
rect 94280 38720 94440 38880
rect 94280 38880 94440 39040
rect 94280 39040 94440 39200
rect 94280 39200 94440 39360
rect 94280 39360 94440 39520
rect 94280 39520 94440 39680
rect 94280 39680 94440 39840
rect 94280 39840 94440 40000
rect 94280 40000 94440 40160
rect 94280 40160 94440 40320
rect 94280 40320 94440 40480
rect 94280 40480 94440 40640
rect 94280 40640 94440 40800
rect 94440 25600 94600 25760
rect 94440 25760 94600 25920
rect 94440 25920 94600 26080
rect 94440 26080 94600 26240
rect 94440 26240 94600 26400
rect 94440 26400 94600 26560
rect 94440 26560 94600 26720
rect 94440 26720 94600 26880
rect 94440 26880 94600 27040
rect 94440 27040 94600 27200
rect 94440 27200 94600 27360
rect 94440 27360 94600 27520
rect 94440 27520 94600 27680
rect 94440 27680 94600 27840
rect 94440 27840 94600 28000
rect 94440 28000 94600 28160
rect 94440 28160 94600 28320
rect 94440 28320 94600 28480
rect 94440 28480 94600 28640
rect 94440 28640 94600 28800
rect 94440 28800 94600 28960
rect 94440 28960 94600 29120
rect 94440 29120 94600 29280
rect 94440 29280 94600 29440
rect 94440 29440 94600 29600
rect 94440 29600 94600 29760
rect 94440 29760 94600 29920
rect 94440 29920 94600 30080
rect 94440 30080 94600 30240
rect 94440 30240 94600 30400
rect 94440 30400 94600 30560
rect 94440 30560 94600 30720
rect 94440 30720 94600 30880
rect 94440 30880 94600 31040
rect 94440 31040 94600 31200
rect 94440 31200 94600 31360
rect 94440 31360 94600 31520
rect 94440 31520 94600 31680
rect 94440 31680 94600 31840
rect 94440 31840 94600 32000
rect 94440 32000 94600 32160
rect 94440 32160 94600 32320
rect 94440 32320 94600 32480
rect 94440 32480 94600 32640
rect 94440 32640 94600 32800
rect 94440 32800 94600 32960
rect 94440 32960 94600 33120
rect 94440 33120 94600 33280
rect 94440 33280 94600 33440
rect 94440 33440 94600 33600
rect 94440 33600 94600 33760
rect 94440 33760 94600 33920
rect 94440 33920 94600 34080
rect 94440 34080 94600 34240
rect 94440 34240 94600 34400
rect 94440 34400 94600 34560
rect 94440 34560 94600 34720
rect 94440 34720 94600 34880
rect 94440 34880 94600 35040
rect 94440 35040 94600 35200
rect 94440 35200 94600 35360
rect 94440 35360 94600 35520
rect 94440 35520 94600 35680
rect 94440 35680 94600 35840
rect 94440 35840 94600 36000
rect 94440 36000 94600 36160
rect 94440 36160 94600 36320
rect 94440 36320 94600 36480
rect 94440 36480 94600 36640
rect 94440 36640 94600 36800
rect 94440 36800 94600 36960
rect 94440 36960 94600 37120
rect 94440 37120 94600 37280
rect 94440 37280 94600 37440
rect 94440 37440 94600 37600
rect 94440 37600 94600 37760
rect 94440 37760 94600 37920
rect 94440 37920 94600 38080
rect 94440 38080 94600 38240
rect 94440 38240 94600 38400
rect 94440 38400 94600 38560
rect 94440 38560 94600 38720
rect 94440 38720 94600 38880
rect 94440 38880 94600 39040
rect 94440 39040 94600 39200
rect 94440 39200 94600 39360
rect 94440 39360 94600 39520
rect 94440 39520 94600 39680
rect 94440 39680 94600 39840
rect 94440 39840 94600 40000
rect 94440 40000 94600 40160
rect 94440 40160 94600 40320
rect 94600 25440 94760 25600
rect 94600 25600 94760 25760
rect 94600 25760 94760 25920
rect 94600 25920 94760 26080
rect 94600 26080 94760 26240
rect 94600 26240 94760 26400
rect 94600 26400 94760 26560
rect 94600 26560 94760 26720
rect 94600 26720 94760 26880
rect 94600 26880 94760 27040
rect 94600 27040 94760 27200
rect 94600 27200 94760 27360
rect 94600 27360 94760 27520
rect 94600 27520 94760 27680
rect 94600 27680 94760 27840
rect 94600 27840 94760 28000
rect 94600 28000 94760 28160
rect 94600 28160 94760 28320
rect 94600 28320 94760 28480
rect 94600 28480 94760 28640
rect 94600 28640 94760 28800
rect 94600 28800 94760 28960
rect 94600 28960 94760 29120
rect 94600 29120 94760 29280
rect 94600 29280 94760 29440
rect 94600 29440 94760 29600
rect 94600 29600 94760 29760
rect 94600 29760 94760 29920
rect 94600 29920 94760 30080
rect 94600 30080 94760 30240
rect 94600 30240 94760 30400
rect 94600 30400 94760 30560
rect 94600 30560 94760 30720
rect 94600 30720 94760 30880
rect 94600 30880 94760 31040
rect 94600 31040 94760 31200
rect 94600 31200 94760 31360
rect 94600 31360 94760 31520
rect 94600 31520 94760 31680
rect 94600 31680 94760 31840
rect 94600 31840 94760 32000
rect 94600 32000 94760 32160
rect 94600 32160 94760 32320
rect 94600 32320 94760 32480
rect 94600 32480 94760 32640
rect 94600 32640 94760 32800
rect 94600 32800 94760 32960
rect 94600 32960 94760 33120
rect 94600 33120 94760 33280
rect 94600 33280 94760 33440
rect 94600 33440 94760 33600
rect 94600 33600 94760 33760
rect 94600 33760 94760 33920
rect 94600 33920 94760 34080
rect 94600 34080 94760 34240
rect 94600 34240 94760 34400
rect 94600 34400 94760 34560
rect 94600 34560 94760 34720
rect 94600 34720 94760 34880
rect 94600 34880 94760 35040
rect 94600 35040 94760 35200
rect 94600 35200 94760 35360
rect 94600 35360 94760 35520
rect 94600 35520 94760 35680
rect 94600 35680 94760 35840
rect 94600 35840 94760 36000
rect 94600 36000 94760 36160
rect 94600 36160 94760 36320
rect 94600 36320 94760 36480
rect 94600 36480 94760 36640
rect 94600 36640 94760 36800
rect 94600 36800 94760 36960
rect 94600 36960 94760 37120
rect 94600 37120 94760 37280
rect 94600 37280 94760 37440
rect 94600 37440 94760 37600
rect 94600 37600 94760 37760
rect 94600 37760 94760 37920
rect 94600 37920 94760 38080
rect 94600 38080 94760 38240
rect 94600 38240 94760 38400
rect 94600 38400 94760 38560
rect 94600 38560 94760 38720
rect 94600 38720 94760 38880
rect 94600 38880 94760 39040
rect 94600 39040 94760 39200
rect 94600 39200 94760 39360
rect 94600 39360 94760 39520
rect 94600 39520 94760 39680
rect 94600 39680 94760 39840
rect 94600 39840 94760 40000
rect 94760 25440 94920 25600
rect 94760 25600 94920 25760
rect 94760 25760 94920 25920
rect 94760 25920 94920 26080
rect 94760 26080 94920 26240
rect 94760 26240 94920 26400
rect 94760 26400 94920 26560
rect 94760 26560 94920 26720
rect 94760 26720 94920 26880
rect 94760 26880 94920 27040
rect 94760 27040 94920 27200
rect 94760 27200 94920 27360
rect 94760 27360 94920 27520
rect 94760 27520 94920 27680
rect 94760 27680 94920 27840
rect 94760 27840 94920 28000
rect 94760 28000 94920 28160
rect 94760 28160 94920 28320
rect 94760 28320 94920 28480
rect 94760 28480 94920 28640
rect 94760 28640 94920 28800
rect 94760 28800 94920 28960
rect 94760 28960 94920 29120
rect 94760 29120 94920 29280
rect 94760 29280 94920 29440
rect 94760 29440 94920 29600
rect 94760 29600 94920 29760
rect 94760 29760 94920 29920
rect 94760 29920 94920 30080
rect 94760 30080 94920 30240
rect 94760 30240 94920 30400
rect 94760 30400 94920 30560
rect 94760 30560 94920 30720
rect 94760 30720 94920 30880
rect 94760 30880 94920 31040
rect 94760 31040 94920 31200
rect 94760 31200 94920 31360
rect 94760 31360 94920 31520
rect 94760 31520 94920 31680
rect 94760 31680 94920 31840
rect 94760 31840 94920 32000
rect 94760 32000 94920 32160
rect 94760 32160 94920 32320
rect 94760 32320 94920 32480
rect 94760 32480 94920 32640
rect 94760 32640 94920 32800
rect 94760 32800 94920 32960
rect 94760 32960 94920 33120
rect 94760 33120 94920 33280
rect 94760 33280 94920 33440
rect 94760 33440 94920 33600
rect 94760 33600 94920 33760
rect 94760 33760 94920 33920
rect 94760 33920 94920 34080
rect 94760 34080 94920 34240
rect 94760 34240 94920 34400
rect 94760 34400 94920 34560
rect 94760 34560 94920 34720
rect 94760 34720 94920 34880
rect 94760 34880 94920 35040
rect 94760 35040 94920 35200
rect 94760 35200 94920 35360
rect 94760 35360 94920 35520
rect 94760 35520 94920 35680
rect 94760 35680 94920 35840
rect 94760 35840 94920 36000
rect 94760 36000 94920 36160
rect 94760 36160 94920 36320
rect 94760 36320 94920 36480
rect 94760 36480 94920 36640
rect 94760 36640 94920 36800
rect 94760 36800 94920 36960
rect 94760 36960 94920 37120
rect 94760 37120 94920 37280
rect 94760 37280 94920 37440
rect 94760 37440 94920 37600
rect 94760 37600 94920 37760
rect 94760 37760 94920 37920
rect 94760 37920 94920 38080
rect 94760 38080 94920 38240
rect 94760 38240 94920 38400
rect 94760 38400 94920 38560
rect 94760 38560 94920 38720
rect 94760 38720 94920 38880
rect 94760 38880 94920 39040
rect 94760 39040 94920 39200
rect 94760 39200 94920 39360
rect 94760 39360 94920 39520
rect 94920 25280 95080 25440
rect 94920 25440 95080 25600
rect 94920 25600 95080 25760
rect 94920 25760 95080 25920
rect 94920 25920 95080 26080
rect 94920 26080 95080 26240
rect 94920 26240 95080 26400
rect 94920 26400 95080 26560
rect 94920 26560 95080 26720
rect 94920 26720 95080 26880
rect 94920 26880 95080 27040
rect 94920 27040 95080 27200
rect 94920 27200 95080 27360
rect 94920 27360 95080 27520
rect 94920 27520 95080 27680
rect 94920 27680 95080 27840
rect 94920 27840 95080 28000
rect 94920 28000 95080 28160
rect 94920 28160 95080 28320
rect 94920 28320 95080 28480
rect 94920 28480 95080 28640
rect 94920 28640 95080 28800
rect 94920 28800 95080 28960
rect 94920 28960 95080 29120
rect 94920 29120 95080 29280
rect 94920 29280 95080 29440
rect 94920 29440 95080 29600
rect 94920 29600 95080 29760
rect 94920 29760 95080 29920
rect 94920 29920 95080 30080
rect 94920 30080 95080 30240
rect 94920 30240 95080 30400
rect 94920 30400 95080 30560
rect 94920 30560 95080 30720
rect 94920 30720 95080 30880
rect 94920 30880 95080 31040
rect 94920 31040 95080 31200
rect 94920 31200 95080 31360
rect 94920 31360 95080 31520
rect 94920 31520 95080 31680
rect 94920 31680 95080 31840
rect 94920 31840 95080 32000
rect 94920 32000 95080 32160
rect 94920 32160 95080 32320
rect 94920 32320 95080 32480
rect 94920 32480 95080 32640
rect 94920 32640 95080 32800
rect 94920 32800 95080 32960
rect 94920 32960 95080 33120
rect 94920 33120 95080 33280
rect 94920 33280 95080 33440
rect 94920 33440 95080 33600
rect 94920 33600 95080 33760
rect 94920 33760 95080 33920
rect 94920 33920 95080 34080
rect 94920 34080 95080 34240
rect 94920 34240 95080 34400
rect 94920 34400 95080 34560
rect 94920 34560 95080 34720
rect 94920 34720 95080 34880
rect 94920 34880 95080 35040
rect 94920 35040 95080 35200
rect 94920 35200 95080 35360
rect 94920 35360 95080 35520
rect 94920 35520 95080 35680
rect 94920 35680 95080 35840
rect 94920 35840 95080 36000
rect 94920 36000 95080 36160
rect 94920 36160 95080 36320
rect 94920 36320 95080 36480
rect 94920 36480 95080 36640
rect 94920 36640 95080 36800
rect 94920 36800 95080 36960
rect 94920 36960 95080 37120
rect 94920 37120 95080 37280
rect 94920 37280 95080 37440
rect 94920 37440 95080 37600
rect 94920 37600 95080 37760
rect 94920 37760 95080 37920
rect 94920 37920 95080 38080
rect 94920 38080 95080 38240
rect 94920 38240 95080 38400
rect 94920 38400 95080 38560
rect 94920 38560 95080 38720
rect 94920 38720 95080 38880
rect 94920 38880 95080 39040
rect 95080 25280 95240 25440
rect 95080 25440 95240 25600
rect 95080 25600 95240 25760
rect 95080 25760 95240 25920
rect 95080 25920 95240 26080
rect 95080 26080 95240 26240
rect 95080 26240 95240 26400
rect 95080 26400 95240 26560
rect 95080 26560 95240 26720
rect 95080 26720 95240 26880
rect 95080 26880 95240 27040
rect 95080 27040 95240 27200
rect 95080 27200 95240 27360
rect 95080 27360 95240 27520
rect 95080 27520 95240 27680
rect 95080 27680 95240 27840
rect 95080 27840 95240 28000
rect 95080 28000 95240 28160
rect 95080 28160 95240 28320
rect 95080 28320 95240 28480
rect 95080 28480 95240 28640
rect 95080 28640 95240 28800
rect 95080 28800 95240 28960
rect 95080 28960 95240 29120
rect 95080 29120 95240 29280
rect 95080 29280 95240 29440
rect 95080 29440 95240 29600
rect 95080 29600 95240 29760
rect 95080 29760 95240 29920
rect 95080 29920 95240 30080
rect 95080 30080 95240 30240
rect 95080 30240 95240 30400
rect 95080 30400 95240 30560
rect 95080 30560 95240 30720
rect 95080 30720 95240 30880
rect 95080 30880 95240 31040
rect 95080 31040 95240 31200
rect 95080 31200 95240 31360
rect 95080 31360 95240 31520
rect 95080 31520 95240 31680
rect 95080 31680 95240 31840
rect 95080 31840 95240 32000
rect 95080 32000 95240 32160
rect 95080 32160 95240 32320
rect 95080 32320 95240 32480
rect 95080 32480 95240 32640
rect 95080 32640 95240 32800
rect 95080 32800 95240 32960
rect 95080 32960 95240 33120
rect 95080 33120 95240 33280
rect 95080 33280 95240 33440
rect 95080 33440 95240 33600
rect 95080 33600 95240 33760
rect 95080 33760 95240 33920
rect 95080 33920 95240 34080
rect 95080 34080 95240 34240
rect 95080 34240 95240 34400
rect 95080 34400 95240 34560
rect 95080 34560 95240 34720
rect 95080 34720 95240 34880
rect 95080 34880 95240 35040
rect 95080 35040 95240 35200
rect 95080 35200 95240 35360
rect 95080 35360 95240 35520
rect 95080 35520 95240 35680
rect 95080 35680 95240 35840
rect 95080 35840 95240 36000
rect 95080 36000 95240 36160
rect 95080 36160 95240 36320
rect 95080 36320 95240 36480
rect 95080 36480 95240 36640
rect 95080 36640 95240 36800
rect 95080 36800 95240 36960
rect 95080 36960 95240 37120
rect 95080 37120 95240 37280
rect 95080 37280 95240 37440
rect 95080 37440 95240 37600
rect 95080 37600 95240 37760
rect 95080 37760 95240 37920
rect 95080 37920 95240 38080
rect 95080 38080 95240 38240
rect 95080 38240 95240 38400
rect 95080 38400 95240 38560
rect 95240 25280 95400 25440
rect 95240 25440 95400 25600
rect 95240 25600 95400 25760
rect 95240 25760 95400 25920
rect 95240 25920 95400 26080
rect 95240 26080 95400 26240
rect 95240 26240 95400 26400
rect 95240 26400 95400 26560
rect 95240 26560 95400 26720
rect 95240 26720 95400 26880
rect 95240 26880 95400 27040
rect 95240 27040 95400 27200
rect 95240 27200 95400 27360
rect 95240 27360 95400 27520
rect 95240 27520 95400 27680
rect 95240 27680 95400 27840
rect 95240 27840 95400 28000
rect 95240 28000 95400 28160
rect 95240 28160 95400 28320
rect 95240 28320 95400 28480
rect 95240 28480 95400 28640
rect 95240 28640 95400 28800
rect 95240 28800 95400 28960
rect 95240 28960 95400 29120
rect 95240 29120 95400 29280
rect 95240 29280 95400 29440
rect 95240 29440 95400 29600
rect 95240 29600 95400 29760
rect 95240 29760 95400 29920
rect 95240 29920 95400 30080
rect 95240 30080 95400 30240
rect 95240 30240 95400 30400
rect 95240 30400 95400 30560
rect 95240 30560 95400 30720
rect 95240 30720 95400 30880
rect 95240 30880 95400 31040
rect 95240 31040 95400 31200
rect 95240 31200 95400 31360
rect 95240 31360 95400 31520
rect 95240 31520 95400 31680
rect 95240 31680 95400 31840
rect 95240 31840 95400 32000
rect 95240 32000 95400 32160
rect 95240 32160 95400 32320
rect 95240 32320 95400 32480
rect 95240 32480 95400 32640
rect 95240 32640 95400 32800
rect 95240 32800 95400 32960
rect 95240 32960 95400 33120
rect 95240 33120 95400 33280
rect 95240 33280 95400 33440
rect 95240 33440 95400 33600
rect 95240 33600 95400 33760
rect 95240 33760 95400 33920
rect 95240 33920 95400 34080
rect 95240 34080 95400 34240
rect 95240 34240 95400 34400
rect 95240 34400 95400 34560
rect 95240 34560 95400 34720
rect 95240 34720 95400 34880
rect 95240 34880 95400 35040
rect 95240 35040 95400 35200
rect 95240 35200 95400 35360
rect 95240 35360 95400 35520
rect 95240 35520 95400 35680
rect 95240 35680 95400 35840
rect 95240 35840 95400 36000
rect 95240 36000 95400 36160
rect 95240 36160 95400 36320
rect 95240 36320 95400 36480
rect 95240 36480 95400 36640
rect 95240 36640 95400 36800
rect 95240 36800 95400 36960
rect 95240 36960 95400 37120
rect 95240 37120 95400 37280
rect 95240 37280 95400 37440
rect 95240 37440 95400 37600
rect 95240 37600 95400 37760
rect 95240 37760 95400 37920
rect 95240 37920 95400 38080
rect 95400 25280 95560 25440
rect 95400 25440 95560 25600
rect 95400 25600 95560 25760
rect 95400 25760 95560 25920
rect 95400 25920 95560 26080
rect 95400 26080 95560 26240
rect 95400 26240 95560 26400
rect 95400 26400 95560 26560
rect 95400 26560 95560 26720
rect 95400 26720 95560 26880
rect 95400 26880 95560 27040
rect 95400 27040 95560 27200
rect 95400 27200 95560 27360
rect 95400 27360 95560 27520
rect 95400 27520 95560 27680
rect 95400 27680 95560 27840
rect 95400 27840 95560 28000
rect 95400 28000 95560 28160
rect 95400 28160 95560 28320
rect 95400 28320 95560 28480
rect 95400 28480 95560 28640
rect 95400 28640 95560 28800
rect 95400 28800 95560 28960
rect 95400 28960 95560 29120
rect 95400 29120 95560 29280
rect 95400 29280 95560 29440
rect 95400 29440 95560 29600
rect 95400 29600 95560 29760
rect 95400 29760 95560 29920
rect 95400 29920 95560 30080
rect 95400 30080 95560 30240
rect 95400 30240 95560 30400
rect 95400 30400 95560 30560
rect 95400 30560 95560 30720
rect 95400 30720 95560 30880
rect 95400 30880 95560 31040
rect 95400 31040 95560 31200
rect 95400 31200 95560 31360
rect 95400 31360 95560 31520
rect 95400 31520 95560 31680
rect 95400 31680 95560 31840
rect 95400 31840 95560 32000
rect 95400 32000 95560 32160
rect 95400 32160 95560 32320
rect 95400 32320 95560 32480
rect 95400 32480 95560 32640
rect 95400 32640 95560 32800
rect 95400 32800 95560 32960
rect 95400 32960 95560 33120
rect 95400 33120 95560 33280
rect 95400 33280 95560 33440
rect 95400 33440 95560 33600
rect 95400 33600 95560 33760
rect 95400 33760 95560 33920
rect 95400 33920 95560 34080
rect 95400 34080 95560 34240
rect 95400 34240 95560 34400
rect 95400 34400 95560 34560
rect 95400 34560 95560 34720
rect 95400 34720 95560 34880
rect 95400 34880 95560 35040
rect 95400 35040 95560 35200
rect 95400 35200 95560 35360
rect 95400 35360 95560 35520
rect 95400 35520 95560 35680
rect 95400 35680 95560 35840
rect 95400 35840 95560 36000
rect 95400 36000 95560 36160
rect 95400 36160 95560 36320
rect 95400 36320 95560 36480
rect 95400 36480 95560 36640
rect 95400 36640 95560 36800
rect 95400 36800 95560 36960
rect 95400 36960 95560 37120
rect 95400 37120 95560 37280
rect 95400 37280 95560 37440
rect 95400 37440 95560 37600
rect 95560 25120 95720 25280
rect 95560 25280 95720 25440
rect 95560 25440 95720 25600
rect 95560 25600 95720 25760
rect 95560 25760 95720 25920
rect 95560 25920 95720 26080
rect 95560 26080 95720 26240
rect 95560 26240 95720 26400
rect 95560 26400 95720 26560
rect 95560 26560 95720 26720
rect 95560 26720 95720 26880
rect 95560 26880 95720 27040
rect 95560 27040 95720 27200
rect 95560 27200 95720 27360
rect 95560 27360 95720 27520
rect 95560 27520 95720 27680
rect 95560 27680 95720 27840
rect 95560 27840 95720 28000
rect 95560 28000 95720 28160
rect 95560 28160 95720 28320
rect 95560 28320 95720 28480
rect 95560 28480 95720 28640
rect 95560 28640 95720 28800
rect 95560 28800 95720 28960
rect 95560 28960 95720 29120
rect 95560 30080 95720 30240
rect 95560 30240 95720 30400
rect 95560 30400 95720 30560
rect 95560 30560 95720 30720
rect 95560 30720 95720 30880
rect 95560 30880 95720 31040
rect 95560 31040 95720 31200
rect 95560 31200 95720 31360
rect 95560 31360 95720 31520
rect 95560 31520 95720 31680
rect 95560 31680 95720 31840
rect 95560 31840 95720 32000
rect 95560 32000 95720 32160
rect 95560 32160 95720 32320
rect 95560 32320 95720 32480
rect 95560 32480 95720 32640
rect 95560 32640 95720 32800
rect 95560 32800 95720 32960
rect 95560 32960 95720 33120
rect 95560 33120 95720 33280
rect 95560 33280 95720 33440
rect 95560 33440 95720 33600
rect 95560 33600 95720 33760
rect 95560 33760 95720 33920
rect 95560 33920 95720 34080
rect 95560 34080 95720 34240
rect 95560 34240 95720 34400
rect 95560 34400 95720 34560
rect 95560 34560 95720 34720
rect 95560 34720 95720 34880
rect 95560 34880 95720 35040
rect 95560 35040 95720 35200
rect 95560 35200 95720 35360
rect 95560 35360 95720 35520
rect 95560 35520 95720 35680
rect 95560 35680 95720 35840
rect 95560 35840 95720 36000
rect 95560 36000 95720 36160
rect 95560 36160 95720 36320
rect 95560 36320 95720 36480
rect 95560 36480 95720 36640
rect 95560 36640 95720 36800
rect 95560 36800 95720 36960
rect 95560 36960 95720 37120
rect 95560 37120 95720 37280
rect 95720 25120 95880 25280
rect 95720 25280 95880 25440
rect 95720 25440 95880 25600
rect 95720 25600 95880 25760
rect 95720 25760 95880 25920
rect 95720 25920 95880 26080
rect 95720 26080 95880 26240
rect 95720 26240 95880 26400
rect 95720 26400 95880 26560
rect 95720 26560 95880 26720
rect 95720 26720 95880 26880
rect 95720 26880 95880 27040
rect 95720 27040 95880 27200
rect 95720 27200 95880 27360
rect 95720 27360 95880 27520
rect 95720 27520 95880 27680
rect 95720 27680 95880 27840
rect 95720 27840 95880 28000
rect 95720 28000 95880 28160
rect 95720 28160 95880 28320
rect 95720 28320 95880 28480
rect 95720 28480 95880 28640
rect 95720 28640 95880 28800
rect 95720 30240 95880 30400
rect 95720 30400 95880 30560
rect 95720 30560 95880 30720
rect 95720 30720 95880 30880
rect 95720 30880 95880 31040
rect 95720 31040 95880 31200
rect 95720 31200 95880 31360
rect 95720 31360 95880 31520
rect 95720 31520 95880 31680
rect 95720 31680 95880 31840
rect 95720 31840 95880 32000
rect 95720 32000 95880 32160
rect 95720 32160 95880 32320
rect 95720 32320 95880 32480
rect 95720 32480 95880 32640
rect 95720 32640 95880 32800
rect 95720 32800 95880 32960
rect 95720 32960 95880 33120
rect 95720 33120 95880 33280
rect 95720 33280 95880 33440
rect 95720 33440 95880 33600
rect 95720 33600 95880 33760
rect 95720 33760 95880 33920
rect 95720 33920 95880 34080
rect 95720 34080 95880 34240
rect 95720 34240 95880 34400
rect 95720 34400 95880 34560
rect 95720 34560 95880 34720
rect 95720 34720 95880 34880
rect 95720 34880 95880 35040
rect 95720 35040 95880 35200
rect 95720 35200 95880 35360
rect 95720 35360 95880 35520
rect 95720 35520 95880 35680
rect 95720 35680 95880 35840
rect 95720 35840 95880 36000
rect 95720 36000 95880 36160
rect 95720 36160 95880 36320
rect 95720 36320 95880 36480
rect 95720 36480 95880 36640
rect 95720 36640 95880 36800
rect 95880 25120 96040 25280
rect 95880 25280 96040 25440
rect 95880 25440 96040 25600
rect 95880 25600 96040 25760
rect 95880 25760 96040 25920
rect 95880 25920 96040 26080
rect 95880 26080 96040 26240
rect 95880 26240 96040 26400
rect 95880 26400 96040 26560
rect 95880 26560 96040 26720
rect 95880 26720 96040 26880
rect 95880 26880 96040 27040
rect 95880 27040 96040 27200
rect 95880 27200 96040 27360
rect 95880 27360 96040 27520
rect 95880 27520 96040 27680
rect 95880 27680 96040 27840
rect 95880 27840 96040 28000
rect 95880 28000 96040 28160
rect 95880 28160 96040 28320
rect 95880 28320 96040 28480
rect 95880 28480 96040 28640
rect 95880 30240 96040 30400
rect 95880 30400 96040 30560
rect 95880 30560 96040 30720
rect 95880 30720 96040 30880
rect 95880 30880 96040 31040
rect 95880 31040 96040 31200
rect 95880 31200 96040 31360
rect 95880 31360 96040 31520
rect 95880 31520 96040 31680
rect 95880 31680 96040 31840
rect 95880 31840 96040 32000
rect 95880 32000 96040 32160
rect 95880 32160 96040 32320
rect 95880 32320 96040 32480
rect 95880 32480 96040 32640
rect 95880 32640 96040 32800
rect 95880 32800 96040 32960
rect 95880 32960 96040 33120
rect 95880 33120 96040 33280
rect 95880 33280 96040 33440
rect 95880 33440 96040 33600
rect 95880 33600 96040 33760
rect 95880 33760 96040 33920
rect 95880 33920 96040 34080
rect 95880 34080 96040 34240
rect 95880 34240 96040 34400
rect 95880 34400 96040 34560
rect 95880 34560 96040 34720
rect 95880 34720 96040 34880
rect 95880 34880 96040 35040
rect 95880 35040 96040 35200
rect 95880 35200 96040 35360
rect 95880 35360 96040 35520
rect 95880 35520 96040 35680
rect 95880 35680 96040 35840
rect 95880 35840 96040 36000
rect 95880 36000 96040 36160
rect 95880 36160 96040 36320
rect 96040 25120 96200 25280
rect 96040 25280 96200 25440
rect 96040 25440 96200 25600
rect 96040 25600 96200 25760
rect 96040 25760 96200 25920
rect 96040 25920 96200 26080
rect 96040 26080 96200 26240
rect 96040 26240 96200 26400
rect 96040 26400 96200 26560
rect 96040 26560 96200 26720
rect 96040 26720 96200 26880
rect 96040 26880 96200 27040
rect 96040 27040 96200 27200
rect 96040 27200 96200 27360
rect 96040 27360 96200 27520
rect 96040 27520 96200 27680
rect 96040 27680 96200 27840
rect 96040 27840 96200 28000
rect 96040 28000 96200 28160
rect 96040 28160 96200 28320
rect 96040 28320 96200 28480
rect 96040 30240 96200 30400
rect 96040 30400 96200 30560
rect 96040 30560 96200 30720
rect 96040 30720 96200 30880
rect 96040 30880 96200 31040
rect 96040 31040 96200 31200
rect 96040 31200 96200 31360
rect 96040 31360 96200 31520
rect 96040 31520 96200 31680
rect 96040 31680 96200 31840
rect 96040 31840 96200 32000
rect 96040 32000 96200 32160
rect 96040 32160 96200 32320
rect 96040 32320 96200 32480
rect 96040 32480 96200 32640
rect 96040 32640 96200 32800
rect 96040 32800 96200 32960
rect 96040 32960 96200 33120
rect 96040 33120 96200 33280
rect 96040 33280 96200 33440
rect 96040 33440 96200 33600
rect 96040 33600 96200 33760
rect 96040 33760 96200 33920
rect 96040 33920 96200 34080
rect 96040 34080 96200 34240
rect 96040 34240 96200 34400
rect 96040 34400 96200 34560
rect 96040 34560 96200 34720
rect 96040 34720 96200 34880
rect 96040 34880 96200 35040
rect 96040 35040 96200 35200
rect 96040 35200 96200 35360
rect 96040 35360 96200 35520
rect 96040 35520 96200 35680
rect 96040 35680 96200 35840
rect 96040 35840 96200 36000
rect 96200 25120 96360 25280
rect 96200 25280 96360 25440
rect 96200 25440 96360 25600
rect 96200 25600 96360 25760
rect 96200 25760 96360 25920
rect 96200 25920 96360 26080
rect 96200 26080 96360 26240
rect 96200 26240 96360 26400
rect 96200 26400 96360 26560
rect 96200 26560 96360 26720
rect 96200 26720 96360 26880
rect 96200 26880 96360 27040
rect 96200 27040 96360 27200
rect 96200 27200 96360 27360
rect 96200 27360 96360 27520
rect 96200 27520 96360 27680
rect 96200 27680 96360 27840
rect 96200 27840 96360 28000
rect 96200 28000 96360 28160
rect 96200 28160 96360 28320
rect 96200 28320 96360 28480
rect 96200 30240 96360 30400
rect 96200 30400 96360 30560
rect 96200 30560 96360 30720
rect 96200 30720 96360 30880
rect 96200 30880 96360 31040
rect 96200 31040 96360 31200
rect 96200 31200 96360 31360
rect 96200 31360 96360 31520
rect 96200 31520 96360 31680
rect 96200 31680 96360 31840
rect 96200 31840 96360 32000
rect 96200 32000 96360 32160
rect 96200 32160 96360 32320
rect 96200 32320 96360 32480
rect 96200 32480 96360 32640
rect 96200 32640 96360 32800
rect 96200 32800 96360 32960
rect 96200 32960 96360 33120
rect 96200 33120 96360 33280
rect 96200 33280 96360 33440
rect 96200 33440 96360 33600
rect 96200 33600 96360 33760
rect 96200 33760 96360 33920
rect 96200 33920 96360 34080
rect 96200 34080 96360 34240
rect 96200 34240 96360 34400
rect 96200 34400 96360 34560
rect 96200 34560 96360 34720
rect 96200 34720 96360 34880
rect 96200 34880 96360 35040
rect 96200 35040 96360 35200
rect 96200 35200 96360 35360
rect 96200 35360 96360 35520
rect 96360 25120 96520 25280
rect 96360 25280 96520 25440
rect 96360 25440 96520 25600
rect 96360 25600 96520 25760
rect 96360 25760 96520 25920
rect 96360 25920 96520 26080
rect 96360 26080 96520 26240
rect 96360 26240 96520 26400
rect 96360 26400 96520 26560
rect 96360 26560 96520 26720
rect 96360 26720 96520 26880
rect 96360 26880 96520 27040
rect 96360 27040 96520 27200
rect 96360 27200 96520 27360
rect 96360 27360 96520 27520
rect 96360 27520 96520 27680
rect 96360 27680 96520 27840
rect 96360 27840 96520 28000
rect 96360 28000 96520 28160
rect 96360 28160 96520 28320
rect 96360 28320 96520 28480
rect 96360 30240 96520 30400
rect 96360 30400 96520 30560
rect 96360 30560 96520 30720
rect 96360 30720 96520 30880
rect 96360 30880 96520 31040
rect 96360 31040 96520 31200
rect 96360 31200 96520 31360
rect 96360 31360 96520 31520
rect 96360 31520 96520 31680
rect 96360 31680 96520 31840
rect 96360 31840 96520 32000
rect 96360 32000 96520 32160
rect 96360 32160 96520 32320
rect 96360 32320 96520 32480
rect 96360 32480 96520 32640
rect 96360 32640 96520 32800
rect 96360 32800 96520 32960
rect 96360 32960 96520 33120
rect 96360 33120 96520 33280
rect 96360 33280 96520 33440
rect 96360 33440 96520 33600
rect 96360 33600 96520 33760
rect 96360 33760 96520 33920
rect 96360 33920 96520 34080
rect 96360 34080 96520 34240
rect 96360 34240 96520 34400
rect 96360 34400 96520 34560
rect 96360 34560 96520 34720
rect 96360 34720 96520 34880
rect 96360 34880 96520 35040
rect 96360 35040 96520 35200
rect 96520 25280 96680 25440
rect 96520 25440 96680 25600
rect 96520 25600 96680 25760
rect 96520 25760 96680 25920
rect 96520 25920 96680 26080
rect 96520 26080 96680 26240
rect 96520 26240 96680 26400
rect 96520 26400 96680 26560
rect 96520 26560 96680 26720
rect 96520 26720 96680 26880
rect 96520 26880 96680 27040
rect 96520 27040 96680 27200
rect 96520 27200 96680 27360
rect 96520 27360 96680 27520
rect 96520 27520 96680 27680
rect 96520 27680 96680 27840
rect 96520 27840 96680 28000
rect 96520 28000 96680 28160
rect 96520 28160 96680 28320
rect 96520 30240 96680 30400
rect 96520 30400 96680 30560
rect 96520 30560 96680 30720
rect 96520 30720 96680 30880
rect 96520 30880 96680 31040
rect 96520 31040 96680 31200
rect 96520 31200 96680 31360
rect 96520 31360 96680 31520
rect 96520 31520 96680 31680
rect 96520 31680 96680 31840
rect 96520 31840 96680 32000
rect 96520 32000 96680 32160
rect 96520 32160 96680 32320
rect 96520 32320 96680 32480
rect 96520 32480 96680 32640
rect 96520 32640 96680 32800
rect 96520 32800 96680 32960
rect 96520 32960 96680 33120
rect 96520 33120 96680 33280
rect 96520 33280 96680 33440
rect 96520 33440 96680 33600
rect 96520 33600 96680 33760
rect 96520 33760 96680 33920
rect 96520 33920 96680 34080
rect 96520 34080 96680 34240
rect 96520 34240 96680 34400
rect 96520 34400 96680 34560
rect 96520 34560 96680 34720
rect 96520 34720 96680 34880
rect 96680 25280 96840 25440
rect 96680 25440 96840 25600
rect 96680 25600 96840 25760
rect 96680 25760 96840 25920
rect 96680 25920 96840 26080
rect 96680 26080 96840 26240
rect 96680 26240 96840 26400
rect 96680 26400 96840 26560
rect 96680 26560 96840 26720
rect 96680 26720 96840 26880
rect 96680 26880 96840 27040
rect 96680 27040 96840 27200
rect 96680 27200 96840 27360
rect 96680 27360 96840 27520
rect 96680 27520 96840 27680
rect 96680 27680 96840 27840
rect 96680 27840 96840 28000
rect 96680 28000 96840 28160
rect 96680 28160 96840 28320
rect 96680 30240 96840 30400
rect 96680 30400 96840 30560
rect 96680 30560 96840 30720
rect 96680 30720 96840 30880
rect 96680 30880 96840 31040
rect 96680 31040 96840 31200
rect 96680 31200 96840 31360
rect 96680 31360 96840 31520
rect 96680 31520 96840 31680
rect 96680 31680 96840 31840
rect 96680 31840 96840 32000
rect 96680 32000 96840 32160
rect 96680 32160 96840 32320
rect 96680 32320 96840 32480
rect 96680 32480 96840 32640
rect 96680 32640 96840 32800
rect 96680 32800 96840 32960
rect 96680 32960 96840 33120
rect 96680 33120 96840 33280
rect 96680 33280 96840 33440
rect 96680 33440 96840 33600
rect 96680 33600 96840 33760
rect 96680 33760 96840 33920
rect 96680 33920 96840 34080
rect 96680 34080 96840 34240
rect 96680 34240 96840 34400
rect 96680 34400 96840 34560
rect 96680 34560 96840 34720
rect 96840 25280 97000 25440
rect 96840 25440 97000 25600
rect 96840 25600 97000 25760
rect 96840 25760 97000 25920
rect 96840 25920 97000 26080
rect 96840 26080 97000 26240
rect 96840 26240 97000 26400
rect 96840 26400 97000 26560
rect 96840 26560 97000 26720
rect 96840 26720 97000 26880
rect 96840 26880 97000 27040
rect 96840 27040 97000 27200
rect 96840 27200 97000 27360
rect 96840 27360 97000 27520
rect 96840 27520 97000 27680
rect 96840 27680 97000 27840
rect 96840 27840 97000 28000
rect 96840 28000 97000 28160
rect 96840 28160 97000 28320
rect 96840 30240 97000 30400
rect 96840 30400 97000 30560
rect 96840 30560 97000 30720
rect 96840 30720 97000 30880
rect 96840 30880 97000 31040
rect 96840 31040 97000 31200
rect 96840 31200 97000 31360
rect 96840 31360 97000 31520
rect 96840 31520 97000 31680
rect 96840 31680 97000 31840
rect 96840 31840 97000 32000
rect 96840 32000 97000 32160
rect 96840 32160 97000 32320
rect 96840 32320 97000 32480
rect 96840 32480 97000 32640
rect 96840 32640 97000 32800
rect 96840 32800 97000 32960
rect 96840 32960 97000 33120
rect 96840 33120 97000 33280
rect 96840 33280 97000 33440
rect 96840 33440 97000 33600
rect 96840 33600 97000 33760
rect 96840 33760 97000 33920
rect 96840 33920 97000 34080
rect 96840 34080 97000 34240
rect 96840 34240 97000 34400
rect 97000 25280 97160 25440
rect 97000 25440 97160 25600
rect 97000 25600 97160 25760
rect 97000 25760 97160 25920
rect 97000 25920 97160 26080
rect 97000 26080 97160 26240
rect 97000 26240 97160 26400
rect 97000 26400 97160 26560
rect 97000 26560 97160 26720
rect 97000 26720 97160 26880
rect 97000 26880 97160 27040
rect 97000 27040 97160 27200
rect 97000 27200 97160 27360
rect 97000 27360 97160 27520
rect 97000 27520 97160 27680
rect 97000 27680 97160 27840
rect 97000 27840 97160 28000
rect 97000 28000 97160 28160
rect 97000 28160 97160 28320
rect 97000 28320 97160 28480
rect 97000 30080 97160 30240
rect 97000 30240 97160 30400
rect 97000 30400 97160 30560
rect 97000 30560 97160 30720
rect 97000 30720 97160 30880
rect 97000 30880 97160 31040
rect 97000 31040 97160 31200
rect 97000 31200 97160 31360
rect 97000 31360 97160 31520
rect 97000 31520 97160 31680
rect 97000 31680 97160 31840
rect 97000 31840 97160 32000
rect 97000 32000 97160 32160
rect 97000 32160 97160 32320
rect 97000 32320 97160 32480
rect 97000 32480 97160 32640
rect 97000 32640 97160 32800
rect 97000 32800 97160 32960
rect 97000 32960 97160 33120
rect 97000 33120 97160 33280
rect 97000 33280 97160 33440
rect 97000 33440 97160 33600
rect 97000 33600 97160 33760
rect 97000 33760 97160 33920
rect 97000 33920 97160 34080
rect 97000 34080 97160 34240
rect 97160 25440 97320 25600
rect 97160 25600 97320 25760
rect 97160 25760 97320 25920
rect 97160 25920 97320 26080
rect 97160 26080 97320 26240
rect 97160 26240 97320 26400
rect 97160 26400 97320 26560
rect 97160 26560 97320 26720
rect 97160 26720 97320 26880
rect 97160 26880 97320 27040
rect 97160 27040 97320 27200
rect 97160 27200 97320 27360
rect 97160 27360 97320 27520
rect 97160 27520 97320 27680
rect 97160 27680 97320 27840
rect 97160 27840 97320 28000
rect 97160 28000 97320 28160
rect 97160 28160 97320 28320
rect 97160 28320 97320 28480
rect 97160 30080 97320 30240
rect 97160 30240 97320 30400
rect 97160 30400 97320 30560
rect 97160 30560 97320 30720
rect 97160 30720 97320 30880
rect 97160 30880 97320 31040
rect 97160 31040 97320 31200
rect 97160 31200 97320 31360
rect 97160 31360 97320 31520
rect 97160 31520 97320 31680
rect 97160 31680 97320 31840
rect 97160 31840 97320 32000
rect 97160 32000 97320 32160
rect 97160 32160 97320 32320
rect 97160 32320 97320 32480
rect 97160 32480 97320 32640
rect 97160 32640 97320 32800
rect 97160 32800 97320 32960
rect 97160 32960 97320 33120
rect 97160 33120 97320 33280
rect 97160 33280 97320 33440
rect 97160 33440 97320 33600
rect 97160 33600 97320 33760
rect 97160 33760 97320 33920
rect 97160 33920 97320 34080
rect 97320 25440 97480 25600
rect 97320 25600 97480 25760
rect 97320 25760 97480 25920
rect 97320 25920 97480 26080
rect 97320 26080 97480 26240
rect 97320 26240 97480 26400
rect 97320 26400 97480 26560
rect 97320 26560 97480 26720
rect 97320 26720 97480 26880
rect 97320 26880 97480 27040
rect 97320 27040 97480 27200
rect 97320 27200 97480 27360
rect 97320 27360 97480 27520
rect 97320 27520 97480 27680
rect 97320 27680 97480 27840
rect 97320 27840 97480 28000
rect 97320 28000 97480 28160
rect 97320 28160 97480 28320
rect 97320 28320 97480 28480
rect 97320 29920 97480 30080
rect 97320 30080 97480 30240
rect 97320 30240 97480 30400
rect 97320 30400 97480 30560
rect 97320 30560 97480 30720
rect 97320 30720 97480 30880
rect 97320 30880 97480 31040
rect 97320 31040 97480 31200
rect 97320 31200 97480 31360
rect 97320 31360 97480 31520
rect 97320 31520 97480 31680
rect 97320 31680 97480 31840
rect 97320 31840 97480 32000
rect 97320 32000 97480 32160
rect 97320 32160 97480 32320
rect 97320 32320 97480 32480
rect 97320 32480 97480 32640
rect 97320 32640 97480 32800
rect 97320 32800 97480 32960
rect 97320 32960 97480 33120
rect 97320 33120 97480 33280
rect 97320 33280 97480 33440
rect 97320 33440 97480 33600
rect 97320 33600 97480 33760
rect 97320 33760 97480 33920
rect 97480 25440 97640 25600
rect 97480 25600 97640 25760
rect 97480 25760 97640 25920
rect 97480 25920 97640 26080
rect 97480 26080 97640 26240
rect 97480 26240 97640 26400
rect 97480 26400 97640 26560
rect 97480 26560 97640 26720
rect 97480 26720 97640 26880
rect 97480 26880 97640 27040
rect 97480 27040 97640 27200
rect 97480 27200 97640 27360
rect 97480 27360 97640 27520
rect 97480 27520 97640 27680
rect 97480 27680 97640 27840
rect 97480 27840 97640 28000
rect 97480 28000 97640 28160
rect 97480 28160 97640 28320
rect 97480 28320 97640 28480
rect 97480 28480 97640 28640
rect 97480 28640 97640 28800
rect 97480 29760 97640 29920
rect 97480 29920 97640 30080
rect 97480 30080 97640 30240
rect 97480 30240 97640 30400
rect 97480 30400 97640 30560
rect 97480 30560 97640 30720
rect 97480 30720 97640 30880
rect 97480 30880 97640 31040
rect 97480 31040 97640 31200
rect 97480 31200 97640 31360
rect 97480 31360 97640 31520
rect 97480 31520 97640 31680
rect 97480 31680 97640 31840
rect 97480 31840 97640 32000
rect 97480 32000 97640 32160
rect 97480 32160 97640 32320
rect 97480 32320 97640 32480
rect 97480 32480 97640 32640
rect 97480 32640 97640 32800
rect 97480 32800 97640 32960
rect 97480 32960 97640 33120
rect 97480 33120 97640 33280
rect 97480 33280 97640 33440
rect 97480 33440 97640 33600
rect 97480 33600 97640 33760
rect 97640 25600 97800 25760
rect 97640 25760 97800 25920
rect 97640 25920 97800 26080
rect 97640 26080 97800 26240
rect 97640 26240 97800 26400
rect 97640 26400 97800 26560
rect 97640 26560 97800 26720
rect 97640 26720 97800 26880
rect 97640 26880 97800 27040
rect 97640 27040 97800 27200
rect 97640 27200 97800 27360
rect 97640 27360 97800 27520
rect 97640 27520 97800 27680
rect 97640 27680 97800 27840
rect 97640 27840 97800 28000
rect 97640 28000 97800 28160
rect 97640 28160 97800 28320
rect 97640 28320 97800 28480
rect 97640 28480 97800 28640
rect 97640 28640 97800 28800
rect 97640 28800 97800 28960
rect 97640 28960 97800 29120
rect 97640 29120 97800 29280
rect 97640 29280 97800 29440
rect 97640 29440 97800 29600
rect 97640 29600 97800 29760
rect 97640 29760 97800 29920
rect 97640 29920 97800 30080
rect 97640 30080 97800 30240
rect 97640 30240 97800 30400
rect 97640 30400 97800 30560
rect 97640 30560 97800 30720
rect 97640 30720 97800 30880
rect 97640 30880 97800 31040
rect 97640 31040 97800 31200
rect 97640 31200 97800 31360
rect 97640 31360 97800 31520
rect 97640 31520 97800 31680
rect 97640 31680 97800 31840
rect 97640 31840 97800 32000
rect 97640 32000 97800 32160
rect 97640 32160 97800 32320
rect 97640 32320 97800 32480
rect 97640 32480 97800 32640
rect 97640 32640 97800 32800
rect 97640 32800 97800 32960
rect 97640 32960 97800 33120
rect 97640 33120 97800 33280
rect 97640 33280 97800 33440
rect 97640 33440 97800 33600
rect 97800 25600 97960 25760
rect 97800 25760 97960 25920
rect 97800 25920 97960 26080
rect 97800 26080 97960 26240
rect 97800 26240 97960 26400
rect 97800 26400 97960 26560
rect 97800 26560 97960 26720
rect 97800 26720 97960 26880
rect 97800 26880 97960 27040
rect 97800 27040 97960 27200
rect 97800 27200 97960 27360
rect 97800 27360 97960 27520
rect 97800 27520 97960 27680
rect 97800 27680 97960 27840
rect 97800 27840 97960 28000
rect 97800 28000 97960 28160
rect 97800 28160 97960 28320
rect 97800 28320 97960 28480
rect 97800 28480 97960 28640
rect 97800 28640 97960 28800
rect 97800 28800 97960 28960
rect 97800 28960 97960 29120
rect 97800 29120 97960 29280
rect 97800 29280 97960 29440
rect 97800 29440 97960 29600
rect 97800 29600 97960 29760
rect 97800 29760 97960 29920
rect 97800 29920 97960 30080
rect 97800 30080 97960 30240
rect 97800 30240 97960 30400
rect 97800 30400 97960 30560
rect 97800 30560 97960 30720
rect 97800 30720 97960 30880
rect 97800 30880 97960 31040
rect 97800 31040 97960 31200
rect 97800 31200 97960 31360
rect 97800 31360 97960 31520
rect 97800 31520 97960 31680
rect 97800 31680 97960 31840
rect 97800 31840 97960 32000
rect 97800 32000 97960 32160
rect 97800 32160 97960 32320
rect 97800 32320 97960 32480
rect 97800 32480 97960 32640
rect 97800 32640 97960 32800
rect 97800 32800 97960 32960
rect 97800 32960 97960 33120
rect 97800 33120 97960 33280
rect 97800 33280 97960 33440
rect 97800 33440 97960 33600
rect 97960 25760 98120 25920
rect 97960 25920 98120 26080
rect 97960 26080 98120 26240
rect 97960 26240 98120 26400
rect 97960 26400 98120 26560
rect 97960 26560 98120 26720
rect 97960 26720 98120 26880
rect 97960 26880 98120 27040
rect 97960 27040 98120 27200
rect 97960 27200 98120 27360
rect 97960 27360 98120 27520
rect 97960 27520 98120 27680
rect 97960 27680 98120 27840
rect 97960 27840 98120 28000
rect 97960 28000 98120 28160
rect 97960 28160 98120 28320
rect 97960 28320 98120 28480
rect 97960 28480 98120 28640
rect 97960 28640 98120 28800
rect 97960 28800 98120 28960
rect 97960 28960 98120 29120
rect 97960 29120 98120 29280
rect 97960 29280 98120 29440
rect 97960 29440 98120 29600
rect 97960 29600 98120 29760
rect 97960 29760 98120 29920
rect 97960 29920 98120 30080
rect 97960 30080 98120 30240
rect 97960 30240 98120 30400
rect 97960 30400 98120 30560
rect 97960 30560 98120 30720
rect 97960 30720 98120 30880
rect 97960 30880 98120 31040
rect 97960 31040 98120 31200
rect 97960 31200 98120 31360
rect 97960 31360 98120 31520
rect 97960 31520 98120 31680
rect 97960 31680 98120 31840
rect 97960 31840 98120 32000
rect 97960 32000 98120 32160
rect 97960 32160 98120 32320
rect 97960 32320 98120 32480
rect 97960 32480 98120 32640
rect 97960 32640 98120 32800
rect 97960 32800 98120 32960
rect 97960 32960 98120 33120
rect 97960 33120 98120 33280
rect 97960 33280 98120 33440
rect 97960 33440 98120 33600
rect 98120 25760 98280 25920
rect 98120 25920 98280 26080
rect 98120 26080 98280 26240
rect 98120 26240 98280 26400
rect 98120 26400 98280 26560
rect 98120 26560 98280 26720
rect 98120 26720 98280 26880
rect 98120 26880 98280 27040
rect 98120 27040 98280 27200
rect 98120 27200 98280 27360
rect 98120 27360 98280 27520
rect 98120 27520 98280 27680
rect 98120 27680 98280 27840
rect 98120 27840 98280 28000
rect 98120 28000 98280 28160
rect 98120 28160 98280 28320
rect 98120 28320 98280 28480
rect 98120 28480 98280 28640
rect 98120 28640 98280 28800
rect 98120 28800 98280 28960
rect 98120 28960 98280 29120
rect 98120 29120 98280 29280
rect 98120 29280 98280 29440
rect 98120 29440 98280 29600
rect 98120 29600 98280 29760
rect 98120 29760 98280 29920
rect 98120 29920 98280 30080
rect 98120 30080 98280 30240
rect 98120 30240 98280 30400
rect 98120 30400 98280 30560
rect 98120 30560 98280 30720
rect 98120 30720 98280 30880
rect 98120 30880 98280 31040
rect 98120 31040 98280 31200
rect 98120 31200 98280 31360
rect 98120 31360 98280 31520
rect 98120 31520 98280 31680
rect 98120 31680 98280 31840
rect 98120 31840 98280 32000
rect 98120 32000 98280 32160
rect 98120 32160 98280 32320
rect 98120 32320 98280 32480
rect 98120 32480 98280 32640
rect 98120 32640 98280 32800
rect 98120 32800 98280 32960
rect 98120 32960 98280 33120
rect 98120 33120 98280 33280
rect 98120 33280 98280 33440
rect 98120 33440 98280 33600
rect 98120 33600 98280 33760
rect 98280 25920 98440 26080
rect 98280 26080 98440 26240
rect 98280 26240 98440 26400
rect 98280 26400 98440 26560
rect 98280 26560 98440 26720
rect 98280 26720 98440 26880
rect 98280 26880 98440 27040
rect 98280 27040 98440 27200
rect 98280 27200 98440 27360
rect 98280 27360 98440 27520
rect 98280 27520 98440 27680
rect 98280 27680 98440 27840
rect 98280 27840 98440 28000
rect 98280 28000 98440 28160
rect 98280 28160 98440 28320
rect 98280 28320 98440 28480
rect 98280 28480 98440 28640
rect 98280 28640 98440 28800
rect 98280 28800 98440 28960
rect 98280 28960 98440 29120
rect 98280 29120 98440 29280
rect 98280 29280 98440 29440
rect 98280 29440 98440 29600
rect 98280 29600 98440 29760
rect 98280 29760 98440 29920
rect 98280 29920 98440 30080
rect 98280 30080 98440 30240
rect 98280 30240 98440 30400
rect 98280 30400 98440 30560
rect 98280 30560 98440 30720
rect 98280 30720 98440 30880
rect 98280 30880 98440 31040
rect 98280 31040 98440 31200
rect 98280 31200 98440 31360
rect 98280 31360 98440 31520
rect 98280 31520 98440 31680
rect 98280 31680 98440 31840
rect 98280 31840 98440 32000
rect 98280 32000 98440 32160
rect 98280 32160 98440 32320
rect 98280 32320 98440 32480
rect 98280 32480 98440 32640
rect 98280 32640 98440 32800
rect 98280 32800 98440 32960
rect 98280 32960 98440 33120
rect 98280 33120 98440 33280
rect 98280 33280 98440 33440
rect 98280 33440 98440 33600
rect 98280 33600 98440 33760
rect 98440 26080 98600 26240
rect 98440 26240 98600 26400
rect 98440 26400 98600 26560
rect 98440 26560 98600 26720
rect 98440 26720 98600 26880
rect 98440 26880 98600 27040
rect 98440 27040 98600 27200
rect 98440 27200 98600 27360
rect 98440 27360 98600 27520
rect 98440 27520 98600 27680
rect 98440 27680 98600 27840
rect 98440 27840 98600 28000
rect 98440 28000 98600 28160
rect 98440 28160 98600 28320
rect 98440 28320 98600 28480
rect 98440 28480 98600 28640
rect 98440 28640 98600 28800
rect 98440 28800 98600 28960
rect 98440 28960 98600 29120
rect 98440 29120 98600 29280
rect 98440 29280 98600 29440
rect 98440 29440 98600 29600
rect 98440 29600 98600 29760
rect 98440 29760 98600 29920
rect 98440 29920 98600 30080
rect 98440 30080 98600 30240
rect 98440 30240 98600 30400
rect 98440 30400 98600 30560
rect 98440 30560 98600 30720
rect 98440 30720 98600 30880
rect 98440 30880 98600 31040
rect 98440 31040 98600 31200
rect 98440 31200 98600 31360
rect 98440 31360 98600 31520
rect 98440 31520 98600 31680
rect 98440 31680 98600 31840
rect 98440 31840 98600 32000
rect 98440 32000 98600 32160
rect 98440 32160 98600 32320
rect 98440 32320 98600 32480
rect 98440 32480 98600 32640
rect 98440 32640 98600 32800
rect 98440 32800 98600 32960
rect 98440 32960 98600 33120
rect 98440 33120 98600 33280
rect 98440 33280 98600 33440
rect 98440 33440 98600 33600
rect 98440 33600 98600 33760
rect 98440 33760 98600 33920
rect 98600 26080 98760 26240
rect 98600 26240 98760 26400
rect 98600 26400 98760 26560
rect 98600 26560 98760 26720
rect 98600 26720 98760 26880
rect 98600 26880 98760 27040
rect 98600 27040 98760 27200
rect 98600 27200 98760 27360
rect 98600 27360 98760 27520
rect 98600 27520 98760 27680
rect 98600 27680 98760 27840
rect 98600 27840 98760 28000
rect 98600 28000 98760 28160
rect 98600 28160 98760 28320
rect 98600 28320 98760 28480
rect 98600 28480 98760 28640
rect 98600 28640 98760 28800
rect 98600 28800 98760 28960
rect 98600 28960 98760 29120
rect 98600 29120 98760 29280
rect 98600 29280 98760 29440
rect 98600 29440 98760 29600
rect 98600 29600 98760 29760
rect 98600 29760 98760 29920
rect 98600 29920 98760 30080
rect 98600 30080 98760 30240
rect 98600 30240 98760 30400
rect 98600 30400 98760 30560
rect 98600 30560 98760 30720
rect 98600 30720 98760 30880
rect 98600 30880 98760 31040
rect 98600 31040 98760 31200
rect 98600 31200 98760 31360
rect 98600 31360 98760 31520
rect 98600 31520 98760 31680
rect 98600 31680 98760 31840
rect 98600 31840 98760 32000
rect 98600 32000 98760 32160
rect 98600 32160 98760 32320
rect 98600 32320 98760 32480
rect 98600 32480 98760 32640
rect 98600 32640 98760 32800
rect 98600 32800 98760 32960
rect 98600 32960 98760 33120
rect 98600 33120 98760 33280
rect 98600 33280 98760 33440
rect 98600 33440 98760 33600
rect 98600 33600 98760 33760
rect 98600 33760 98760 33920
rect 98600 33920 98760 34080
rect 98760 26240 98920 26400
rect 98760 26400 98920 26560
rect 98760 26560 98920 26720
rect 98760 26720 98920 26880
rect 98760 26880 98920 27040
rect 98760 27040 98920 27200
rect 98760 27200 98920 27360
rect 98760 27360 98920 27520
rect 98760 27520 98920 27680
rect 98760 27680 98920 27840
rect 98760 27840 98920 28000
rect 98760 28000 98920 28160
rect 98760 28160 98920 28320
rect 98760 28320 98920 28480
rect 98760 28480 98920 28640
rect 98760 28640 98920 28800
rect 98760 28800 98920 28960
rect 98760 28960 98920 29120
rect 98760 29120 98920 29280
rect 98760 29280 98920 29440
rect 98760 29440 98920 29600
rect 98760 29600 98920 29760
rect 98760 29760 98920 29920
rect 98760 29920 98920 30080
rect 98760 30080 98920 30240
rect 98760 30240 98920 30400
rect 98760 30400 98920 30560
rect 98760 30560 98920 30720
rect 98760 30720 98920 30880
rect 98760 30880 98920 31040
rect 98760 31040 98920 31200
rect 98760 31200 98920 31360
rect 98760 31360 98920 31520
rect 98760 31520 98920 31680
rect 98760 31680 98920 31840
rect 98760 31840 98920 32000
rect 98760 32000 98920 32160
rect 98760 32160 98920 32320
rect 98760 32320 98920 32480
rect 98760 32480 98920 32640
rect 98760 32640 98920 32800
rect 98760 32800 98920 32960
rect 98760 32960 98920 33120
rect 98760 33120 98920 33280
rect 98760 33280 98920 33440
rect 98760 33440 98920 33600
rect 98760 33600 98920 33760
rect 98760 33760 98920 33920
rect 98760 33920 98920 34080
rect 98760 34080 98920 34240
rect 98920 26400 99080 26560
rect 98920 26560 99080 26720
rect 98920 26720 99080 26880
rect 98920 26880 99080 27040
rect 98920 27040 99080 27200
rect 98920 27200 99080 27360
rect 98920 27360 99080 27520
rect 98920 27520 99080 27680
rect 98920 27680 99080 27840
rect 98920 27840 99080 28000
rect 98920 28000 99080 28160
rect 98920 28160 99080 28320
rect 98920 28320 99080 28480
rect 98920 28480 99080 28640
rect 98920 28640 99080 28800
rect 98920 28800 99080 28960
rect 98920 28960 99080 29120
rect 98920 29120 99080 29280
rect 98920 29280 99080 29440
rect 98920 29440 99080 29600
rect 98920 29600 99080 29760
rect 98920 29760 99080 29920
rect 98920 29920 99080 30080
rect 98920 30080 99080 30240
rect 98920 30240 99080 30400
rect 98920 30400 99080 30560
rect 98920 30560 99080 30720
rect 98920 30720 99080 30880
rect 98920 30880 99080 31040
rect 98920 31040 99080 31200
rect 98920 31200 99080 31360
rect 98920 31360 99080 31520
rect 98920 31520 99080 31680
rect 98920 31680 99080 31840
rect 98920 31840 99080 32000
rect 98920 32000 99080 32160
rect 98920 32160 99080 32320
rect 98920 32320 99080 32480
rect 98920 32480 99080 32640
rect 98920 32640 99080 32800
rect 98920 32800 99080 32960
rect 98920 32960 99080 33120
rect 98920 33120 99080 33280
rect 98920 33280 99080 33440
rect 98920 33440 99080 33600
rect 98920 33600 99080 33760
rect 98920 33760 99080 33920
rect 98920 33920 99080 34080
rect 98920 34080 99080 34240
rect 98920 34240 99080 34400
rect 99080 26560 99240 26720
rect 99080 26720 99240 26880
rect 99080 26880 99240 27040
rect 99080 27040 99240 27200
rect 99080 27200 99240 27360
rect 99080 27360 99240 27520
rect 99080 27520 99240 27680
rect 99080 27680 99240 27840
rect 99080 27840 99240 28000
rect 99080 28000 99240 28160
rect 99080 28160 99240 28320
rect 99080 28320 99240 28480
rect 99080 28480 99240 28640
rect 99080 28640 99240 28800
rect 99080 28800 99240 28960
rect 99080 28960 99240 29120
rect 99080 29120 99240 29280
rect 99080 29280 99240 29440
rect 99080 29440 99240 29600
rect 99080 29600 99240 29760
rect 99080 29760 99240 29920
rect 99080 29920 99240 30080
rect 99080 30080 99240 30240
rect 99080 30240 99240 30400
rect 99080 30400 99240 30560
rect 99080 30560 99240 30720
rect 99080 30720 99240 30880
rect 99080 30880 99240 31040
rect 99080 31040 99240 31200
rect 99080 31200 99240 31360
rect 99080 31360 99240 31520
rect 99080 31520 99240 31680
rect 99080 31680 99240 31840
rect 99080 31840 99240 32000
rect 99080 32000 99240 32160
rect 99080 32160 99240 32320
rect 99080 32320 99240 32480
rect 99080 32480 99240 32640
rect 99080 32640 99240 32800
rect 99080 32800 99240 32960
rect 99080 32960 99240 33120
rect 99080 33120 99240 33280
rect 99080 33280 99240 33440
rect 99080 33440 99240 33600
rect 99080 33600 99240 33760
rect 99080 33760 99240 33920
rect 99080 33920 99240 34080
rect 99080 34080 99240 34240
rect 99080 34240 99240 34400
rect 99080 34400 99240 34560
rect 99240 26720 99400 26880
rect 99240 26880 99400 27040
rect 99240 27040 99400 27200
rect 99240 27200 99400 27360
rect 99240 27360 99400 27520
rect 99240 27520 99400 27680
rect 99240 27680 99400 27840
rect 99240 27840 99400 28000
rect 99240 28000 99400 28160
rect 99240 28160 99400 28320
rect 99240 28320 99400 28480
rect 99240 28480 99400 28640
rect 99240 28640 99400 28800
rect 99240 28800 99400 28960
rect 99240 28960 99400 29120
rect 99240 29120 99400 29280
rect 99240 29280 99400 29440
rect 99240 29440 99400 29600
rect 99240 29600 99400 29760
rect 99240 29760 99400 29920
rect 99240 29920 99400 30080
rect 99240 30080 99400 30240
rect 99240 30240 99400 30400
rect 99240 30400 99400 30560
rect 99240 30560 99400 30720
rect 99240 30720 99400 30880
rect 99240 30880 99400 31040
rect 99240 31040 99400 31200
rect 99240 31200 99400 31360
rect 99240 31360 99400 31520
rect 99240 31520 99400 31680
rect 99240 31680 99400 31840
rect 99240 31840 99400 32000
rect 99240 32000 99400 32160
rect 99240 32160 99400 32320
rect 99240 32320 99400 32480
rect 99240 32480 99400 32640
rect 99240 32640 99400 32800
rect 99240 32800 99400 32960
rect 99240 32960 99400 33120
rect 99240 33120 99400 33280
rect 99240 33280 99400 33440
rect 99240 33440 99400 33600
rect 99240 33600 99400 33760
rect 99240 33760 99400 33920
rect 99240 33920 99400 34080
rect 99240 34080 99400 34240
rect 99240 34240 99400 34400
rect 99240 34400 99400 34560
rect 99240 34560 99400 34720
rect 99400 26880 99560 27040
rect 99400 27040 99560 27200
rect 99400 27200 99560 27360
rect 99400 27360 99560 27520
rect 99400 27520 99560 27680
rect 99400 27680 99560 27840
rect 99400 27840 99560 28000
rect 99400 28000 99560 28160
rect 99400 28160 99560 28320
rect 99400 28320 99560 28480
rect 99400 28480 99560 28640
rect 99400 28640 99560 28800
rect 99400 28800 99560 28960
rect 99400 28960 99560 29120
rect 99400 29120 99560 29280
rect 99400 29280 99560 29440
rect 99400 29440 99560 29600
rect 99400 29600 99560 29760
rect 99400 29760 99560 29920
rect 99400 29920 99560 30080
rect 99400 30080 99560 30240
rect 99400 30240 99560 30400
rect 99400 30400 99560 30560
rect 99400 30560 99560 30720
rect 99400 30720 99560 30880
rect 99400 30880 99560 31040
rect 99400 31040 99560 31200
rect 99400 31200 99560 31360
rect 99400 31360 99560 31520
rect 99400 31520 99560 31680
rect 99400 31680 99560 31840
rect 99400 31840 99560 32000
rect 99400 32000 99560 32160
rect 99400 32160 99560 32320
rect 99400 32320 99560 32480
rect 99400 32480 99560 32640
rect 99400 32640 99560 32800
rect 99400 32800 99560 32960
rect 99400 32960 99560 33120
rect 99400 33120 99560 33280
rect 99400 33280 99560 33440
rect 99400 33440 99560 33600
rect 99400 33600 99560 33760
rect 99400 33760 99560 33920
rect 99400 33920 99560 34080
rect 99400 34080 99560 34240
rect 99400 34240 99560 34400
rect 99400 34400 99560 34560
rect 99400 34560 99560 34720
rect 99400 34720 99560 34880
rect 99560 27040 99720 27200
rect 99560 27200 99720 27360
rect 99560 27360 99720 27520
rect 99560 27520 99720 27680
rect 99560 27680 99720 27840
rect 99560 27840 99720 28000
rect 99560 28000 99720 28160
rect 99560 28160 99720 28320
rect 99560 28320 99720 28480
rect 99560 28480 99720 28640
rect 99560 28640 99720 28800
rect 99560 28800 99720 28960
rect 99560 28960 99720 29120
rect 99560 29120 99720 29280
rect 99560 29280 99720 29440
rect 99560 29440 99720 29600
rect 99560 29600 99720 29760
rect 99560 29760 99720 29920
rect 99560 29920 99720 30080
rect 99560 30080 99720 30240
rect 99560 30240 99720 30400
rect 99560 30400 99720 30560
rect 99560 30560 99720 30720
rect 99560 30720 99720 30880
rect 99560 30880 99720 31040
rect 99560 31040 99720 31200
rect 99560 31200 99720 31360
rect 99560 31360 99720 31520
rect 99560 31520 99720 31680
rect 99560 31680 99720 31840
rect 99560 31840 99720 32000
rect 99560 32000 99720 32160
rect 99560 32160 99720 32320
rect 99560 32320 99720 32480
rect 99560 32480 99720 32640
rect 99560 32640 99720 32800
rect 99560 32800 99720 32960
rect 99560 32960 99720 33120
rect 99560 33120 99720 33280
rect 99560 33280 99720 33440
rect 99560 33440 99720 33600
rect 99560 33600 99720 33760
rect 99560 33760 99720 33920
rect 99560 33920 99720 34080
rect 99560 34080 99720 34240
rect 99560 34240 99720 34400
rect 99560 34400 99720 34560
rect 99560 34560 99720 34720
rect 99560 34720 99720 34880
rect 99560 34880 99720 35040
rect 99720 27200 99880 27360
rect 99720 27360 99880 27520
rect 99720 27520 99880 27680
rect 99720 27680 99880 27840
rect 99720 27840 99880 28000
rect 99720 28000 99880 28160
rect 99720 28160 99880 28320
rect 99720 28320 99880 28480
rect 99720 28480 99880 28640
rect 99720 28640 99880 28800
rect 99720 28800 99880 28960
rect 99720 28960 99880 29120
rect 99720 29120 99880 29280
rect 99720 29280 99880 29440
rect 99720 29440 99880 29600
rect 99720 29600 99880 29760
rect 99720 29760 99880 29920
rect 99720 29920 99880 30080
rect 99720 30080 99880 30240
rect 99720 30240 99880 30400
rect 99720 30400 99880 30560
rect 99720 30560 99880 30720
rect 99720 30720 99880 30880
rect 99720 30880 99880 31040
rect 99720 31040 99880 31200
rect 99720 31200 99880 31360
rect 99720 31360 99880 31520
rect 99720 31520 99880 31680
rect 99720 31680 99880 31840
rect 99720 31840 99880 32000
rect 99720 32000 99880 32160
rect 99720 32160 99880 32320
rect 99720 32320 99880 32480
rect 99720 32480 99880 32640
rect 99720 32640 99880 32800
rect 99720 32800 99880 32960
rect 99720 32960 99880 33120
rect 99720 33120 99880 33280
rect 99720 33280 99880 33440
rect 99720 33440 99880 33600
rect 99720 33600 99880 33760
rect 99720 33760 99880 33920
rect 99720 33920 99880 34080
rect 99720 34080 99880 34240
rect 99720 34240 99880 34400
rect 99720 34400 99880 34560
rect 99720 34560 99880 34720
rect 99720 34720 99880 34880
rect 99720 34880 99880 35040
rect 99720 35040 99880 35200
rect 99880 27520 100040 27680
rect 99880 27680 100040 27840
rect 99880 27840 100040 28000
rect 99880 28000 100040 28160
rect 99880 28160 100040 28320
rect 99880 28320 100040 28480
rect 99880 28480 100040 28640
rect 99880 28640 100040 28800
rect 99880 28800 100040 28960
rect 99880 28960 100040 29120
rect 99880 29120 100040 29280
rect 99880 29280 100040 29440
rect 99880 29440 100040 29600
rect 99880 29600 100040 29760
rect 99880 29760 100040 29920
rect 99880 29920 100040 30080
rect 99880 30080 100040 30240
rect 99880 30240 100040 30400
rect 99880 30400 100040 30560
rect 99880 30560 100040 30720
rect 99880 30720 100040 30880
rect 99880 30880 100040 31040
rect 99880 31040 100040 31200
rect 99880 31200 100040 31360
rect 99880 31360 100040 31520
rect 99880 31520 100040 31680
rect 99880 31680 100040 31840
rect 99880 31840 100040 32000
rect 99880 32000 100040 32160
rect 99880 32160 100040 32320
rect 99880 32320 100040 32480
rect 99880 32480 100040 32640
rect 99880 32640 100040 32800
rect 99880 32800 100040 32960
rect 99880 32960 100040 33120
rect 99880 33120 100040 33280
rect 99880 33280 100040 33440
rect 99880 33440 100040 33600
rect 99880 33600 100040 33760
rect 99880 33760 100040 33920
rect 99880 33920 100040 34080
rect 99880 34080 100040 34240
rect 99880 34240 100040 34400
rect 99880 34400 100040 34560
rect 99880 34560 100040 34720
rect 99880 34720 100040 34880
rect 99880 34880 100040 35040
rect 99880 35040 100040 35200
rect 99880 35200 100040 35360
rect 100040 27680 100200 27840
rect 100040 27840 100200 28000
rect 100040 28000 100200 28160
rect 100040 28160 100200 28320
rect 100040 28320 100200 28480
rect 100040 28480 100200 28640
rect 100040 28640 100200 28800
rect 100040 28800 100200 28960
rect 100040 28960 100200 29120
rect 100040 29120 100200 29280
rect 100040 29280 100200 29440
rect 100040 29440 100200 29600
rect 100040 29600 100200 29760
rect 100040 29760 100200 29920
rect 100040 29920 100200 30080
rect 100040 30080 100200 30240
rect 100040 30240 100200 30400
rect 100040 30400 100200 30560
rect 100040 30560 100200 30720
rect 100040 30720 100200 30880
rect 100040 30880 100200 31040
rect 100040 31040 100200 31200
rect 100040 31200 100200 31360
rect 100040 31360 100200 31520
rect 100040 31520 100200 31680
rect 100040 31680 100200 31840
rect 100040 31840 100200 32000
rect 100040 32000 100200 32160
rect 100040 32160 100200 32320
rect 100040 32320 100200 32480
rect 100040 32480 100200 32640
rect 100040 32640 100200 32800
rect 100040 32800 100200 32960
rect 100040 32960 100200 33120
rect 100040 33120 100200 33280
rect 100040 33280 100200 33440
rect 100040 33440 100200 33600
rect 100040 33600 100200 33760
rect 100040 33760 100200 33920
rect 100040 33920 100200 34080
rect 100040 34080 100200 34240
rect 100040 34240 100200 34400
rect 100040 34400 100200 34560
rect 100040 34560 100200 34720
rect 100040 34720 100200 34880
rect 100040 34880 100200 35040
rect 100040 35040 100200 35200
rect 100040 35200 100200 35360
rect 100040 35360 100200 35520
rect 100200 28000 100360 28160
rect 100200 28160 100360 28320
rect 100200 28320 100360 28480
rect 100200 28480 100360 28640
rect 100200 28640 100360 28800
rect 100200 28800 100360 28960
rect 100200 28960 100360 29120
rect 100200 29120 100360 29280
rect 100200 29280 100360 29440
rect 100200 29440 100360 29600
rect 100200 29600 100360 29760
rect 100200 29760 100360 29920
rect 100200 29920 100360 30080
rect 100200 30080 100360 30240
rect 100200 30240 100360 30400
rect 100200 30400 100360 30560
rect 100200 30560 100360 30720
rect 100200 30720 100360 30880
rect 100200 30880 100360 31040
rect 100200 31040 100360 31200
rect 100200 31200 100360 31360
rect 100200 31360 100360 31520
rect 100200 31520 100360 31680
rect 100200 31680 100360 31840
rect 100200 31840 100360 32000
rect 100200 32000 100360 32160
rect 100200 32160 100360 32320
rect 100200 32320 100360 32480
rect 100200 32480 100360 32640
rect 100200 32640 100360 32800
rect 100200 32800 100360 32960
rect 100200 32960 100360 33120
rect 100200 33120 100360 33280
rect 100200 33280 100360 33440
rect 100200 33440 100360 33600
rect 100200 33600 100360 33760
rect 100200 33760 100360 33920
rect 100200 33920 100360 34080
rect 100200 34080 100360 34240
rect 100200 34240 100360 34400
rect 100200 34400 100360 34560
rect 100200 34560 100360 34720
rect 100200 34720 100360 34880
rect 100200 34880 100360 35040
rect 100200 35040 100360 35200
rect 100200 35200 100360 35360
rect 100200 35360 100360 35520
rect 100200 35520 100360 35680
rect 100360 28320 100520 28480
rect 100360 28480 100520 28640
rect 100360 28640 100520 28800
rect 100360 28800 100520 28960
rect 100360 28960 100520 29120
rect 100360 29120 100520 29280
rect 100360 29280 100520 29440
rect 100360 29440 100520 29600
rect 100360 29600 100520 29760
rect 100360 29760 100520 29920
rect 100360 29920 100520 30080
rect 100360 30080 100520 30240
rect 100360 30240 100520 30400
rect 100360 30400 100520 30560
rect 100360 30560 100520 30720
rect 100360 30720 100520 30880
rect 100360 30880 100520 31040
rect 100360 31040 100520 31200
rect 100360 31200 100520 31360
rect 100360 31360 100520 31520
rect 100360 31520 100520 31680
rect 100360 31680 100520 31840
rect 100360 31840 100520 32000
rect 100360 32000 100520 32160
rect 100360 32160 100520 32320
rect 100360 32320 100520 32480
rect 100360 32480 100520 32640
rect 100360 32640 100520 32800
rect 100360 32800 100520 32960
rect 100360 32960 100520 33120
rect 100360 33120 100520 33280
rect 100360 33280 100520 33440
rect 100360 33440 100520 33600
rect 100360 33600 100520 33760
rect 100360 33760 100520 33920
rect 100360 33920 100520 34080
rect 100360 34080 100520 34240
rect 100360 34240 100520 34400
rect 100360 34400 100520 34560
rect 100360 34560 100520 34720
rect 100360 34720 100520 34880
rect 100360 34880 100520 35040
rect 100360 35040 100520 35200
rect 100360 35200 100520 35360
rect 100360 35360 100520 35520
rect 100360 35520 100520 35680
rect 100360 35680 100520 35840
rect 100520 28960 100680 29120
rect 100520 29120 100680 29280
rect 100520 29280 100680 29440
rect 100520 29440 100680 29600
rect 100520 29600 100680 29760
rect 100520 29760 100680 29920
rect 100520 29920 100680 30080
rect 100520 30080 100680 30240
rect 100520 30240 100680 30400
rect 100520 30400 100680 30560
rect 100520 30560 100680 30720
rect 100520 31520 100680 31680
rect 100520 31680 100680 31840
rect 100520 31840 100680 32000
rect 100520 32000 100680 32160
rect 100520 32160 100680 32320
rect 100520 32320 100680 32480
rect 100520 32480 100680 32640
rect 100520 32640 100680 32800
rect 100520 32800 100680 32960
rect 100520 32960 100680 33120
rect 100520 33120 100680 33280
rect 100520 33280 100680 33440
rect 100520 33440 100680 33600
rect 100520 33600 100680 33760
rect 100520 33760 100680 33920
rect 100520 33920 100680 34080
rect 100520 34080 100680 34240
rect 100520 34240 100680 34400
rect 100520 34400 100680 34560
rect 100520 34560 100680 34720
rect 100520 34720 100680 34880
rect 100520 34880 100680 35040
rect 100520 35040 100680 35200
rect 100520 35200 100680 35360
rect 100520 35360 100680 35520
rect 100520 35520 100680 35680
rect 100520 35680 100680 35840
rect 100520 35840 100680 36000
rect 100520 48960 100680 49120
rect 100520 49120 100680 49280
rect 100520 49280 100680 49440
rect 100520 49440 100680 49600
rect 100520 49600 100680 49760
rect 100520 49760 100680 49920
rect 100520 49920 100680 50080
rect 100520 50080 100680 50240
rect 100520 50240 100680 50400
rect 100680 31840 100840 32000
rect 100680 32000 100840 32160
rect 100680 32160 100840 32320
rect 100680 32320 100840 32480
rect 100680 32480 100840 32640
rect 100680 32640 100840 32800
rect 100680 32800 100840 32960
rect 100680 32960 100840 33120
rect 100680 33120 100840 33280
rect 100680 33280 100840 33440
rect 100680 33440 100840 33600
rect 100680 33600 100840 33760
rect 100680 33760 100840 33920
rect 100680 33920 100840 34080
rect 100680 34080 100840 34240
rect 100680 34240 100840 34400
rect 100680 34400 100840 34560
rect 100680 34560 100840 34720
rect 100680 34720 100840 34880
rect 100680 34880 100840 35040
rect 100680 35040 100840 35200
rect 100680 35200 100840 35360
rect 100680 35360 100840 35520
rect 100680 35520 100840 35680
rect 100680 35680 100840 35840
rect 100680 35840 100840 36000
rect 100680 48320 100840 48480
rect 100680 48480 100840 48640
rect 100680 48640 100840 48800
rect 100680 48800 100840 48960
rect 100680 48960 100840 49120
rect 100680 49120 100840 49280
rect 100680 49280 100840 49440
rect 100680 49440 100840 49600
rect 100680 49600 100840 49760
rect 100680 49760 100840 49920
rect 100680 49920 100840 50080
rect 100680 50080 100840 50240
rect 100680 50240 100840 50400
rect 100680 50400 100840 50560
rect 100680 50560 100840 50720
rect 100680 50720 100840 50880
rect 100680 50880 100840 51040
rect 100840 32160 101000 32320
rect 100840 32320 101000 32480
rect 100840 32480 101000 32640
rect 100840 32640 101000 32800
rect 100840 32800 101000 32960
rect 100840 32960 101000 33120
rect 100840 33120 101000 33280
rect 100840 33280 101000 33440
rect 100840 33440 101000 33600
rect 100840 33600 101000 33760
rect 100840 33760 101000 33920
rect 100840 33920 101000 34080
rect 100840 34080 101000 34240
rect 100840 34240 101000 34400
rect 100840 34400 101000 34560
rect 100840 34560 101000 34720
rect 100840 34720 101000 34880
rect 100840 34880 101000 35040
rect 100840 35040 101000 35200
rect 100840 35200 101000 35360
rect 100840 35360 101000 35520
rect 100840 35520 101000 35680
rect 100840 35680 101000 35840
rect 100840 35840 101000 36000
rect 100840 36000 101000 36160
rect 100840 48000 101000 48160
rect 100840 48160 101000 48320
rect 100840 48320 101000 48480
rect 100840 48480 101000 48640
rect 100840 48640 101000 48800
rect 100840 48800 101000 48960
rect 100840 48960 101000 49120
rect 100840 49120 101000 49280
rect 100840 49280 101000 49440
rect 100840 49440 101000 49600
rect 100840 49600 101000 49760
rect 100840 49760 101000 49920
rect 100840 49920 101000 50080
rect 100840 50080 101000 50240
rect 100840 50240 101000 50400
rect 100840 50400 101000 50560
rect 100840 50560 101000 50720
rect 100840 50720 101000 50880
rect 100840 50880 101000 51040
rect 100840 51040 101000 51200
rect 100840 51200 101000 51360
rect 101000 32320 101160 32480
rect 101000 32480 101160 32640
rect 101000 32640 101160 32800
rect 101000 32800 101160 32960
rect 101000 32960 101160 33120
rect 101000 33120 101160 33280
rect 101000 33280 101160 33440
rect 101000 33440 101160 33600
rect 101000 33600 101160 33760
rect 101000 33760 101160 33920
rect 101000 33920 101160 34080
rect 101000 34080 101160 34240
rect 101000 34240 101160 34400
rect 101000 34400 101160 34560
rect 101000 34560 101160 34720
rect 101000 34720 101160 34880
rect 101000 34880 101160 35040
rect 101000 35040 101160 35200
rect 101000 35200 101160 35360
rect 101000 35360 101160 35520
rect 101000 35520 101160 35680
rect 101000 35680 101160 35840
rect 101000 35840 101160 36000
rect 101000 36000 101160 36160
rect 101000 36160 101160 36320
rect 101000 47680 101160 47840
rect 101000 47840 101160 48000
rect 101000 48000 101160 48160
rect 101000 48160 101160 48320
rect 101000 48320 101160 48480
rect 101000 48480 101160 48640
rect 101000 48640 101160 48800
rect 101000 48800 101160 48960
rect 101000 48960 101160 49120
rect 101000 49120 101160 49280
rect 101000 49280 101160 49440
rect 101000 49440 101160 49600
rect 101000 49600 101160 49760
rect 101000 49760 101160 49920
rect 101000 49920 101160 50080
rect 101000 50080 101160 50240
rect 101000 50240 101160 50400
rect 101000 50400 101160 50560
rect 101000 50560 101160 50720
rect 101000 50720 101160 50880
rect 101000 50880 101160 51040
rect 101000 51040 101160 51200
rect 101000 51200 101160 51360
rect 101000 51360 101160 51520
rect 101000 51520 101160 51680
rect 101160 32480 101320 32640
rect 101160 32640 101320 32800
rect 101160 32800 101320 32960
rect 101160 32960 101320 33120
rect 101160 33120 101320 33280
rect 101160 33280 101320 33440
rect 101160 33440 101320 33600
rect 101160 33600 101320 33760
rect 101160 33760 101320 33920
rect 101160 33920 101320 34080
rect 101160 34080 101320 34240
rect 101160 34240 101320 34400
rect 101160 34400 101320 34560
rect 101160 34560 101320 34720
rect 101160 34720 101320 34880
rect 101160 34880 101320 35040
rect 101160 35040 101320 35200
rect 101160 35200 101320 35360
rect 101160 35360 101320 35520
rect 101160 35520 101320 35680
rect 101160 35680 101320 35840
rect 101160 35840 101320 36000
rect 101160 36000 101320 36160
rect 101160 36160 101320 36320
rect 101160 36320 101320 36480
rect 101160 47520 101320 47680
rect 101160 47680 101320 47840
rect 101160 47840 101320 48000
rect 101160 48000 101320 48160
rect 101160 48160 101320 48320
rect 101160 48320 101320 48480
rect 101160 48480 101320 48640
rect 101160 48640 101320 48800
rect 101160 48800 101320 48960
rect 101160 48960 101320 49120
rect 101160 49120 101320 49280
rect 101160 49280 101320 49440
rect 101160 49440 101320 49600
rect 101160 49600 101320 49760
rect 101160 49760 101320 49920
rect 101160 49920 101320 50080
rect 101160 50080 101320 50240
rect 101160 50240 101320 50400
rect 101160 50400 101320 50560
rect 101160 50560 101320 50720
rect 101160 50720 101320 50880
rect 101160 50880 101320 51040
rect 101160 51040 101320 51200
rect 101160 51200 101320 51360
rect 101160 51360 101320 51520
rect 101160 51520 101320 51680
rect 101160 51680 101320 51840
rect 101320 32800 101480 32960
rect 101320 32960 101480 33120
rect 101320 33120 101480 33280
rect 101320 33280 101480 33440
rect 101320 33440 101480 33600
rect 101320 33600 101480 33760
rect 101320 33760 101480 33920
rect 101320 33920 101480 34080
rect 101320 34080 101480 34240
rect 101320 34240 101480 34400
rect 101320 34400 101480 34560
rect 101320 34560 101480 34720
rect 101320 34720 101480 34880
rect 101320 34880 101480 35040
rect 101320 35040 101480 35200
rect 101320 35200 101480 35360
rect 101320 35360 101480 35520
rect 101320 35520 101480 35680
rect 101320 35680 101480 35840
rect 101320 35840 101480 36000
rect 101320 36000 101480 36160
rect 101320 36160 101480 36320
rect 101320 36320 101480 36480
rect 101320 36480 101480 36640
rect 101320 47200 101480 47360
rect 101320 47360 101480 47520
rect 101320 47520 101480 47680
rect 101320 47680 101480 47840
rect 101320 47840 101480 48000
rect 101320 48000 101480 48160
rect 101320 48160 101480 48320
rect 101320 48320 101480 48480
rect 101320 48480 101480 48640
rect 101320 48640 101480 48800
rect 101320 48800 101480 48960
rect 101320 48960 101480 49120
rect 101320 49120 101480 49280
rect 101320 49280 101480 49440
rect 101320 49440 101480 49600
rect 101320 49600 101480 49760
rect 101320 49760 101480 49920
rect 101320 49920 101480 50080
rect 101320 50080 101480 50240
rect 101320 50240 101480 50400
rect 101320 50400 101480 50560
rect 101320 50560 101480 50720
rect 101320 50720 101480 50880
rect 101320 50880 101480 51040
rect 101320 51040 101480 51200
rect 101320 51200 101480 51360
rect 101320 51360 101480 51520
rect 101320 51520 101480 51680
rect 101320 51680 101480 51840
rect 101320 51840 101480 52000
rect 101480 32960 101640 33120
rect 101480 33120 101640 33280
rect 101480 33280 101640 33440
rect 101480 33440 101640 33600
rect 101480 33600 101640 33760
rect 101480 33760 101640 33920
rect 101480 33920 101640 34080
rect 101480 34080 101640 34240
rect 101480 34240 101640 34400
rect 101480 34400 101640 34560
rect 101480 34560 101640 34720
rect 101480 34720 101640 34880
rect 101480 34880 101640 35040
rect 101480 35040 101640 35200
rect 101480 35200 101640 35360
rect 101480 35360 101640 35520
rect 101480 35520 101640 35680
rect 101480 35680 101640 35840
rect 101480 35840 101640 36000
rect 101480 36000 101640 36160
rect 101480 36160 101640 36320
rect 101480 36320 101640 36480
rect 101480 36480 101640 36640
rect 101480 36640 101640 36800
rect 101480 47040 101640 47200
rect 101480 47200 101640 47360
rect 101480 47360 101640 47520
rect 101480 47520 101640 47680
rect 101480 47680 101640 47840
rect 101480 47840 101640 48000
rect 101480 48000 101640 48160
rect 101480 48160 101640 48320
rect 101480 48320 101640 48480
rect 101480 48480 101640 48640
rect 101480 48640 101640 48800
rect 101480 48800 101640 48960
rect 101480 48960 101640 49120
rect 101480 49120 101640 49280
rect 101480 49280 101640 49440
rect 101480 49440 101640 49600
rect 101480 49600 101640 49760
rect 101480 49760 101640 49920
rect 101480 49920 101640 50080
rect 101480 50080 101640 50240
rect 101480 50240 101640 50400
rect 101480 50400 101640 50560
rect 101480 50560 101640 50720
rect 101480 50720 101640 50880
rect 101480 50880 101640 51040
rect 101480 51040 101640 51200
rect 101480 51200 101640 51360
rect 101480 51360 101640 51520
rect 101480 51520 101640 51680
rect 101480 51680 101640 51840
rect 101480 51840 101640 52000
rect 101480 52000 101640 52160
rect 101640 33120 101800 33280
rect 101640 33280 101800 33440
rect 101640 33440 101800 33600
rect 101640 33600 101800 33760
rect 101640 33760 101800 33920
rect 101640 33920 101800 34080
rect 101640 34080 101800 34240
rect 101640 34240 101800 34400
rect 101640 34400 101800 34560
rect 101640 34560 101800 34720
rect 101640 34720 101800 34880
rect 101640 34880 101800 35040
rect 101640 35040 101800 35200
rect 101640 35200 101800 35360
rect 101640 35360 101800 35520
rect 101640 35520 101800 35680
rect 101640 35680 101800 35840
rect 101640 35840 101800 36000
rect 101640 36000 101800 36160
rect 101640 36160 101800 36320
rect 101640 36320 101800 36480
rect 101640 36480 101800 36640
rect 101640 36640 101800 36800
rect 101640 36800 101800 36960
rect 101640 46880 101800 47040
rect 101640 47040 101800 47200
rect 101640 47200 101800 47360
rect 101640 47360 101800 47520
rect 101640 47520 101800 47680
rect 101640 47680 101800 47840
rect 101640 47840 101800 48000
rect 101640 48000 101800 48160
rect 101640 48160 101800 48320
rect 101640 48320 101800 48480
rect 101640 48480 101800 48640
rect 101640 48640 101800 48800
rect 101640 48800 101800 48960
rect 101640 48960 101800 49120
rect 101640 49120 101800 49280
rect 101640 49280 101800 49440
rect 101640 49440 101800 49600
rect 101640 49600 101800 49760
rect 101640 49760 101800 49920
rect 101640 49920 101800 50080
rect 101640 50080 101800 50240
rect 101640 50240 101800 50400
rect 101640 50400 101800 50560
rect 101640 50560 101800 50720
rect 101640 50720 101800 50880
rect 101640 50880 101800 51040
rect 101640 51040 101800 51200
rect 101640 51200 101800 51360
rect 101640 51360 101800 51520
rect 101640 51520 101800 51680
rect 101640 51680 101800 51840
rect 101640 51840 101800 52000
rect 101640 52000 101800 52160
rect 101640 52160 101800 52320
rect 101800 33440 101960 33600
rect 101800 33600 101960 33760
rect 101800 33760 101960 33920
rect 101800 33920 101960 34080
rect 101800 34080 101960 34240
rect 101800 34240 101960 34400
rect 101800 34400 101960 34560
rect 101800 34560 101960 34720
rect 101800 34720 101960 34880
rect 101800 34880 101960 35040
rect 101800 35040 101960 35200
rect 101800 35200 101960 35360
rect 101800 35360 101960 35520
rect 101800 35520 101960 35680
rect 101800 35680 101960 35840
rect 101800 35840 101960 36000
rect 101800 36000 101960 36160
rect 101800 36160 101960 36320
rect 101800 36320 101960 36480
rect 101800 36480 101960 36640
rect 101800 36640 101960 36800
rect 101800 36800 101960 36960
rect 101800 36960 101960 37120
rect 101800 46720 101960 46880
rect 101800 46880 101960 47040
rect 101800 47040 101960 47200
rect 101800 47200 101960 47360
rect 101800 47360 101960 47520
rect 101800 47520 101960 47680
rect 101800 47680 101960 47840
rect 101800 47840 101960 48000
rect 101800 48000 101960 48160
rect 101800 48160 101960 48320
rect 101800 48320 101960 48480
rect 101800 48480 101960 48640
rect 101800 48640 101960 48800
rect 101800 48800 101960 48960
rect 101800 48960 101960 49120
rect 101800 49120 101960 49280
rect 101800 49280 101960 49440
rect 101800 49440 101960 49600
rect 101800 49600 101960 49760
rect 101800 49760 101960 49920
rect 101800 49920 101960 50080
rect 101800 50080 101960 50240
rect 101800 50240 101960 50400
rect 101800 50400 101960 50560
rect 101800 50560 101960 50720
rect 101800 50720 101960 50880
rect 101800 50880 101960 51040
rect 101800 51040 101960 51200
rect 101800 51200 101960 51360
rect 101800 51360 101960 51520
rect 101800 51520 101960 51680
rect 101800 51680 101960 51840
rect 101800 51840 101960 52000
rect 101800 52000 101960 52160
rect 101800 52160 101960 52320
rect 101800 52320 101960 52480
rect 101960 33600 102120 33760
rect 101960 33760 102120 33920
rect 101960 33920 102120 34080
rect 101960 34080 102120 34240
rect 101960 34240 102120 34400
rect 101960 34400 102120 34560
rect 101960 34560 102120 34720
rect 101960 34720 102120 34880
rect 101960 34880 102120 35040
rect 101960 35040 102120 35200
rect 101960 35200 102120 35360
rect 101960 35360 102120 35520
rect 101960 35520 102120 35680
rect 101960 35680 102120 35840
rect 101960 35840 102120 36000
rect 101960 36000 102120 36160
rect 101960 36160 102120 36320
rect 101960 36320 102120 36480
rect 101960 36480 102120 36640
rect 101960 36640 102120 36800
rect 101960 36800 102120 36960
rect 101960 36960 102120 37120
rect 101960 37120 102120 37280
rect 101960 46560 102120 46720
rect 101960 46720 102120 46880
rect 101960 46880 102120 47040
rect 101960 47040 102120 47200
rect 101960 47200 102120 47360
rect 101960 47360 102120 47520
rect 101960 47520 102120 47680
rect 101960 47680 102120 47840
rect 101960 47840 102120 48000
rect 101960 48000 102120 48160
rect 101960 48160 102120 48320
rect 101960 48320 102120 48480
rect 101960 48480 102120 48640
rect 101960 48640 102120 48800
rect 101960 48800 102120 48960
rect 101960 48960 102120 49120
rect 101960 49120 102120 49280
rect 101960 49280 102120 49440
rect 101960 49440 102120 49600
rect 101960 49600 102120 49760
rect 101960 49760 102120 49920
rect 101960 49920 102120 50080
rect 101960 50080 102120 50240
rect 101960 50240 102120 50400
rect 101960 50400 102120 50560
rect 101960 50560 102120 50720
rect 101960 50720 102120 50880
rect 101960 50880 102120 51040
rect 101960 51040 102120 51200
rect 101960 51200 102120 51360
rect 101960 51360 102120 51520
rect 101960 51520 102120 51680
rect 101960 51680 102120 51840
rect 101960 51840 102120 52000
rect 101960 52000 102120 52160
rect 101960 52160 102120 52320
rect 101960 52320 102120 52480
rect 101960 52480 102120 52640
rect 102120 33760 102280 33920
rect 102120 33920 102280 34080
rect 102120 34080 102280 34240
rect 102120 34240 102280 34400
rect 102120 34400 102280 34560
rect 102120 34560 102280 34720
rect 102120 34720 102280 34880
rect 102120 34880 102280 35040
rect 102120 35040 102280 35200
rect 102120 35200 102280 35360
rect 102120 35360 102280 35520
rect 102120 35520 102280 35680
rect 102120 35680 102280 35840
rect 102120 35840 102280 36000
rect 102120 36000 102280 36160
rect 102120 36160 102280 36320
rect 102120 36320 102280 36480
rect 102120 36480 102280 36640
rect 102120 36640 102280 36800
rect 102120 36800 102280 36960
rect 102120 36960 102280 37120
rect 102120 37120 102280 37280
rect 102120 37280 102280 37440
rect 102120 46400 102280 46560
rect 102120 46560 102280 46720
rect 102120 46720 102280 46880
rect 102120 46880 102280 47040
rect 102120 47040 102280 47200
rect 102120 47200 102280 47360
rect 102120 47360 102280 47520
rect 102120 47520 102280 47680
rect 102120 47680 102280 47840
rect 102120 47840 102280 48000
rect 102120 48000 102280 48160
rect 102120 48160 102280 48320
rect 102120 48320 102280 48480
rect 102120 48480 102280 48640
rect 102120 48640 102280 48800
rect 102120 48800 102280 48960
rect 102120 48960 102280 49120
rect 102120 49120 102280 49280
rect 102120 49280 102280 49440
rect 102120 49440 102280 49600
rect 102120 49600 102280 49760
rect 102120 49760 102280 49920
rect 102120 49920 102280 50080
rect 102120 50080 102280 50240
rect 102120 50240 102280 50400
rect 102120 50400 102280 50560
rect 102120 50560 102280 50720
rect 102120 50720 102280 50880
rect 102120 50880 102280 51040
rect 102120 51040 102280 51200
rect 102120 51200 102280 51360
rect 102120 51360 102280 51520
rect 102120 51520 102280 51680
rect 102120 51680 102280 51840
rect 102120 51840 102280 52000
rect 102120 52000 102280 52160
rect 102120 52160 102280 52320
rect 102120 52320 102280 52480
rect 102120 52480 102280 52640
rect 102120 52640 102280 52800
rect 102280 33920 102440 34080
rect 102280 34080 102440 34240
rect 102280 34240 102440 34400
rect 102280 34400 102440 34560
rect 102280 34560 102440 34720
rect 102280 34720 102440 34880
rect 102280 34880 102440 35040
rect 102280 35040 102440 35200
rect 102280 35200 102440 35360
rect 102280 35360 102440 35520
rect 102280 35520 102440 35680
rect 102280 35680 102440 35840
rect 102280 35840 102440 36000
rect 102280 36000 102440 36160
rect 102280 36160 102440 36320
rect 102280 36320 102440 36480
rect 102280 36480 102440 36640
rect 102280 36640 102440 36800
rect 102280 36800 102440 36960
rect 102280 36960 102440 37120
rect 102280 37120 102440 37280
rect 102280 37280 102440 37440
rect 102280 37440 102440 37600
rect 102280 46400 102440 46560
rect 102280 46560 102440 46720
rect 102280 46720 102440 46880
rect 102280 46880 102440 47040
rect 102280 47040 102440 47200
rect 102280 47200 102440 47360
rect 102280 47360 102440 47520
rect 102280 47520 102440 47680
rect 102280 47680 102440 47840
rect 102280 47840 102440 48000
rect 102280 48000 102440 48160
rect 102280 48160 102440 48320
rect 102280 48320 102440 48480
rect 102280 48480 102440 48640
rect 102280 48640 102440 48800
rect 102280 48800 102440 48960
rect 102280 48960 102440 49120
rect 102280 49120 102440 49280
rect 102280 49280 102440 49440
rect 102280 49440 102440 49600
rect 102280 49600 102440 49760
rect 102280 49760 102440 49920
rect 102280 49920 102440 50080
rect 102280 50080 102440 50240
rect 102280 50240 102440 50400
rect 102280 50400 102440 50560
rect 102280 50560 102440 50720
rect 102280 50720 102440 50880
rect 102280 50880 102440 51040
rect 102280 51040 102440 51200
rect 102280 51200 102440 51360
rect 102280 51360 102440 51520
rect 102280 51520 102440 51680
rect 102280 51680 102440 51840
rect 102280 51840 102440 52000
rect 102280 52000 102440 52160
rect 102280 52160 102440 52320
rect 102280 52320 102440 52480
rect 102280 52480 102440 52640
rect 102280 52640 102440 52800
rect 102440 34080 102600 34240
rect 102440 34240 102600 34400
rect 102440 34400 102600 34560
rect 102440 34560 102600 34720
rect 102440 34720 102600 34880
rect 102440 34880 102600 35040
rect 102440 35040 102600 35200
rect 102440 35200 102600 35360
rect 102440 35360 102600 35520
rect 102440 35520 102600 35680
rect 102440 35680 102600 35840
rect 102440 35840 102600 36000
rect 102440 36000 102600 36160
rect 102440 36160 102600 36320
rect 102440 36320 102600 36480
rect 102440 36480 102600 36640
rect 102440 36640 102600 36800
rect 102440 36800 102600 36960
rect 102440 36960 102600 37120
rect 102440 37120 102600 37280
rect 102440 37280 102600 37440
rect 102440 37440 102600 37600
rect 102440 46240 102600 46400
rect 102440 46400 102600 46560
rect 102440 46560 102600 46720
rect 102440 46720 102600 46880
rect 102440 46880 102600 47040
rect 102440 47040 102600 47200
rect 102440 47200 102600 47360
rect 102440 47360 102600 47520
rect 102440 47520 102600 47680
rect 102440 47680 102600 47840
rect 102440 47840 102600 48000
rect 102440 48000 102600 48160
rect 102440 48160 102600 48320
rect 102440 48320 102600 48480
rect 102440 48480 102600 48640
rect 102440 48640 102600 48800
rect 102440 48800 102600 48960
rect 102440 48960 102600 49120
rect 102440 49120 102600 49280
rect 102440 49280 102600 49440
rect 102440 49440 102600 49600
rect 102440 49600 102600 49760
rect 102440 49760 102600 49920
rect 102440 49920 102600 50080
rect 102440 50080 102600 50240
rect 102440 50240 102600 50400
rect 102440 50400 102600 50560
rect 102440 50560 102600 50720
rect 102440 50720 102600 50880
rect 102440 50880 102600 51040
rect 102440 51040 102600 51200
rect 102440 51200 102600 51360
rect 102440 51360 102600 51520
rect 102440 51520 102600 51680
rect 102440 51680 102600 51840
rect 102440 51840 102600 52000
rect 102440 52000 102600 52160
rect 102440 52160 102600 52320
rect 102440 52320 102600 52480
rect 102440 52480 102600 52640
rect 102440 52640 102600 52800
rect 102440 52800 102600 52960
rect 102600 34240 102760 34400
rect 102600 34400 102760 34560
rect 102600 34560 102760 34720
rect 102600 34720 102760 34880
rect 102600 34880 102760 35040
rect 102600 35040 102760 35200
rect 102600 35200 102760 35360
rect 102600 35360 102760 35520
rect 102600 35520 102760 35680
rect 102600 35680 102760 35840
rect 102600 35840 102760 36000
rect 102600 36000 102760 36160
rect 102600 36160 102760 36320
rect 102600 36320 102760 36480
rect 102600 36480 102760 36640
rect 102600 36640 102760 36800
rect 102600 36800 102760 36960
rect 102600 36960 102760 37120
rect 102600 37120 102760 37280
rect 102600 37280 102760 37440
rect 102600 37440 102760 37600
rect 102600 37600 102760 37760
rect 102600 46080 102760 46240
rect 102600 46240 102760 46400
rect 102600 46400 102760 46560
rect 102600 46560 102760 46720
rect 102600 46720 102760 46880
rect 102600 46880 102760 47040
rect 102600 47040 102760 47200
rect 102600 47200 102760 47360
rect 102600 47360 102760 47520
rect 102600 47520 102760 47680
rect 102600 47680 102760 47840
rect 102600 47840 102760 48000
rect 102600 48000 102760 48160
rect 102600 48160 102760 48320
rect 102600 48320 102760 48480
rect 102600 48480 102760 48640
rect 102600 48640 102760 48800
rect 102600 48800 102760 48960
rect 102600 48960 102760 49120
rect 102600 49120 102760 49280
rect 102600 49280 102760 49440
rect 102600 49440 102760 49600
rect 102600 49600 102760 49760
rect 102600 49760 102760 49920
rect 102600 49920 102760 50080
rect 102600 50080 102760 50240
rect 102600 50240 102760 50400
rect 102600 50400 102760 50560
rect 102600 50560 102760 50720
rect 102600 50720 102760 50880
rect 102600 50880 102760 51040
rect 102600 51040 102760 51200
rect 102600 51200 102760 51360
rect 102600 51360 102760 51520
rect 102600 51520 102760 51680
rect 102600 51680 102760 51840
rect 102600 51840 102760 52000
rect 102600 52000 102760 52160
rect 102600 52160 102760 52320
rect 102600 52320 102760 52480
rect 102600 52480 102760 52640
rect 102600 52640 102760 52800
rect 102600 52800 102760 52960
rect 102760 34400 102920 34560
rect 102760 34560 102920 34720
rect 102760 34720 102920 34880
rect 102760 34880 102920 35040
rect 102760 35040 102920 35200
rect 102760 35200 102920 35360
rect 102760 35360 102920 35520
rect 102760 35520 102920 35680
rect 102760 35680 102920 35840
rect 102760 35840 102920 36000
rect 102760 36000 102920 36160
rect 102760 36160 102920 36320
rect 102760 36320 102920 36480
rect 102760 36480 102920 36640
rect 102760 36640 102920 36800
rect 102760 36800 102920 36960
rect 102760 36960 102920 37120
rect 102760 37120 102920 37280
rect 102760 37280 102920 37440
rect 102760 37440 102920 37600
rect 102760 37600 102920 37760
rect 102760 37760 102920 37920
rect 102760 46080 102920 46240
rect 102760 46240 102920 46400
rect 102760 46400 102920 46560
rect 102760 46560 102920 46720
rect 102760 46720 102920 46880
rect 102760 46880 102920 47040
rect 102760 47040 102920 47200
rect 102760 47200 102920 47360
rect 102760 47360 102920 47520
rect 102760 47520 102920 47680
rect 102760 47680 102920 47840
rect 102760 47840 102920 48000
rect 102760 48000 102920 48160
rect 102760 48160 102920 48320
rect 102760 48320 102920 48480
rect 102760 48480 102920 48640
rect 102760 48640 102920 48800
rect 102760 48800 102920 48960
rect 102760 48960 102920 49120
rect 102760 49120 102920 49280
rect 102760 49280 102920 49440
rect 102760 49440 102920 49600
rect 102760 49600 102920 49760
rect 102760 49760 102920 49920
rect 102760 49920 102920 50080
rect 102760 50080 102920 50240
rect 102760 50240 102920 50400
rect 102760 50400 102920 50560
rect 102760 50560 102920 50720
rect 102760 50720 102920 50880
rect 102760 50880 102920 51040
rect 102760 51040 102920 51200
rect 102760 51200 102920 51360
rect 102760 51360 102920 51520
rect 102760 51520 102920 51680
rect 102760 51680 102920 51840
rect 102760 51840 102920 52000
rect 102760 52000 102920 52160
rect 102760 52160 102920 52320
rect 102760 52320 102920 52480
rect 102760 52480 102920 52640
rect 102760 52640 102920 52800
rect 102760 52800 102920 52960
rect 102760 52960 102920 53120
rect 102920 34560 103080 34720
rect 102920 34720 103080 34880
rect 102920 34880 103080 35040
rect 102920 35040 103080 35200
rect 102920 35200 103080 35360
rect 102920 35360 103080 35520
rect 102920 35520 103080 35680
rect 102920 35680 103080 35840
rect 102920 35840 103080 36000
rect 102920 36000 103080 36160
rect 102920 36160 103080 36320
rect 102920 36320 103080 36480
rect 102920 36480 103080 36640
rect 102920 36640 103080 36800
rect 102920 36800 103080 36960
rect 102920 36960 103080 37120
rect 102920 37120 103080 37280
rect 102920 37280 103080 37440
rect 102920 37440 103080 37600
rect 102920 37600 103080 37760
rect 102920 37760 103080 37920
rect 102920 37920 103080 38080
rect 102920 45920 103080 46080
rect 102920 46080 103080 46240
rect 102920 46240 103080 46400
rect 102920 46400 103080 46560
rect 102920 46560 103080 46720
rect 102920 46720 103080 46880
rect 102920 46880 103080 47040
rect 102920 47040 103080 47200
rect 102920 47200 103080 47360
rect 102920 47360 103080 47520
rect 102920 47520 103080 47680
rect 102920 47680 103080 47840
rect 102920 47840 103080 48000
rect 102920 48000 103080 48160
rect 102920 48160 103080 48320
rect 102920 48320 103080 48480
rect 102920 48480 103080 48640
rect 102920 48640 103080 48800
rect 102920 48800 103080 48960
rect 102920 48960 103080 49120
rect 102920 49120 103080 49280
rect 102920 49280 103080 49440
rect 102920 49440 103080 49600
rect 102920 49600 103080 49760
rect 102920 49760 103080 49920
rect 102920 49920 103080 50080
rect 102920 50080 103080 50240
rect 102920 50240 103080 50400
rect 102920 50400 103080 50560
rect 102920 50560 103080 50720
rect 102920 50720 103080 50880
rect 102920 50880 103080 51040
rect 102920 51040 103080 51200
rect 102920 51200 103080 51360
rect 102920 51360 103080 51520
rect 102920 51520 103080 51680
rect 102920 51680 103080 51840
rect 102920 51840 103080 52000
rect 102920 52000 103080 52160
rect 102920 52160 103080 52320
rect 102920 52320 103080 52480
rect 102920 52480 103080 52640
rect 102920 52640 103080 52800
rect 102920 52800 103080 52960
rect 102920 52960 103080 53120
rect 103080 34720 103240 34880
rect 103080 34880 103240 35040
rect 103080 35040 103240 35200
rect 103080 35200 103240 35360
rect 103080 35360 103240 35520
rect 103080 35520 103240 35680
rect 103080 35680 103240 35840
rect 103080 35840 103240 36000
rect 103080 36000 103240 36160
rect 103080 36160 103240 36320
rect 103080 36320 103240 36480
rect 103080 36480 103240 36640
rect 103080 36640 103240 36800
rect 103080 36800 103240 36960
rect 103080 36960 103240 37120
rect 103080 37120 103240 37280
rect 103080 37280 103240 37440
rect 103080 37440 103240 37600
rect 103080 37600 103240 37760
rect 103080 37760 103240 37920
rect 103080 37920 103240 38080
rect 103080 38080 103240 38240
rect 103080 45920 103240 46080
rect 103080 46080 103240 46240
rect 103080 46240 103240 46400
rect 103080 46400 103240 46560
rect 103080 46560 103240 46720
rect 103080 46720 103240 46880
rect 103080 46880 103240 47040
rect 103080 47040 103240 47200
rect 103080 47200 103240 47360
rect 103080 47360 103240 47520
rect 103080 47520 103240 47680
rect 103080 47680 103240 47840
rect 103080 47840 103240 48000
rect 103080 48000 103240 48160
rect 103080 48160 103240 48320
rect 103080 48320 103240 48480
rect 103080 48480 103240 48640
rect 103080 48640 103240 48800
rect 103080 48800 103240 48960
rect 103080 48960 103240 49120
rect 103080 49120 103240 49280
rect 103080 49280 103240 49440
rect 103080 49440 103240 49600
rect 103080 49600 103240 49760
rect 103080 49760 103240 49920
rect 103080 49920 103240 50080
rect 103080 50080 103240 50240
rect 103080 50240 103240 50400
rect 103080 50400 103240 50560
rect 103080 50560 103240 50720
rect 103080 50720 103240 50880
rect 103080 50880 103240 51040
rect 103080 51040 103240 51200
rect 103080 51200 103240 51360
rect 103080 51360 103240 51520
rect 103080 51520 103240 51680
rect 103080 51680 103240 51840
rect 103080 51840 103240 52000
rect 103080 52000 103240 52160
rect 103080 52160 103240 52320
rect 103080 52320 103240 52480
rect 103080 52480 103240 52640
rect 103080 52640 103240 52800
rect 103080 52800 103240 52960
rect 103080 52960 103240 53120
rect 103080 53120 103240 53280
rect 103240 34880 103400 35040
rect 103240 35040 103400 35200
rect 103240 35200 103400 35360
rect 103240 35360 103400 35520
rect 103240 35520 103400 35680
rect 103240 35680 103400 35840
rect 103240 35840 103400 36000
rect 103240 36000 103400 36160
rect 103240 36160 103400 36320
rect 103240 36320 103400 36480
rect 103240 36480 103400 36640
rect 103240 36640 103400 36800
rect 103240 36800 103400 36960
rect 103240 36960 103400 37120
rect 103240 37120 103400 37280
rect 103240 37280 103400 37440
rect 103240 37440 103400 37600
rect 103240 37600 103400 37760
rect 103240 37760 103400 37920
rect 103240 37920 103400 38080
rect 103240 38080 103400 38240
rect 103240 38240 103400 38400
rect 103240 45760 103400 45920
rect 103240 45920 103400 46080
rect 103240 46080 103400 46240
rect 103240 46240 103400 46400
rect 103240 46400 103400 46560
rect 103240 46560 103400 46720
rect 103240 46720 103400 46880
rect 103240 46880 103400 47040
rect 103240 47040 103400 47200
rect 103240 47200 103400 47360
rect 103240 47360 103400 47520
rect 103240 47520 103400 47680
rect 103240 47680 103400 47840
rect 103240 47840 103400 48000
rect 103240 48000 103400 48160
rect 103240 48160 103400 48320
rect 103240 48320 103400 48480
rect 103240 48480 103400 48640
rect 103240 48640 103400 48800
rect 103240 48800 103400 48960
rect 103240 48960 103400 49120
rect 103240 49120 103400 49280
rect 103240 50080 103400 50240
rect 103240 50240 103400 50400
rect 103240 50400 103400 50560
rect 103240 50560 103400 50720
rect 103240 50720 103400 50880
rect 103240 50880 103400 51040
rect 103240 51040 103400 51200
rect 103240 51200 103400 51360
rect 103240 51360 103400 51520
rect 103240 51520 103400 51680
rect 103240 51680 103400 51840
rect 103240 51840 103400 52000
rect 103240 52000 103400 52160
rect 103240 52160 103400 52320
rect 103240 52320 103400 52480
rect 103240 52480 103400 52640
rect 103240 52640 103400 52800
rect 103240 52800 103400 52960
rect 103240 52960 103400 53120
rect 103240 53120 103400 53280
rect 103400 35040 103560 35200
rect 103400 35200 103560 35360
rect 103400 35360 103560 35520
rect 103400 35520 103560 35680
rect 103400 35680 103560 35840
rect 103400 35840 103560 36000
rect 103400 36000 103560 36160
rect 103400 36160 103560 36320
rect 103400 36320 103560 36480
rect 103400 36480 103560 36640
rect 103400 36640 103560 36800
rect 103400 36800 103560 36960
rect 103400 36960 103560 37120
rect 103400 37120 103560 37280
rect 103400 37280 103560 37440
rect 103400 37440 103560 37600
rect 103400 37600 103560 37760
rect 103400 37760 103560 37920
rect 103400 37920 103560 38080
rect 103400 38080 103560 38240
rect 103400 38240 103560 38400
rect 103400 38400 103560 38560
rect 103400 45760 103560 45920
rect 103400 45920 103560 46080
rect 103400 46080 103560 46240
rect 103400 46240 103560 46400
rect 103400 46400 103560 46560
rect 103400 46560 103560 46720
rect 103400 46720 103560 46880
rect 103400 46880 103560 47040
rect 103400 47040 103560 47200
rect 103400 47200 103560 47360
rect 103400 47360 103560 47520
rect 103400 47520 103560 47680
rect 103400 47680 103560 47840
rect 103400 47840 103560 48000
rect 103400 48000 103560 48160
rect 103400 48160 103560 48320
rect 103400 48320 103560 48480
rect 103400 48480 103560 48640
rect 103400 48640 103560 48800
rect 103400 48800 103560 48960
rect 103400 48960 103560 49120
rect 103400 50400 103560 50560
rect 103400 50560 103560 50720
rect 103400 50720 103560 50880
rect 103400 50880 103560 51040
rect 103400 51040 103560 51200
rect 103400 51200 103560 51360
rect 103400 51360 103560 51520
rect 103400 51520 103560 51680
rect 103400 51680 103560 51840
rect 103400 51840 103560 52000
rect 103400 52000 103560 52160
rect 103400 52160 103560 52320
rect 103400 52320 103560 52480
rect 103400 52480 103560 52640
rect 103400 52640 103560 52800
rect 103400 52800 103560 52960
rect 103400 52960 103560 53120
rect 103400 53120 103560 53280
rect 103560 35200 103720 35360
rect 103560 35360 103720 35520
rect 103560 35520 103720 35680
rect 103560 35680 103720 35840
rect 103560 35840 103720 36000
rect 103560 36000 103720 36160
rect 103560 36160 103720 36320
rect 103560 36320 103720 36480
rect 103560 36480 103720 36640
rect 103560 36640 103720 36800
rect 103560 36800 103720 36960
rect 103560 36960 103720 37120
rect 103560 37120 103720 37280
rect 103560 37280 103720 37440
rect 103560 37440 103720 37600
rect 103560 37600 103720 37760
rect 103560 37760 103720 37920
rect 103560 37920 103720 38080
rect 103560 38080 103720 38240
rect 103560 38240 103720 38400
rect 103560 38400 103720 38560
rect 103560 45600 103720 45760
rect 103560 45760 103720 45920
rect 103560 45920 103720 46080
rect 103560 46080 103720 46240
rect 103560 46240 103720 46400
rect 103560 46400 103720 46560
rect 103560 46560 103720 46720
rect 103560 46720 103720 46880
rect 103560 46880 103720 47040
rect 103560 47040 103720 47200
rect 103560 47200 103720 47360
rect 103560 47360 103720 47520
rect 103560 47520 103720 47680
rect 103560 47680 103720 47840
rect 103560 47840 103720 48000
rect 103560 48000 103720 48160
rect 103560 48160 103720 48320
rect 103560 48320 103720 48480
rect 103560 48480 103720 48640
rect 103560 48640 103720 48800
rect 103560 48800 103720 48960
rect 103560 50560 103720 50720
rect 103560 50720 103720 50880
rect 103560 50880 103720 51040
rect 103560 51040 103720 51200
rect 103560 51200 103720 51360
rect 103560 51360 103720 51520
rect 103560 51520 103720 51680
rect 103560 51680 103720 51840
rect 103560 51840 103720 52000
rect 103560 52000 103720 52160
rect 103560 52160 103720 52320
rect 103560 52320 103720 52480
rect 103560 52480 103720 52640
rect 103560 52640 103720 52800
rect 103560 52800 103720 52960
rect 103560 52960 103720 53120
rect 103560 53120 103720 53280
rect 103720 35200 103880 35360
rect 103720 35360 103880 35520
rect 103720 35520 103880 35680
rect 103720 35680 103880 35840
rect 103720 35840 103880 36000
rect 103720 36000 103880 36160
rect 103720 36160 103880 36320
rect 103720 36320 103880 36480
rect 103720 36480 103880 36640
rect 103720 36640 103880 36800
rect 103720 36800 103880 36960
rect 103720 36960 103880 37120
rect 103720 37120 103880 37280
rect 103720 37280 103880 37440
rect 103720 37440 103880 37600
rect 103720 37600 103880 37760
rect 103720 37760 103880 37920
rect 103720 37920 103880 38080
rect 103720 38080 103880 38240
rect 103720 38240 103880 38400
rect 103720 38400 103880 38560
rect 103720 38560 103880 38720
rect 103720 45440 103880 45600
rect 103720 45600 103880 45760
rect 103720 45760 103880 45920
rect 103720 45920 103880 46080
rect 103720 46080 103880 46240
rect 103720 46240 103880 46400
rect 103720 46400 103880 46560
rect 103720 46560 103880 46720
rect 103720 46720 103880 46880
rect 103720 46880 103880 47040
rect 103720 47040 103880 47200
rect 103720 47200 103880 47360
rect 103720 47360 103880 47520
rect 103720 47520 103880 47680
rect 103720 47680 103880 47840
rect 103720 47840 103880 48000
rect 103720 48000 103880 48160
rect 103720 48160 103880 48320
rect 103720 48320 103880 48480
rect 103720 48480 103880 48640
rect 103720 48640 103880 48800
rect 103720 50720 103880 50880
rect 103720 50880 103880 51040
rect 103720 51040 103880 51200
rect 103720 51200 103880 51360
rect 103720 51360 103880 51520
rect 103720 51520 103880 51680
rect 103720 51680 103880 51840
rect 103720 51840 103880 52000
rect 103720 52000 103880 52160
rect 103720 52160 103880 52320
rect 103720 52320 103880 52480
rect 103720 52480 103880 52640
rect 103720 52640 103880 52800
rect 103720 52800 103880 52960
rect 103720 52960 103880 53120
rect 103720 53120 103880 53280
rect 103720 53280 103880 53440
rect 103880 35360 104040 35520
rect 103880 35520 104040 35680
rect 103880 35680 104040 35840
rect 103880 35840 104040 36000
rect 103880 36000 104040 36160
rect 103880 36160 104040 36320
rect 103880 36320 104040 36480
rect 103880 36480 104040 36640
rect 103880 36640 104040 36800
rect 103880 36800 104040 36960
rect 103880 36960 104040 37120
rect 103880 37120 104040 37280
rect 103880 37280 104040 37440
rect 103880 37440 104040 37600
rect 103880 37600 104040 37760
rect 103880 37760 104040 37920
rect 103880 37920 104040 38080
rect 103880 38080 104040 38240
rect 103880 38240 104040 38400
rect 103880 38400 104040 38560
rect 103880 38560 104040 38720
rect 103880 38720 104040 38880
rect 103880 45280 104040 45440
rect 103880 45440 104040 45600
rect 103880 45600 104040 45760
rect 103880 45760 104040 45920
rect 103880 45920 104040 46080
rect 103880 46080 104040 46240
rect 103880 46240 104040 46400
rect 103880 46400 104040 46560
rect 103880 46560 104040 46720
rect 103880 46720 104040 46880
rect 103880 46880 104040 47040
rect 103880 47040 104040 47200
rect 103880 47200 104040 47360
rect 103880 47360 104040 47520
rect 103880 47520 104040 47680
rect 103880 47680 104040 47840
rect 103880 47840 104040 48000
rect 103880 48000 104040 48160
rect 103880 48160 104040 48320
rect 103880 48320 104040 48480
rect 103880 48480 104040 48640
rect 103880 50720 104040 50880
rect 103880 50880 104040 51040
rect 103880 51040 104040 51200
rect 103880 51200 104040 51360
rect 103880 51360 104040 51520
rect 103880 51520 104040 51680
rect 103880 51680 104040 51840
rect 103880 51840 104040 52000
rect 103880 52000 104040 52160
rect 103880 52160 104040 52320
rect 103880 52320 104040 52480
rect 103880 52480 104040 52640
rect 103880 52640 104040 52800
rect 103880 52800 104040 52960
rect 103880 52960 104040 53120
rect 103880 53120 104040 53280
rect 103880 53280 104040 53440
rect 104040 35520 104200 35680
rect 104040 35680 104200 35840
rect 104040 35840 104200 36000
rect 104040 36000 104200 36160
rect 104040 36160 104200 36320
rect 104040 36320 104200 36480
rect 104040 36480 104200 36640
rect 104040 36640 104200 36800
rect 104040 36800 104200 36960
rect 104040 36960 104200 37120
rect 104040 37120 104200 37280
rect 104040 37280 104200 37440
rect 104040 37440 104200 37600
rect 104040 37600 104200 37760
rect 104040 37760 104200 37920
rect 104040 37920 104200 38080
rect 104040 38080 104200 38240
rect 104040 38240 104200 38400
rect 104040 38400 104200 38560
rect 104040 38560 104200 38720
rect 104040 38720 104200 38880
rect 104040 38880 104200 39040
rect 104040 45280 104200 45440
rect 104040 45440 104200 45600
rect 104040 45600 104200 45760
rect 104040 45760 104200 45920
rect 104040 45920 104200 46080
rect 104040 46080 104200 46240
rect 104040 46240 104200 46400
rect 104040 46400 104200 46560
rect 104040 46560 104200 46720
rect 104040 46720 104200 46880
rect 104040 46880 104200 47040
rect 104040 47040 104200 47200
rect 104040 47200 104200 47360
rect 104040 47360 104200 47520
rect 104040 47520 104200 47680
rect 104040 47680 104200 47840
rect 104040 47840 104200 48000
rect 104040 48000 104200 48160
rect 104040 48160 104200 48320
rect 104040 48320 104200 48480
rect 104040 48480 104200 48640
rect 104040 50880 104200 51040
rect 104040 51040 104200 51200
rect 104040 51200 104200 51360
rect 104040 51360 104200 51520
rect 104040 51520 104200 51680
rect 104040 51680 104200 51840
rect 104040 51840 104200 52000
rect 104040 52000 104200 52160
rect 104040 52160 104200 52320
rect 104040 52320 104200 52480
rect 104040 52480 104200 52640
rect 104040 52640 104200 52800
rect 104040 52800 104200 52960
rect 104040 52960 104200 53120
rect 104040 53120 104200 53280
rect 104040 53280 104200 53440
rect 104200 35680 104360 35840
rect 104200 35840 104360 36000
rect 104200 36000 104360 36160
rect 104200 36160 104360 36320
rect 104200 36320 104360 36480
rect 104200 36480 104360 36640
rect 104200 36640 104360 36800
rect 104200 36800 104360 36960
rect 104200 36960 104360 37120
rect 104200 37120 104360 37280
rect 104200 37280 104360 37440
rect 104200 37440 104360 37600
rect 104200 37600 104360 37760
rect 104200 37760 104360 37920
rect 104200 37920 104360 38080
rect 104200 38080 104360 38240
rect 104200 38240 104360 38400
rect 104200 38400 104360 38560
rect 104200 38560 104360 38720
rect 104200 38720 104360 38880
rect 104200 38880 104360 39040
rect 104200 39040 104360 39200
rect 104200 44960 104360 45120
rect 104200 45120 104360 45280
rect 104200 45280 104360 45440
rect 104200 45440 104360 45600
rect 104200 45600 104360 45760
rect 104200 45760 104360 45920
rect 104200 45920 104360 46080
rect 104200 46080 104360 46240
rect 104200 46240 104360 46400
rect 104200 46400 104360 46560
rect 104200 46560 104360 46720
rect 104200 46720 104360 46880
rect 104200 46880 104360 47040
rect 104200 47040 104360 47200
rect 104200 47200 104360 47360
rect 104200 47360 104360 47520
rect 104200 47520 104360 47680
rect 104200 47680 104360 47840
rect 104200 47840 104360 48000
rect 104200 48000 104360 48160
rect 104200 48160 104360 48320
rect 104200 48320 104360 48480
rect 104200 48480 104360 48640
rect 104200 50880 104360 51040
rect 104200 51040 104360 51200
rect 104200 51200 104360 51360
rect 104200 51360 104360 51520
rect 104200 51520 104360 51680
rect 104200 51680 104360 51840
rect 104200 51840 104360 52000
rect 104200 52000 104360 52160
rect 104200 52160 104360 52320
rect 104200 52320 104360 52480
rect 104200 52480 104360 52640
rect 104200 52640 104360 52800
rect 104200 52800 104360 52960
rect 104200 52960 104360 53120
rect 104200 53120 104360 53280
rect 104200 53280 104360 53440
rect 104360 35840 104520 36000
rect 104360 36000 104520 36160
rect 104360 36160 104520 36320
rect 104360 36320 104520 36480
rect 104360 36480 104520 36640
rect 104360 36640 104520 36800
rect 104360 36800 104520 36960
rect 104360 36960 104520 37120
rect 104360 37120 104520 37280
rect 104360 37280 104520 37440
rect 104360 37440 104520 37600
rect 104360 37600 104520 37760
rect 104360 37760 104520 37920
rect 104360 37920 104520 38080
rect 104360 38080 104520 38240
rect 104360 38240 104520 38400
rect 104360 38400 104520 38560
rect 104360 38560 104520 38720
rect 104360 38720 104520 38880
rect 104360 38880 104520 39040
rect 104360 39040 104520 39200
rect 104360 44800 104520 44960
rect 104360 44960 104520 45120
rect 104360 45120 104520 45280
rect 104360 45280 104520 45440
rect 104360 45440 104520 45600
rect 104360 45600 104520 45760
rect 104360 45760 104520 45920
rect 104360 45920 104520 46080
rect 104360 46080 104520 46240
rect 104360 46240 104520 46400
rect 104360 46400 104520 46560
rect 104360 46560 104520 46720
rect 104360 46720 104520 46880
rect 104360 46880 104520 47040
rect 104360 47040 104520 47200
rect 104360 47200 104520 47360
rect 104360 47360 104520 47520
rect 104360 47520 104520 47680
rect 104360 47680 104520 47840
rect 104360 47840 104520 48000
rect 104360 48000 104520 48160
rect 104360 48160 104520 48320
rect 104360 48320 104520 48480
rect 104360 50880 104520 51040
rect 104360 51040 104520 51200
rect 104360 51200 104520 51360
rect 104360 51360 104520 51520
rect 104360 51520 104520 51680
rect 104360 51680 104520 51840
rect 104360 51840 104520 52000
rect 104360 52000 104520 52160
rect 104360 52160 104520 52320
rect 104360 52320 104520 52480
rect 104360 52480 104520 52640
rect 104360 52640 104520 52800
rect 104360 52800 104520 52960
rect 104360 52960 104520 53120
rect 104360 53120 104520 53280
rect 104360 53280 104520 53440
rect 104520 35840 104680 36000
rect 104520 36000 104680 36160
rect 104520 36160 104680 36320
rect 104520 36320 104680 36480
rect 104520 36480 104680 36640
rect 104520 36640 104680 36800
rect 104520 36800 104680 36960
rect 104520 36960 104680 37120
rect 104520 37120 104680 37280
rect 104520 37280 104680 37440
rect 104520 37440 104680 37600
rect 104520 37600 104680 37760
rect 104520 37760 104680 37920
rect 104520 37920 104680 38080
rect 104520 38080 104680 38240
rect 104520 38240 104680 38400
rect 104520 38400 104680 38560
rect 104520 38560 104680 38720
rect 104520 38720 104680 38880
rect 104520 38880 104680 39040
rect 104520 39040 104680 39200
rect 104520 39200 104680 39360
rect 104520 44480 104680 44640
rect 104520 44640 104680 44800
rect 104520 44800 104680 44960
rect 104520 44960 104680 45120
rect 104520 45120 104680 45280
rect 104520 45280 104680 45440
rect 104520 45440 104680 45600
rect 104520 45600 104680 45760
rect 104520 45760 104680 45920
rect 104520 45920 104680 46080
rect 104520 46080 104680 46240
rect 104520 46240 104680 46400
rect 104520 46400 104680 46560
rect 104520 46560 104680 46720
rect 104520 46720 104680 46880
rect 104520 46880 104680 47040
rect 104520 47040 104680 47200
rect 104520 47200 104680 47360
rect 104520 47360 104680 47520
rect 104520 47520 104680 47680
rect 104520 47680 104680 47840
rect 104520 47840 104680 48000
rect 104520 48000 104680 48160
rect 104520 48160 104680 48320
rect 104520 48320 104680 48480
rect 104520 51040 104680 51200
rect 104520 51200 104680 51360
rect 104520 51360 104680 51520
rect 104520 51520 104680 51680
rect 104520 51680 104680 51840
rect 104520 51840 104680 52000
rect 104520 52000 104680 52160
rect 104520 52160 104680 52320
rect 104520 52320 104680 52480
rect 104520 52480 104680 52640
rect 104520 52640 104680 52800
rect 104520 52800 104680 52960
rect 104520 52960 104680 53120
rect 104520 53120 104680 53280
rect 104520 53280 104680 53440
rect 104680 36000 104840 36160
rect 104680 36160 104840 36320
rect 104680 36320 104840 36480
rect 104680 36480 104840 36640
rect 104680 36640 104840 36800
rect 104680 36800 104840 36960
rect 104680 36960 104840 37120
rect 104680 37120 104840 37280
rect 104680 37280 104840 37440
rect 104680 37440 104840 37600
rect 104680 37600 104840 37760
rect 104680 37760 104840 37920
rect 104680 37920 104840 38080
rect 104680 38080 104840 38240
rect 104680 38240 104840 38400
rect 104680 38400 104840 38560
rect 104680 38560 104840 38720
rect 104680 38720 104840 38880
rect 104680 38880 104840 39040
rect 104680 39040 104840 39200
rect 104680 39200 104840 39360
rect 104680 39360 104840 39520
rect 104680 44320 104840 44480
rect 104680 44480 104840 44640
rect 104680 44640 104840 44800
rect 104680 44800 104840 44960
rect 104680 44960 104840 45120
rect 104680 45120 104840 45280
rect 104680 45280 104840 45440
rect 104680 45440 104840 45600
rect 104680 45600 104840 45760
rect 104680 45760 104840 45920
rect 104680 45920 104840 46080
rect 104680 46080 104840 46240
rect 104680 46240 104840 46400
rect 104680 46400 104840 46560
rect 104680 46560 104840 46720
rect 104680 46720 104840 46880
rect 104680 46880 104840 47040
rect 104680 47040 104840 47200
rect 104680 47200 104840 47360
rect 104680 47360 104840 47520
rect 104680 47520 104840 47680
rect 104680 47680 104840 47840
rect 104680 47840 104840 48000
rect 104680 48000 104840 48160
rect 104680 48160 104840 48320
rect 104680 48320 104840 48480
rect 104680 50880 104840 51040
rect 104680 51040 104840 51200
rect 104680 51200 104840 51360
rect 104680 51360 104840 51520
rect 104680 51520 104840 51680
rect 104680 51680 104840 51840
rect 104680 51840 104840 52000
rect 104680 52000 104840 52160
rect 104680 52160 104840 52320
rect 104680 52320 104840 52480
rect 104680 52480 104840 52640
rect 104680 52640 104840 52800
rect 104680 52800 104840 52960
rect 104680 52960 104840 53120
rect 104680 53120 104840 53280
rect 104680 53280 104840 53440
rect 104840 36160 105000 36320
rect 104840 36320 105000 36480
rect 104840 36480 105000 36640
rect 104840 36640 105000 36800
rect 104840 36800 105000 36960
rect 104840 36960 105000 37120
rect 104840 37120 105000 37280
rect 104840 37280 105000 37440
rect 104840 37440 105000 37600
rect 104840 37600 105000 37760
rect 104840 37760 105000 37920
rect 104840 37920 105000 38080
rect 104840 38080 105000 38240
rect 104840 38240 105000 38400
rect 104840 38400 105000 38560
rect 104840 38560 105000 38720
rect 104840 38720 105000 38880
rect 104840 38880 105000 39040
rect 104840 39040 105000 39200
rect 104840 39200 105000 39360
rect 104840 39360 105000 39520
rect 104840 39520 105000 39680
rect 104840 44000 105000 44160
rect 104840 44160 105000 44320
rect 104840 44320 105000 44480
rect 104840 44480 105000 44640
rect 104840 44640 105000 44800
rect 104840 44800 105000 44960
rect 104840 44960 105000 45120
rect 104840 45120 105000 45280
rect 104840 45280 105000 45440
rect 104840 45440 105000 45600
rect 104840 45600 105000 45760
rect 104840 45760 105000 45920
rect 104840 45920 105000 46080
rect 104840 46080 105000 46240
rect 104840 46240 105000 46400
rect 104840 46400 105000 46560
rect 104840 46560 105000 46720
rect 104840 46720 105000 46880
rect 104840 46880 105000 47040
rect 104840 47040 105000 47200
rect 104840 47200 105000 47360
rect 104840 47360 105000 47520
rect 104840 47520 105000 47680
rect 104840 47680 105000 47840
rect 104840 47840 105000 48000
rect 104840 48000 105000 48160
rect 104840 48160 105000 48320
rect 104840 48320 105000 48480
rect 104840 50880 105000 51040
rect 104840 51040 105000 51200
rect 104840 51200 105000 51360
rect 104840 51360 105000 51520
rect 104840 51520 105000 51680
rect 104840 51680 105000 51840
rect 104840 51840 105000 52000
rect 104840 52000 105000 52160
rect 104840 52160 105000 52320
rect 104840 52320 105000 52480
rect 104840 52480 105000 52640
rect 104840 52640 105000 52800
rect 104840 52800 105000 52960
rect 104840 52960 105000 53120
rect 104840 53120 105000 53280
rect 104840 53280 105000 53440
rect 105000 36320 105160 36480
rect 105000 36480 105160 36640
rect 105000 36640 105160 36800
rect 105000 36800 105160 36960
rect 105000 36960 105160 37120
rect 105000 37120 105160 37280
rect 105000 37280 105160 37440
rect 105000 37440 105160 37600
rect 105000 37600 105160 37760
rect 105000 37760 105160 37920
rect 105000 37920 105160 38080
rect 105000 38080 105160 38240
rect 105000 38240 105160 38400
rect 105000 38400 105160 38560
rect 105000 38560 105160 38720
rect 105000 38720 105160 38880
rect 105000 38880 105160 39040
rect 105000 39040 105160 39200
rect 105000 39200 105160 39360
rect 105000 39360 105160 39520
rect 105000 39520 105160 39680
rect 105000 43520 105160 43680
rect 105000 43680 105160 43840
rect 105000 43840 105160 44000
rect 105000 44000 105160 44160
rect 105000 44160 105160 44320
rect 105000 44320 105160 44480
rect 105000 44480 105160 44640
rect 105000 44640 105160 44800
rect 105000 44800 105160 44960
rect 105000 44960 105160 45120
rect 105000 45120 105160 45280
rect 105000 45280 105160 45440
rect 105000 45440 105160 45600
rect 105000 45600 105160 45760
rect 105000 45760 105160 45920
rect 105000 45920 105160 46080
rect 105000 46080 105160 46240
rect 105000 46240 105160 46400
rect 105000 46400 105160 46560
rect 105000 46560 105160 46720
rect 105000 46720 105160 46880
rect 105000 46880 105160 47040
rect 105000 47040 105160 47200
rect 105000 47200 105160 47360
rect 105000 47360 105160 47520
rect 105000 47520 105160 47680
rect 105000 47680 105160 47840
rect 105000 47840 105160 48000
rect 105000 48000 105160 48160
rect 105000 48160 105160 48320
rect 105000 48320 105160 48480
rect 105000 50880 105160 51040
rect 105000 51040 105160 51200
rect 105000 51200 105160 51360
rect 105000 51360 105160 51520
rect 105000 51520 105160 51680
rect 105000 51680 105160 51840
rect 105000 51840 105160 52000
rect 105000 52000 105160 52160
rect 105000 52160 105160 52320
rect 105000 52320 105160 52480
rect 105000 52480 105160 52640
rect 105000 52640 105160 52800
rect 105000 52800 105160 52960
rect 105000 52960 105160 53120
rect 105000 53120 105160 53280
rect 105000 53280 105160 53440
rect 105160 36480 105320 36640
rect 105160 36640 105320 36800
rect 105160 36800 105320 36960
rect 105160 36960 105320 37120
rect 105160 37120 105320 37280
rect 105160 37280 105320 37440
rect 105160 37440 105320 37600
rect 105160 37600 105320 37760
rect 105160 37760 105320 37920
rect 105160 37920 105320 38080
rect 105160 38080 105320 38240
rect 105160 38240 105320 38400
rect 105160 38400 105320 38560
rect 105160 38560 105320 38720
rect 105160 38720 105320 38880
rect 105160 38880 105320 39040
rect 105160 39040 105320 39200
rect 105160 39200 105320 39360
rect 105160 39360 105320 39520
rect 105160 39520 105320 39680
rect 105160 39680 105320 39840
rect 105160 43200 105320 43360
rect 105160 43360 105320 43520
rect 105160 43520 105320 43680
rect 105160 43680 105320 43840
rect 105160 43840 105320 44000
rect 105160 44000 105320 44160
rect 105160 44160 105320 44320
rect 105160 44320 105320 44480
rect 105160 44480 105320 44640
rect 105160 44640 105320 44800
rect 105160 44800 105320 44960
rect 105160 44960 105320 45120
rect 105160 45120 105320 45280
rect 105160 45280 105320 45440
rect 105160 45440 105320 45600
rect 105160 45600 105320 45760
rect 105160 45760 105320 45920
rect 105160 45920 105320 46080
rect 105160 46080 105320 46240
rect 105160 46240 105320 46400
rect 105160 46400 105320 46560
rect 105160 46560 105320 46720
rect 105160 46720 105320 46880
rect 105160 46880 105320 47040
rect 105160 47040 105320 47200
rect 105160 47200 105320 47360
rect 105160 47360 105320 47520
rect 105160 47520 105320 47680
rect 105160 47680 105320 47840
rect 105160 47840 105320 48000
rect 105160 48000 105320 48160
rect 105160 48160 105320 48320
rect 105160 48320 105320 48480
rect 105160 50720 105320 50880
rect 105160 50880 105320 51040
rect 105160 51040 105320 51200
rect 105160 51200 105320 51360
rect 105160 51360 105320 51520
rect 105160 51520 105320 51680
rect 105160 51680 105320 51840
rect 105160 51840 105320 52000
rect 105160 52000 105320 52160
rect 105160 52160 105320 52320
rect 105160 52320 105320 52480
rect 105160 52480 105320 52640
rect 105160 52640 105320 52800
rect 105160 52800 105320 52960
rect 105160 52960 105320 53120
rect 105160 53120 105320 53280
rect 105160 53280 105320 53440
rect 105320 36480 105480 36640
rect 105320 36640 105480 36800
rect 105320 36800 105480 36960
rect 105320 36960 105480 37120
rect 105320 37120 105480 37280
rect 105320 37280 105480 37440
rect 105320 37440 105480 37600
rect 105320 37600 105480 37760
rect 105320 37760 105480 37920
rect 105320 37920 105480 38080
rect 105320 38080 105480 38240
rect 105320 38240 105480 38400
rect 105320 38400 105480 38560
rect 105320 38560 105480 38720
rect 105320 38720 105480 38880
rect 105320 38880 105480 39040
rect 105320 39040 105480 39200
rect 105320 39200 105480 39360
rect 105320 39360 105480 39520
rect 105320 39520 105480 39680
rect 105320 39680 105480 39840
rect 105320 39840 105480 40000
rect 105320 42880 105480 43040
rect 105320 43040 105480 43200
rect 105320 43200 105480 43360
rect 105320 43360 105480 43520
rect 105320 43520 105480 43680
rect 105320 43680 105480 43840
rect 105320 43840 105480 44000
rect 105320 44000 105480 44160
rect 105320 44160 105480 44320
rect 105320 44320 105480 44480
rect 105320 44480 105480 44640
rect 105320 44640 105480 44800
rect 105320 44800 105480 44960
rect 105320 44960 105480 45120
rect 105320 45120 105480 45280
rect 105320 45280 105480 45440
rect 105320 45440 105480 45600
rect 105320 45600 105480 45760
rect 105320 45760 105480 45920
rect 105320 45920 105480 46080
rect 105320 46080 105480 46240
rect 105320 46240 105480 46400
rect 105320 46400 105480 46560
rect 105320 46560 105480 46720
rect 105320 46720 105480 46880
rect 105320 46880 105480 47040
rect 105320 47040 105480 47200
rect 105320 47200 105480 47360
rect 105320 47360 105480 47520
rect 105320 47520 105480 47680
rect 105320 47680 105480 47840
rect 105320 47840 105480 48000
rect 105320 48000 105480 48160
rect 105320 48160 105480 48320
rect 105320 48320 105480 48480
rect 105320 48480 105480 48640
rect 105320 50400 105480 50560
rect 105320 50560 105480 50720
rect 105320 50720 105480 50880
rect 105320 50880 105480 51040
rect 105320 51040 105480 51200
rect 105320 51200 105480 51360
rect 105320 51360 105480 51520
rect 105320 51520 105480 51680
rect 105320 51680 105480 51840
rect 105320 51840 105480 52000
rect 105320 52000 105480 52160
rect 105320 52160 105480 52320
rect 105320 52320 105480 52480
rect 105320 52480 105480 52640
rect 105320 52640 105480 52800
rect 105320 52800 105480 52960
rect 105320 52960 105480 53120
rect 105320 53120 105480 53280
rect 105320 53280 105480 53440
rect 105480 36640 105640 36800
rect 105480 36800 105640 36960
rect 105480 36960 105640 37120
rect 105480 37120 105640 37280
rect 105480 37280 105640 37440
rect 105480 37440 105640 37600
rect 105480 37600 105640 37760
rect 105480 37760 105640 37920
rect 105480 37920 105640 38080
rect 105480 38080 105640 38240
rect 105480 38240 105640 38400
rect 105480 38400 105640 38560
rect 105480 38560 105640 38720
rect 105480 38720 105640 38880
rect 105480 38880 105640 39040
rect 105480 39040 105640 39200
rect 105480 39200 105640 39360
rect 105480 39360 105640 39520
rect 105480 39520 105640 39680
rect 105480 39680 105640 39840
rect 105480 39840 105640 40000
rect 105480 40000 105640 40160
rect 105480 42400 105640 42560
rect 105480 42560 105640 42720
rect 105480 42720 105640 42880
rect 105480 42880 105640 43040
rect 105480 43040 105640 43200
rect 105480 43200 105640 43360
rect 105480 43360 105640 43520
rect 105480 43520 105640 43680
rect 105480 43680 105640 43840
rect 105480 43840 105640 44000
rect 105480 44000 105640 44160
rect 105480 44160 105640 44320
rect 105480 44320 105640 44480
rect 105480 44480 105640 44640
rect 105480 44640 105640 44800
rect 105480 44800 105640 44960
rect 105480 44960 105640 45120
rect 105480 45120 105640 45280
rect 105480 45280 105640 45440
rect 105480 45440 105640 45600
rect 105480 45600 105640 45760
rect 105480 45760 105640 45920
rect 105480 45920 105640 46080
rect 105480 46080 105640 46240
rect 105480 46240 105640 46400
rect 105480 46400 105640 46560
rect 105480 46560 105640 46720
rect 105480 46720 105640 46880
rect 105480 46880 105640 47040
rect 105480 47040 105640 47200
rect 105480 47200 105640 47360
rect 105480 47360 105640 47520
rect 105480 47520 105640 47680
rect 105480 47680 105640 47840
rect 105480 47840 105640 48000
rect 105480 48000 105640 48160
rect 105480 48160 105640 48320
rect 105480 48320 105640 48480
rect 105480 48480 105640 48640
rect 105480 48640 105640 48800
rect 105480 50080 105640 50240
rect 105480 50240 105640 50400
rect 105480 50400 105640 50560
rect 105480 50560 105640 50720
rect 105480 50720 105640 50880
rect 105480 50880 105640 51040
rect 105480 51040 105640 51200
rect 105480 51200 105640 51360
rect 105480 51360 105640 51520
rect 105480 51520 105640 51680
rect 105480 51680 105640 51840
rect 105480 51840 105640 52000
rect 105480 52000 105640 52160
rect 105480 52160 105640 52320
rect 105480 52320 105640 52480
rect 105480 52480 105640 52640
rect 105480 52640 105640 52800
rect 105480 52800 105640 52960
rect 105480 52960 105640 53120
rect 105480 53120 105640 53280
rect 105640 36800 105800 36960
rect 105640 36960 105800 37120
rect 105640 37120 105800 37280
rect 105640 37280 105800 37440
rect 105640 37440 105800 37600
rect 105640 37600 105800 37760
rect 105640 37760 105800 37920
rect 105640 37920 105800 38080
rect 105640 38080 105800 38240
rect 105640 38240 105800 38400
rect 105640 38400 105800 38560
rect 105640 38560 105800 38720
rect 105640 38720 105800 38880
rect 105640 38880 105800 39040
rect 105640 39040 105800 39200
rect 105640 39200 105800 39360
rect 105640 39360 105800 39520
rect 105640 39520 105800 39680
rect 105640 39680 105800 39840
rect 105640 39840 105800 40000
rect 105640 40000 105800 40160
rect 105640 41920 105800 42080
rect 105640 42080 105800 42240
rect 105640 42240 105800 42400
rect 105640 42400 105800 42560
rect 105640 42560 105800 42720
rect 105640 42720 105800 42880
rect 105640 42880 105800 43040
rect 105640 43040 105800 43200
rect 105640 43200 105800 43360
rect 105640 43360 105800 43520
rect 105640 43520 105800 43680
rect 105640 43680 105800 43840
rect 105640 43840 105800 44000
rect 105640 44000 105800 44160
rect 105640 44160 105800 44320
rect 105640 44320 105800 44480
rect 105640 44480 105800 44640
rect 105640 44640 105800 44800
rect 105640 44800 105800 44960
rect 105640 44960 105800 45120
rect 105640 45120 105800 45280
rect 105640 45280 105800 45440
rect 105640 45440 105800 45600
rect 105640 45600 105800 45760
rect 105640 45760 105800 45920
rect 105640 45920 105800 46080
rect 105640 46080 105800 46240
rect 105640 46240 105800 46400
rect 105640 46400 105800 46560
rect 105640 46560 105800 46720
rect 105640 46720 105800 46880
rect 105640 46880 105800 47040
rect 105640 47040 105800 47200
rect 105640 47200 105800 47360
rect 105640 47360 105800 47520
rect 105640 47520 105800 47680
rect 105640 47680 105800 47840
rect 105640 47840 105800 48000
rect 105640 48000 105800 48160
rect 105640 48160 105800 48320
rect 105640 48320 105800 48480
rect 105640 48480 105800 48640
rect 105640 48640 105800 48800
rect 105640 48800 105800 48960
rect 105640 48960 105800 49120
rect 105640 49120 105800 49280
rect 105640 49280 105800 49440
rect 105640 49440 105800 49600
rect 105640 49600 105800 49760
rect 105640 49760 105800 49920
rect 105640 49920 105800 50080
rect 105640 50080 105800 50240
rect 105640 50240 105800 50400
rect 105640 50400 105800 50560
rect 105640 50560 105800 50720
rect 105640 50720 105800 50880
rect 105640 50880 105800 51040
rect 105640 51040 105800 51200
rect 105640 51200 105800 51360
rect 105640 51360 105800 51520
rect 105640 51520 105800 51680
rect 105640 51680 105800 51840
rect 105640 51840 105800 52000
rect 105640 52000 105800 52160
rect 105640 52160 105800 52320
rect 105640 52320 105800 52480
rect 105640 52480 105800 52640
rect 105640 52640 105800 52800
rect 105640 52800 105800 52960
rect 105640 52960 105800 53120
rect 105640 53120 105800 53280
rect 105800 36800 105960 36960
rect 105800 36960 105960 37120
rect 105800 37120 105960 37280
rect 105800 37280 105960 37440
rect 105800 37440 105960 37600
rect 105800 37600 105960 37760
rect 105800 37760 105960 37920
rect 105800 37920 105960 38080
rect 105800 38080 105960 38240
rect 105800 38240 105960 38400
rect 105800 38400 105960 38560
rect 105800 38560 105960 38720
rect 105800 38720 105960 38880
rect 105800 38880 105960 39040
rect 105800 39040 105960 39200
rect 105800 39200 105960 39360
rect 105800 39360 105960 39520
rect 105800 39520 105960 39680
rect 105800 39680 105960 39840
rect 105800 39840 105960 40000
rect 105800 40000 105960 40160
rect 105800 40160 105960 40320
rect 105800 41440 105960 41600
rect 105800 41600 105960 41760
rect 105800 41760 105960 41920
rect 105800 41920 105960 42080
rect 105800 42080 105960 42240
rect 105800 42240 105960 42400
rect 105800 42400 105960 42560
rect 105800 42560 105960 42720
rect 105800 42720 105960 42880
rect 105800 42880 105960 43040
rect 105800 43040 105960 43200
rect 105800 43200 105960 43360
rect 105800 43360 105960 43520
rect 105800 43520 105960 43680
rect 105800 43680 105960 43840
rect 105800 43840 105960 44000
rect 105800 44000 105960 44160
rect 105800 44160 105960 44320
rect 105800 44320 105960 44480
rect 105800 44480 105960 44640
rect 105800 44640 105960 44800
rect 105800 44800 105960 44960
rect 105800 44960 105960 45120
rect 105800 45120 105960 45280
rect 105800 45280 105960 45440
rect 105800 45440 105960 45600
rect 105800 45600 105960 45760
rect 105800 45760 105960 45920
rect 105800 45920 105960 46080
rect 105800 46080 105960 46240
rect 105800 46240 105960 46400
rect 105800 46400 105960 46560
rect 105800 46560 105960 46720
rect 105800 46720 105960 46880
rect 105800 46880 105960 47040
rect 105800 47040 105960 47200
rect 105800 47200 105960 47360
rect 105800 47360 105960 47520
rect 105800 47520 105960 47680
rect 105800 47680 105960 47840
rect 105800 47840 105960 48000
rect 105800 48000 105960 48160
rect 105800 48160 105960 48320
rect 105800 48320 105960 48480
rect 105800 48480 105960 48640
rect 105800 48640 105960 48800
rect 105800 48800 105960 48960
rect 105800 48960 105960 49120
rect 105800 49120 105960 49280
rect 105800 49280 105960 49440
rect 105800 49440 105960 49600
rect 105800 49600 105960 49760
rect 105800 49760 105960 49920
rect 105800 49920 105960 50080
rect 105800 50080 105960 50240
rect 105800 50240 105960 50400
rect 105800 50400 105960 50560
rect 105800 50560 105960 50720
rect 105800 50720 105960 50880
rect 105800 50880 105960 51040
rect 105800 51040 105960 51200
rect 105800 51200 105960 51360
rect 105800 51360 105960 51520
rect 105800 51520 105960 51680
rect 105800 51680 105960 51840
rect 105800 51840 105960 52000
rect 105800 52000 105960 52160
rect 105800 52160 105960 52320
rect 105800 52320 105960 52480
rect 105800 52480 105960 52640
rect 105800 52640 105960 52800
rect 105800 52800 105960 52960
rect 105800 52960 105960 53120
rect 105800 53120 105960 53280
rect 105960 36960 106120 37120
rect 105960 37120 106120 37280
rect 105960 37280 106120 37440
rect 105960 37440 106120 37600
rect 105960 37600 106120 37760
rect 105960 37760 106120 37920
rect 105960 37920 106120 38080
rect 105960 38080 106120 38240
rect 105960 38240 106120 38400
rect 105960 38400 106120 38560
rect 105960 38560 106120 38720
rect 105960 38720 106120 38880
rect 105960 38880 106120 39040
rect 105960 39040 106120 39200
rect 105960 39200 106120 39360
rect 105960 39360 106120 39520
rect 105960 39520 106120 39680
rect 105960 39680 106120 39840
rect 105960 39840 106120 40000
rect 105960 40000 106120 40160
rect 105960 40160 106120 40320
rect 105960 40320 106120 40480
rect 105960 41120 106120 41280
rect 105960 41280 106120 41440
rect 105960 41440 106120 41600
rect 105960 41600 106120 41760
rect 105960 41760 106120 41920
rect 105960 41920 106120 42080
rect 105960 42080 106120 42240
rect 105960 42240 106120 42400
rect 105960 42400 106120 42560
rect 105960 42560 106120 42720
rect 105960 42720 106120 42880
rect 105960 42880 106120 43040
rect 105960 43040 106120 43200
rect 105960 43200 106120 43360
rect 105960 43360 106120 43520
rect 105960 43520 106120 43680
rect 105960 43680 106120 43840
rect 105960 43840 106120 44000
rect 105960 44000 106120 44160
rect 105960 44160 106120 44320
rect 105960 44320 106120 44480
rect 105960 44480 106120 44640
rect 105960 44640 106120 44800
rect 105960 44800 106120 44960
rect 105960 44960 106120 45120
rect 105960 45120 106120 45280
rect 105960 45280 106120 45440
rect 105960 45440 106120 45600
rect 105960 45600 106120 45760
rect 105960 45760 106120 45920
rect 105960 45920 106120 46080
rect 105960 46080 106120 46240
rect 105960 46240 106120 46400
rect 105960 46400 106120 46560
rect 105960 46560 106120 46720
rect 105960 46720 106120 46880
rect 105960 46880 106120 47040
rect 105960 47040 106120 47200
rect 105960 47200 106120 47360
rect 105960 47360 106120 47520
rect 105960 47520 106120 47680
rect 105960 47680 106120 47840
rect 105960 47840 106120 48000
rect 105960 48000 106120 48160
rect 105960 48160 106120 48320
rect 105960 48320 106120 48480
rect 105960 48480 106120 48640
rect 105960 48640 106120 48800
rect 105960 48800 106120 48960
rect 105960 48960 106120 49120
rect 105960 49120 106120 49280
rect 105960 49280 106120 49440
rect 105960 49440 106120 49600
rect 105960 49600 106120 49760
rect 105960 49760 106120 49920
rect 105960 49920 106120 50080
rect 105960 50080 106120 50240
rect 105960 50240 106120 50400
rect 105960 50400 106120 50560
rect 105960 50560 106120 50720
rect 105960 50720 106120 50880
rect 105960 50880 106120 51040
rect 105960 51040 106120 51200
rect 105960 51200 106120 51360
rect 105960 51360 106120 51520
rect 105960 51520 106120 51680
rect 105960 51680 106120 51840
rect 105960 51840 106120 52000
rect 105960 52000 106120 52160
rect 105960 52160 106120 52320
rect 105960 52320 106120 52480
rect 105960 52480 106120 52640
rect 105960 52640 106120 52800
rect 105960 52800 106120 52960
rect 105960 52960 106120 53120
rect 106120 37120 106280 37280
rect 106120 37280 106280 37440
rect 106120 37440 106280 37600
rect 106120 37600 106280 37760
rect 106120 37760 106280 37920
rect 106120 37920 106280 38080
rect 106120 38080 106280 38240
rect 106120 38240 106280 38400
rect 106120 38400 106280 38560
rect 106120 38560 106280 38720
rect 106120 38720 106280 38880
rect 106120 38880 106280 39040
rect 106120 39040 106280 39200
rect 106120 39200 106280 39360
rect 106120 39360 106280 39520
rect 106120 39520 106280 39680
rect 106120 39680 106280 39840
rect 106120 39840 106280 40000
rect 106120 40000 106280 40160
rect 106120 40160 106280 40320
rect 106120 40320 106280 40480
rect 106120 40480 106280 40640
rect 106120 40640 106280 40800
rect 106120 40800 106280 40960
rect 106120 40960 106280 41120
rect 106120 41120 106280 41280
rect 106120 41280 106280 41440
rect 106120 41440 106280 41600
rect 106120 41600 106280 41760
rect 106120 41760 106280 41920
rect 106120 41920 106280 42080
rect 106120 42080 106280 42240
rect 106120 42240 106280 42400
rect 106120 42400 106280 42560
rect 106120 42560 106280 42720
rect 106120 42720 106280 42880
rect 106120 42880 106280 43040
rect 106120 43040 106280 43200
rect 106120 43200 106280 43360
rect 106120 43360 106280 43520
rect 106120 43520 106280 43680
rect 106120 43680 106280 43840
rect 106120 43840 106280 44000
rect 106120 44000 106280 44160
rect 106120 44160 106280 44320
rect 106120 44320 106280 44480
rect 106120 44480 106280 44640
rect 106120 44640 106280 44800
rect 106120 44800 106280 44960
rect 106120 44960 106280 45120
rect 106120 45120 106280 45280
rect 106120 45280 106280 45440
rect 106120 45440 106280 45600
rect 106120 45600 106280 45760
rect 106120 45760 106280 45920
rect 106120 45920 106280 46080
rect 106120 46080 106280 46240
rect 106120 46240 106280 46400
rect 106120 46400 106280 46560
rect 106120 46560 106280 46720
rect 106120 46720 106280 46880
rect 106120 46880 106280 47040
rect 106120 47040 106280 47200
rect 106120 47200 106280 47360
rect 106120 47360 106280 47520
rect 106120 47520 106280 47680
rect 106120 47680 106280 47840
rect 106120 47840 106280 48000
rect 106120 48000 106280 48160
rect 106120 48160 106280 48320
rect 106120 48320 106280 48480
rect 106120 48480 106280 48640
rect 106120 48640 106280 48800
rect 106120 48800 106280 48960
rect 106120 48960 106280 49120
rect 106120 49120 106280 49280
rect 106120 49280 106280 49440
rect 106120 49440 106280 49600
rect 106120 49600 106280 49760
rect 106120 49760 106280 49920
rect 106120 49920 106280 50080
rect 106120 50080 106280 50240
rect 106120 50240 106280 50400
rect 106120 50400 106280 50560
rect 106120 50560 106280 50720
rect 106120 50720 106280 50880
rect 106120 50880 106280 51040
rect 106120 51040 106280 51200
rect 106120 51200 106280 51360
rect 106120 51360 106280 51520
rect 106120 51520 106280 51680
rect 106120 51680 106280 51840
rect 106120 51840 106280 52000
rect 106120 52000 106280 52160
rect 106120 52160 106280 52320
rect 106120 52320 106280 52480
rect 106120 52480 106280 52640
rect 106120 52640 106280 52800
rect 106120 52800 106280 52960
rect 106120 52960 106280 53120
rect 106280 37120 106440 37280
rect 106280 37280 106440 37440
rect 106280 37440 106440 37600
rect 106280 37600 106440 37760
rect 106280 37760 106440 37920
rect 106280 37920 106440 38080
rect 106280 38080 106440 38240
rect 106280 38240 106440 38400
rect 106280 38400 106440 38560
rect 106280 38560 106440 38720
rect 106280 38720 106440 38880
rect 106280 38880 106440 39040
rect 106280 39040 106440 39200
rect 106280 39200 106440 39360
rect 106280 39360 106440 39520
rect 106280 39520 106440 39680
rect 106280 39680 106440 39840
rect 106280 39840 106440 40000
rect 106280 40000 106440 40160
rect 106280 40160 106440 40320
rect 106280 40320 106440 40480
rect 106280 40480 106440 40640
rect 106280 40640 106440 40800
rect 106280 40800 106440 40960
rect 106280 40960 106440 41120
rect 106280 41120 106440 41280
rect 106280 41280 106440 41440
rect 106280 41440 106440 41600
rect 106280 41600 106440 41760
rect 106280 41760 106440 41920
rect 106280 41920 106440 42080
rect 106280 42080 106440 42240
rect 106280 42240 106440 42400
rect 106280 42400 106440 42560
rect 106280 42560 106440 42720
rect 106280 42720 106440 42880
rect 106280 42880 106440 43040
rect 106280 43040 106440 43200
rect 106280 43200 106440 43360
rect 106280 43360 106440 43520
rect 106280 43520 106440 43680
rect 106280 43680 106440 43840
rect 106280 43840 106440 44000
rect 106280 44000 106440 44160
rect 106280 44160 106440 44320
rect 106280 44320 106440 44480
rect 106280 44480 106440 44640
rect 106280 44640 106440 44800
rect 106280 44800 106440 44960
rect 106280 44960 106440 45120
rect 106280 45120 106440 45280
rect 106280 45280 106440 45440
rect 106280 45440 106440 45600
rect 106280 45600 106440 45760
rect 106280 45760 106440 45920
rect 106280 45920 106440 46080
rect 106280 46080 106440 46240
rect 106280 46240 106440 46400
rect 106280 46400 106440 46560
rect 106280 46560 106440 46720
rect 106280 46720 106440 46880
rect 106280 46880 106440 47040
rect 106280 47040 106440 47200
rect 106280 47200 106440 47360
rect 106280 47360 106440 47520
rect 106280 47520 106440 47680
rect 106280 47680 106440 47840
rect 106280 47840 106440 48000
rect 106280 48000 106440 48160
rect 106280 48160 106440 48320
rect 106280 48320 106440 48480
rect 106280 48480 106440 48640
rect 106280 48640 106440 48800
rect 106280 48800 106440 48960
rect 106280 48960 106440 49120
rect 106280 49120 106440 49280
rect 106280 49280 106440 49440
rect 106280 49440 106440 49600
rect 106280 49600 106440 49760
rect 106280 49760 106440 49920
rect 106280 49920 106440 50080
rect 106280 50080 106440 50240
rect 106280 50240 106440 50400
rect 106280 50400 106440 50560
rect 106280 50560 106440 50720
rect 106280 50720 106440 50880
rect 106280 50880 106440 51040
rect 106280 51040 106440 51200
rect 106280 51200 106440 51360
rect 106280 51360 106440 51520
rect 106280 51520 106440 51680
rect 106280 51680 106440 51840
rect 106280 51840 106440 52000
rect 106280 52000 106440 52160
rect 106280 52160 106440 52320
rect 106280 52320 106440 52480
rect 106280 52480 106440 52640
rect 106280 52640 106440 52800
rect 106280 52800 106440 52960
rect 106440 37280 106600 37440
rect 106440 37440 106600 37600
rect 106440 37600 106600 37760
rect 106440 37760 106600 37920
rect 106440 37920 106600 38080
rect 106440 38080 106600 38240
rect 106440 38240 106600 38400
rect 106440 38400 106600 38560
rect 106440 38560 106600 38720
rect 106440 38720 106600 38880
rect 106440 38880 106600 39040
rect 106440 39040 106600 39200
rect 106440 39200 106600 39360
rect 106440 39360 106600 39520
rect 106440 39520 106600 39680
rect 106440 39680 106600 39840
rect 106440 39840 106600 40000
rect 106440 40000 106600 40160
rect 106440 40160 106600 40320
rect 106440 40320 106600 40480
rect 106440 40480 106600 40640
rect 106440 40640 106600 40800
rect 106440 40800 106600 40960
rect 106440 40960 106600 41120
rect 106440 41120 106600 41280
rect 106440 41280 106600 41440
rect 106440 41440 106600 41600
rect 106440 41600 106600 41760
rect 106440 41760 106600 41920
rect 106440 41920 106600 42080
rect 106440 42080 106600 42240
rect 106440 42240 106600 42400
rect 106440 42400 106600 42560
rect 106440 42560 106600 42720
rect 106440 42720 106600 42880
rect 106440 42880 106600 43040
rect 106440 43040 106600 43200
rect 106440 43200 106600 43360
rect 106440 43360 106600 43520
rect 106440 43520 106600 43680
rect 106440 43680 106600 43840
rect 106440 43840 106600 44000
rect 106440 44000 106600 44160
rect 106440 44160 106600 44320
rect 106440 44320 106600 44480
rect 106440 44480 106600 44640
rect 106440 44640 106600 44800
rect 106440 44800 106600 44960
rect 106440 44960 106600 45120
rect 106440 45120 106600 45280
rect 106440 45280 106600 45440
rect 106440 45440 106600 45600
rect 106440 45600 106600 45760
rect 106440 45760 106600 45920
rect 106440 45920 106600 46080
rect 106440 46080 106600 46240
rect 106440 46240 106600 46400
rect 106440 46400 106600 46560
rect 106440 46560 106600 46720
rect 106440 46720 106600 46880
rect 106440 46880 106600 47040
rect 106440 47040 106600 47200
rect 106440 47200 106600 47360
rect 106440 47360 106600 47520
rect 106440 47520 106600 47680
rect 106440 47680 106600 47840
rect 106440 47840 106600 48000
rect 106440 48000 106600 48160
rect 106440 48160 106600 48320
rect 106440 48320 106600 48480
rect 106440 48480 106600 48640
rect 106440 48640 106600 48800
rect 106440 48800 106600 48960
rect 106440 48960 106600 49120
rect 106440 49120 106600 49280
rect 106440 49280 106600 49440
rect 106440 49440 106600 49600
rect 106440 49600 106600 49760
rect 106440 49760 106600 49920
rect 106440 49920 106600 50080
rect 106440 50080 106600 50240
rect 106440 50240 106600 50400
rect 106440 50400 106600 50560
rect 106440 50560 106600 50720
rect 106440 50720 106600 50880
rect 106440 50880 106600 51040
rect 106440 51040 106600 51200
rect 106440 51200 106600 51360
rect 106440 51360 106600 51520
rect 106440 51520 106600 51680
rect 106440 51680 106600 51840
rect 106440 51840 106600 52000
rect 106440 52000 106600 52160
rect 106440 52160 106600 52320
rect 106440 52320 106600 52480
rect 106440 52480 106600 52640
rect 106440 52640 106600 52800
rect 106440 52800 106600 52960
rect 106600 37280 106760 37440
rect 106600 37440 106760 37600
rect 106600 37600 106760 37760
rect 106600 37760 106760 37920
rect 106600 37920 106760 38080
rect 106600 38080 106760 38240
rect 106600 38240 106760 38400
rect 106600 38400 106760 38560
rect 106600 38560 106760 38720
rect 106600 38720 106760 38880
rect 106600 38880 106760 39040
rect 106600 39040 106760 39200
rect 106600 39200 106760 39360
rect 106600 39360 106760 39520
rect 106600 39520 106760 39680
rect 106600 39680 106760 39840
rect 106600 39840 106760 40000
rect 106600 40000 106760 40160
rect 106600 40160 106760 40320
rect 106600 40320 106760 40480
rect 106600 40480 106760 40640
rect 106600 40640 106760 40800
rect 106600 40800 106760 40960
rect 106600 40960 106760 41120
rect 106600 41120 106760 41280
rect 106600 41280 106760 41440
rect 106600 41440 106760 41600
rect 106600 41600 106760 41760
rect 106600 41760 106760 41920
rect 106600 41920 106760 42080
rect 106600 42080 106760 42240
rect 106600 42240 106760 42400
rect 106600 42400 106760 42560
rect 106600 42560 106760 42720
rect 106600 42720 106760 42880
rect 106600 42880 106760 43040
rect 106600 43040 106760 43200
rect 106600 43200 106760 43360
rect 106600 43360 106760 43520
rect 106600 43520 106760 43680
rect 106600 43680 106760 43840
rect 106600 43840 106760 44000
rect 106600 44000 106760 44160
rect 106600 44160 106760 44320
rect 106600 44320 106760 44480
rect 106600 44480 106760 44640
rect 106600 44640 106760 44800
rect 106600 44800 106760 44960
rect 106600 44960 106760 45120
rect 106600 45120 106760 45280
rect 106600 45280 106760 45440
rect 106600 45440 106760 45600
rect 106600 45600 106760 45760
rect 106600 45760 106760 45920
rect 106600 45920 106760 46080
rect 106600 46080 106760 46240
rect 106600 46240 106760 46400
rect 106600 46400 106760 46560
rect 106600 46560 106760 46720
rect 106600 46720 106760 46880
rect 106600 46880 106760 47040
rect 106600 47040 106760 47200
rect 106600 47200 106760 47360
rect 106600 47360 106760 47520
rect 106600 47520 106760 47680
rect 106600 47680 106760 47840
rect 106600 47840 106760 48000
rect 106600 48000 106760 48160
rect 106600 48160 106760 48320
rect 106600 48320 106760 48480
rect 106600 48480 106760 48640
rect 106600 48640 106760 48800
rect 106600 48800 106760 48960
rect 106600 48960 106760 49120
rect 106600 49120 106760 49280
rect 106600 49280 106760 49440
rect 106600 49440 106760 49600
rect 106600 49600 106760 49760
rect 106600 49760 106760 49920
rect 106600 49920 106760 50080
rect 106600 50080 106760 50240
rect 106600 50240 106760 50400
rect 106600 50400 106760 50560
rect 106600 50560 106760 50720
rect 106600 50720 106760 50880
rect 106600 50880 106760 51040
rect 106600 51040 106760 51200
rect 106600 51200 106760 51360
rect 106600 51360 106760 51520
rect 106600 51520 106760 51680
rect 106600 51680 106760 51840
rect 106600 51840 106760 52000
rect 106600 52000 106760 52160
rect 106600 52160 106760 52320
rect 106600 52320 106760 52480
rect 106600 52480 106760 52640
rect 106600 52640 106760 52800
rect 106760 37440 106920 37600
rect 106760 37600 106920 37760
rect 106760 37760 106920 37920
rect 106760 37920 106920 38080
rect 106760 38080 106920 38240
rect 106760 38240 106920 38400
rect 106760 38400 106920 38560
rect 106760 38560 106920 38720
rect 106760 38720 106920 38880
rect 106760 38880 106920 39040
rect 106760 39040 106920 39200
rect 106760 39200 106920 39360
rect 106760 39360 106920 39520
rect 106760 39520 106920 39680
rect 106760 39680 106920 39840
rect 106760 39840 106920 40000
rect 106760 40000 106920 40160
rect 106760 40160 106920 40320
rect 106760 40320 106920 40480
rect 106760 40480 106920 40640
rect 106760 40640 106920 40800
rect 106760 40800 106920 40960
rect 106760 40960 106920 41120
rect 106760 41120 106920 41280
rect 106760 41280 106920 41440
rect 106760 41440 106920 41600
rect 106760 41600 106920 41760
rect 106760 41760 106920 41920
rect 106760 41920 106920 42080
rect 106760 42080 106920 42240
rect 106760 42240 106920 42400
rect 106760 42400 106920 42560
rect 106760 42560 106920 42720
rect 106760 42720 106920 42880
rect 106760 42880 106920 43040
rect 106760 43040 106920 43200
rect 106760 43200 106920 43360
rect 106760 43360 106920 43520
rect 106760 43520 106920 43680
rect 106760 43680 106920 43840
rect 106760 43840 106920 44000
rect 106760 44000 106920 44160
rect 106760 44160 106920 44320
rect 106760 44320 106920 44480
rect 106760 44480 106920 44640
rect 106760 44640 106920 44800
rect 106760 44800 106920 44960
rect 106760 44960 106920 45120
rect 106760 45120 106920 45280
rect 106760 45280 106920 45440
rect 106760 45440 106920 45600
rect 106760 45600 106920 45760
rect 106760 45760 106920 45920
rect 106760 45920 106920 46080
rect 106760 46080 106920 46240
rect 106760 46240 106920 46400
rect 106760 46400 106920 46560
rect 106760 46560 106920 46720
rect 106760 46720 106920 46880
rect 106760 46880 106920 47040
rect 106760 47040 106920 47200
rect 106760 47200 106920 47360
rect 106760 47360 106920 47520
rect 106760 47520 106920 47680
rect 106760 47680 106920 47840
rect 106760 47840 106920 48000
rect 106760 48000 106920 48160
rect 106760 48160 106920 48320
rect 106760 48320 106920 48480
rect 106760 48480 106920 48640
rect 106760 48640 106920 48800
rect 106760 48800 106920 48960
rect 106760 48960 106920 49120
rect 106760 49120 106920 49280
rect 106760 49280 106920 49440
rect 106760 49440 106920 49600
rect 106760 49600 106920 49760
rect 106760 49760 106920 49920
rect 106760 49920 106920 50080
rect 106760 50080 106920 50240
rect 106760 50240 106920 50400
rect 106760 50400 106920 50560
rect 106760 50560 106920 50720
rect 106760 50720 106920 50880
rect 106760 50880 106920 51040
rect 106760 51040 106920 51200
rect 106760 51200 106920 51360
rect 106760 51360 106920 51520
rect 106760 51520 106920 51680
rect 106760 51680 106920 51840
rect 106760 51840 106920 52000
rect 106760 52000 106920 52160
rect 106760 52160 106920 52320
rect 106760 52320 106920 52480
rect 106760 52480 106920 52640
rect 106760 52640 106920 52800
rect 106920 37440 107080 37600
rect 106920 37600 107080 37760
rect 106920 37760 107080 37920
rect 106920 37920 107080 38080
rect 106920 38080 107080 38240
rect 106920 38240 107080 38400
rect 106920 38400 107080 38560
rect 106920 38560 107080 38720
rect 106920 38720 107080 38880
rect 106920 38880 107080 39040
rect 106920 39040 107080 39200
rect 106920 39200 107080 39360
rect 106920 39360 107080 39520
rect 106920 39520 107080 39680
rect 106920 39680 107080 39840
rect 106920 39840 107080 40000
rect 106920 40000 107080 40160
rect 106920 40160 107080 40320
rect 106920 40320 107080 40480
rect 106920 40480 107080 40640
rect 106920 40640 107080 40800
rect 106920 40800 107080 40960
rect 106920 40960 107080 41120
rect 106920 41120 107080 41280
rect 106920 41280 107080 41440
rect 106920 41440 107080 41600
rect 106920 41600 107080 41760
rect 106920 41760 107080 41920
rect 106920 41920 107080 42080
rect 106920 42080 107080 42240
rect 106920 42240 107080 42400
rect 106920 42400 107080 42560
rect 106920 42560 107080 42720
rect 106920 42720 107080 42880
rect 106920 42880 107080 43040
rect 106920 43040 107080 43200
rect 106920 43200 107080 43360
rect 106920 43360 107080 43520
rect 106920 43520 107080 43680
rect 106920 43680 107080 43840
rect 106920 43840 107080 44000
rect 106920 44000 107080 44160
rect 106920 44160 107080 44320
rect 106920 44320 107080 44480
rect 106920 44480 107080 44640
rect 106920 44640 107080 44800
rect 106920 44800 107080 44960
rect 106920 44960 107080 45120
rect 106920 45120 107080 45280
rect 106920 45280 107080 45440
rect 106920 45440 107080 45600
rect 106920 45600 107080 45760
rect 106920 45760 107080 45920
rect 106920 45920 107080 46080
rect 106920 46080 107080 46240
rect 106920 46240 107080 46400
rect 106920 46400 107080 46560
rect 106920 46560 107080 46720
rect 106920 46720 107080 46880
rect 106920 46880 107080 47040
rect 106920 47040 107080 47200
rect 106920 47200 107080 47360
rect 106920 47360 107080 47520
rect 106920 47520 107080 47680
rect 106920 47680 107080 47840
rect 106920 47840 107080 48000
rect 106920 48000 107080 48160
rect 106920 48160 107080 48320
rect 106920 48320 107080 48480
rect 106920 48480 107080 48640
rect 106920 48640 107080 48800
rect 106920 48800 107080 48960
rect 106920 48960 107080 49120
rect 106920 49120 107080 49280
rect 106920 49280 107080 49440
rect 106920 49440 107080 49600
rect 106920 49600 107080 49760
rect 106920 49760 107080 49920
rect 106920 49920 107080 50080
rect 106920 50080 107080 50240
rect 106920 50240 107080 50400
rect 106920 50400 107080 50560
rect 106920 50560 107080 50720
rect 106920 50720 107080 50880
rect 106920 50880 107080 51040
rect 106920 51040 107080 51200
rect 106920 51200 107080 51360
rect 106920 51360 107080 51520
rect 106920 51520 107080 51680
rect 106920 51680 107080 51840
rect 106920 51840 107080 52000
rect 106920 52000 107080 52160
rect 106920 52160 107080 52320
rect 106920 52320 107080 52480
rect 106920 52480 107080 52640
rect 107080 30080 107240 30240
rect 107080 30240 107240 30400
rect 107080 30400 107240 30560
rect 107080 30560 107240 30720
rect 107080 30720 107240 30880
rect 107080 30880 107240 31040
rect 107080 31040 107240 31200
rect 107080 31200 107240 31360
rect 107080 37600 107240 37760
rect 107080 37760 107240 37920
rect 107080 37920 107240 38080
rect 107080 38080 107240 38240
rect 107080 38240 107240 38400
rect 107080 38400 107240 38560
rect 107080 38560 107240 38720
rect 107080 38720 107240 38880
rect 107080 38880 107240 39040
rect 107080 39040 107240 39200
rect 107080 39200 107240 39360
rect 107080 39360 107240 39520
rect 107080 39520 107240 39680
rect 107080 39680 107240 39840
rect 107080 39840 107240 40000
rect 107080 40000 107240 40160
rect 107080 40160 107240 40320
rect 107080 40320 107240 40480
rect 107080 40480 107240 40640
rect 107080 40640 107240 40800
rect 107080 40800 107240 40960
rect 107080 40960 107240 41120
rect 107080 41120 107240 41280
rect 107080 41280 107240 41440
rect 107080 41440 107240 41600
rect 107080 41600 107240 41760
rect 107080 41760 107240 41920
rect 107080 41920 107240 42080
rect 107080 42080 107240 42240
rect 107080 42240 107240 42400
rect 107080 42400 107240 42560
rect 107080 42560 107240 42720
rect 107080 42720 107240 42880
rect 107080 42880 107240 43040
rect 107080 43040 107240 43200
rect 107080 43200 107240 43360
rect 107080 43360 107240 43520
rect 107080 43520 107240 43680
rect 107080 43680 107240 43840
rect 107080 43840 107240 44000
rect 107080 44000 107240 44160
rect 107080 44160 107240 44320
rect 107080 44320 107240 44480
rect 107080 44480 107240 44640
rect 107080 44640 107240 44800
rect 107080 44800 107240 44960
rect 107080 44960 107240 45120
rect 107080 45120 107240 45280
rect 107080 45280 107240 45440
rect 107080 45440 107240 45600
rect 107080 45600 107240 45760
rect 107080 45760 107240 45920
rect 107080 45920 107240 46080
rect 107080 46080 107240 46240
rect 107080 46240 107240 46400
rect 107080 46400 107240 46560
rect 107080 46560 107240 46720
rect 107080 46720 107240 46880
rect 107080 46880 107240 47040
rect 107080 47040 107240 47200
rect 107080 47200 107240 47360
rect 107080 47360 107240 47520
rect 107080 47520 107240 47680
rect 107080 47680 107240 47840
rect 107080 47840 107240 48000
rect 107080 48000 107240 48160
rect 107080 48160 107240 48320
rect 107080 48320 107240 48480
rect 107080 48480 107240 48640
rect 107080 48640 107240 48800
rect 107080 48800 107240 48960
rect 107080 48960 107240 49120
rect 107080 49120 107240 49280
rect 107080 49280 107240 49440
rect 107080 49440 107240 49600
rect 107080 49600 107240 49760
rect 107080 49760 107240 49920
rect 107080 49920 107240 50080
rect 107080 50080 107240 50240
rect 107080 50240 107240 50400
rect 107080 50400 107240 50560
rect 107080 50560 107240 50720
rect 107080 50720 107240 50880
rect 107080 50880 107240 51040
rect 107080 51040 107240 51200
rect 107080 51200 107240 51360
rect 107080 51360 107240 51520
rect 107080 51520 107240 51680
rect 107080 51680 107240 51840
rect 107080 51840 107240 52000
rect 107080 52000 107240 52160
rect 107080 52160 107240 52320
rect 107080 52320 107240 52480
rect 107240 29280 107400 29440
rect 107240 29440 107400 29600
rect 107240 29600 107400 29760
rect 107240 29760 107400 29920
rect 107240 29920 107400 30080
rect 107240 30080 107400 30240
rect 107240 30240 107400 30400
rect 107240 30400 107400 30560
rect 107240 30560 107400 30720
rect 107240 30720 107400 30880
rect 107240 30880 107400 31040
rect 107240 31040 107400 31200
rect 107240 31200 107400 31360
rect 107240 31360 107400 31520
rect 107240 31520 107400 31680
rect 107240 31680 107400 31840
rect 107240 31840 107400 32000
rect 107240 37280 107400 37440
rect 107240 37440 107400 37600
rect 107240 37600 107400 37760
rect 107240 37760 107400 37920
rect 107240 37920 107400 38080
rect 107240 38080 107400 38240
rect 107240 38240 107400 38400
rect 107240 38400 107400 38560
rect 107240 38560 107400 38720
rect 107240 38720 107400 38880
rect 107240 38880 107400 39040
rect 107240 39040 107400 39200
rect 107240 39200 107400 39360
rect 107240 39360 107400 39520
rect 107240 39520 107400 39680
rect 107240 39680 107400 39840
rect 107240 39840 107400 40000
rect 107240 40000 107400 40160
rect 107240 40160 107400 40320
rect 107240 40320 107400 40480
rect 107240 40480 107400 40640
rect 107240 40640 107400 40800
rect 107240 40800 107400 40960
rect 107240 40960 107400 41120
rect 107240 41120 107400 41280
rect 107240 41280 107400 41440
rect 107240 41440 107400 41600
rect 107240 41600 107400 41760
rect 107240 41760 107400 41920
rect 107240 41920 107400 42080
rect 107240 42080 107400 42240
rect 107240 42240 107400 42400
rect 107240 42400 107400 42560
rect 107240 42560 107400 42720
rect 107240 42720 107400 42880
rect 107240 42880 107400 43040
rect 107240 43040 107400 43200
rect 107240 43200 107400 43360
rect 107240 43360 107400 43520
rect 107240 43520 107400 43680
rect 107240 43680 107400 43840
rect 107240 43840 107400 44000
rect 107240 44000 107400 44160
rect 107240 44160 107400 44320
rect 107240 44320 107400 44480
rect 107240 44480 107400 44640
rect 107240 44640 107400 44800
rect 107240 44800 107400 44960
rect 107240 44960 107400 45120
rect 107240 45120 107400 45280
rect 107240 45280 107400 45440
rect 107240 45440 107400 45600
rect 107240 45600 107400 45760
rect 107240 45760 107400 45920
rect 107240 45920 107400 46080
rect 107240 46080 107400 46240
rect 107240 46240 107400 46400
rect 107240 46400 107400 46560
rect 107240 46560 107400 46720
rect 107240 46720 107400 46880
rect 107240 46880 107400 47040
rect 107240 47040 107400 47200
rect 107240 47200 107400 47360
rect 107240 47360 107400 47520
rect 107240 47520 107400 47680
rect 107240 47680 107400 47840
rect 107240 47840 107400 48000
rect 107240 48000 107400 48160
rect 107240 48160 107400 48320
rect 107240 48320 107400 48480
rect 107240 48480 107400 48640
rect 107240 48640 107400 48800
rect 107240 48800 107400 48960
rect 107240 48960 107400 49120
rect 107240 49120 107400 49280
rect 107240 49280 107400 49440
rect 107240 49440 107400 49600
rect 107240 49600 107400 49760
rect 107240 49760 107400 49920
rect 107240 49920 107400 50080
rect 107240 50080 107400 50240
rect 107240 50240 107400 50400
rect 107240 50400 107400 50560
rect 107240 50560 107400 50720
rect 107240 50720 107400 50880
rect 107240 50880 107400 51040
rect 107240 51040 107400 51200
rect 107240 51200 107400 51360
rect 107240 51360 107400 51520
rect 107240 51520 107400 51680
rect 107240 51680 107400 51840
rect 107240 51840 107400 52000
rect 107240 52000 107400 52160
rect 107240 52160 107400 52320
rect 107400 28960 107560 29120
rect 107400 29120 107560 29280
rect 107400 29280 107560 29440
rect 107400 29440 107560 29600
rect 107400 29600 107560 29760
rect 107400 29760 107560 29920
rect 107400 29920 107560 30080
rect 107400 30080 107560 30240
rect 107400 30240 107560 30400
rect 107400 30400 107560 30560
rect 107400 30560 107560 30720
rect 107400 30720 107560 30880
rect 107400 30880 107560 31040
rect 107400 31040 107560 31200
rect 107400 31200 107560 31360
rect 107400 31360 107560 31520
rect 107400 31520 107560 31680
rect 107400 31680 107560 31840
rect 107400 31840 107560 32000
rect 107400 32000 107560 32160
rect 107400 32160 107560 32320
rect 107400 32320 107560 32480
rect 107400 36800 107560 36960
rect 107400 36960 107560 37120
rect 107400 37120 107560 37280
rect 107400 37280 107560 37440
rect 107400 37440 107560 37600
rect 107400 37600 107560 37760
rect 107400 37760 107560 37920
rect 107400 37920 107560 38080
rect 107400 38080 107560 38240
rect 107400 38240 107560 38400
rect 107400 38400 107560 38560
rect 107400 38560 107560 38720
rect 107400 38720 107560 38880
rect 107400 38880 107560 39040
rect 107400 39040 107560 39200
rect 107400 39200 107560 39360
rect 107400 39360 107560 39520
rect 107400 39520 107560 39680
rect 107400 39680 107560 39840
rect 107400 39840 107560 40000
rect 107400 40000 107560 40160
rect 107400 40160 107560 40320
rect 107400 40320 107560 40480
rect 107400 40480 107560 40640
rect 107400 40640 107560 40800
rect 107400 40800 107560 40960
rect 107400 40960 107560 41120
rect 107400 41120 107560 41280
rect 107400 41280 107560 41440
rect 107400 41440 107560 41600
rect 107400 41600 107560 41760
rect 107400 41760 107560 41920
rect 107400 41920 107560 42080
rect 107400 42080 107560 42240
rect 107400 42240 107560 42400
rect 107400 42400 107560 42560
rect 107400 42560 107560 42720
rect 107400 42720 107560 42880
rect 107400 42880 107560 43040
rect 107400 43040 107560 43200
rect 107400 43200 107560 43360
rect 107400 43360 107560 43520
rect 107400 43520 107560 43680
rect 107400 43680 107560 43840
rect 107400 43840 107560 44000
rect 107400 44000 107560 44160
rect 107400 44160 107560 44320
rect 107400 44320 107560 44480
rect 107400 44480 107560 44640
rect 107400 44640 107560 44800
rect 107400 44800 107560 44960
rect 107400 44960 107560 45120
rect 107400 45120 107560 45280
rect 107400 45280 107560 45440
rect 107400 46720 107560 46880
rect 107400 46880 107560 47040
rect 107400 47040 107560 47200
rect 107400 47200 107560 47360
rect 107400 47360 107560 47520
rect 107400 47520 107560 47680
rect 107400 47680 107560 47840
rect 107400 47840 107560 48000
rect 107400 48000 107560 48160
rect 107400 48160 107560 48320
rect 107400 48320 107560 48480
rect 107400 48480 107560 48640
rect 107400 48640 107560 48800
rect 107400 48800 107560 48960
rect 107400 48960 107560 49120
rect 107400 49120 107560 49280
rect 107400 49280 107560 49440
rect 107400 49440 107560 49600
rect 107400 49600 107560 49760
rect 107400 49760 107560 49920
rect 107400 49920 107560 50080
rect 107400 50080 107560 50240
rect 107400 50240 107560 50400
rect 107400 50400 107560 50560
rect 107400 50560 107560 50720
rect 107400 50720 107560 50880
rect 107400 50880 107560 51040
rect 107400 51040 107560 51200
rect 107400 51200 107560 51360
rect 107400 51360 107560 51520
rect 107400 51520 107560 51680
rect 107400 51680 107560 51840
rect 107400 51840 107560 52000
rect 107400 52000 107560 52160
rect 107560 28480 107720 28640
rect 107560 28640 107720 28800
rect 107560 28800 107720 28960
rect 107560 28960 107720 29120
rect 107560 29120 107720 29280
rect 107560 29280 107720 29440
rect 107560 29440 107720 29600
rect 107560 29600 107720 29760
rect 107560 29760 107720 29920
rect 107560 29920 107720 30080
rect 107560 30080 107720 30240
rect 107560 30240 107720 30400
rect 107560 30400 107720 30560
rect 107560 30560 107720 30720
rect 107560 30720 107720 30880
rect 107560 30880 107720 31040
rect 107560 31040 107720 31200
rect 107560 31200 107720 31360
rect 107560 31360 107720 31520
rect 107560 31520 107720 31680
rect 107560 31680 107720 31840
rect 107560 31840 107720 32000
rect 107560 32000 107720 32160
rect 107560 32160 107720 32320
rect 107560 32320 107720 32480
rect 107560 32480 107720 32640
rect 107560 32640 107720 32800
rect 107560 36160 107720 36320
rect 107560 36320 107720 36480
rect 107560 36480 107720 36640
rect 107560 36640 107720 36800
rect 107560 36800 107720 36960
rect 107560 36960 107720 37120
rect 107560 37120 107720 37280
rect 107560 37280 107720 37440
rect 107560 37440 107720 37600
rect 107560 37600 107720 37760
rect 107560 37760 107720 37920
rect 107560 37920 107720 38080
rect 107560 38080 107720 38240
rect 107560 38240 107720 38400
rect 107560 38400 107720 38560
rect 107560 38560 107720 38720
rect 107560 38720 107720 38880
rect 107560 38880 107720 39040
rect 107560 39040 107720 39200
rect 107560 39200 107720 39360
rect 107560 39360 107720 39520
rect 107560 39520 107720 39680
rect 107560 39680 107720 39840
rect 107560 39840 107720 40000
rect 107560 40000 107720 40160
rect 107560 40160 107720 40320
rect 107560 40320 107720 40480
rect 107560 40480 107720 40640
rect 107560 40640 107720 40800
rect 107560 40800 107720 40960
rect 107560 40960 107720 41120
rect 107560 41120 107720 41280
rect 107560 41280 107720 41440
rect 107560 41440 107720 41600
rect 107560 41600 107720 41760
rect 107560 41760 107720 41920
rect 107560 41920 107720 42080
rect 107560 42080 107720 42240
rect 107560 42240 107720 42400
rect 107560 42400 107720 42560
rect 107560 42560 107720 42720
rect 107560 42720 107720 42880
rect 107560 42880 107720 43040
rect 107560 43040 107720 43200
rect 107560 43200 107720 43360
rect 107560 43360 107720 43520
rect 107560 43520 107720 43680
rect 107560 43680 107720 43840
rect 107560 43840 107720 44000
rect 107560 44000 107720 44160
rect 107560 44160 107720 44320
rect 107560 44320 107720 44480
rect 107560 44480 107720 44640
rect 107560 47200 107720 47360
rect 107560 47360 107720 47520
rect 107560 47520 107720 47680
rect 107560 47680 107720 47840
rect 107560 47840 107720 48000
rect 107560 48000 107720 48160
rect 107560 48160 107720 48320
rect 107560 48320 107720 48480
rect 107560 48480 107720 48640
rect 107560 48640 107720 48800
rect 107560 48800 107720 48960
rect 107560 48960 107720 49120
rect 107560 49120 107720 49280
rect 107560 49280 107720 49440
rect 107560 49440 107720 49600
rect 107560 49600 107720 49760
rect 107560 49760 107720 49920
rect 107560 49920 107720 50080
rect 107560 50080 107720 50240
rect 107560 50240 107720 50400
rect 107560 50400 107720 50560
rect 107560 50560 107720 50720
rect 107560 50720 107720 50880
rect 107560 50880 107720 51040
rect 107560 51040 107720 51200
rect 107560 51200 107720 51360
rect 107560 51360 107720 51520
rect 107560 51520 107720 51680
rect 107560 51680 107720 51840
rect 107560 51840 107720 52000
rect 107720 28320 107880 28480
rect 107720 28480 107880 28640
rect 107720 28640 107880 28800
rect 107720 28800 107880 28960
rect 107720 28960 107880 29120
rect 107720 29120 107880 29280
rect 107720 29280 107880 29440
rect 107720 29440 107880 29600
rect 107720 29600 107880 29760
rect 107720 29760 107880 29920
rect 107720 29920 107880 30080
rect 107720 30080 107880 30240
rect 107720 30240 107880 30400
rect 107720 30400 107880 30560
rect 107720 30560 107880 30720
rect 107720 30720 107880 30880
rect 107720 30880 107880 31040
rect 107720 31040 107880 31200
rect 107720 31200 107880 31360
rect 107720 31360 107880 31520
rect 107720 31520 107880 31680
rect 107720 31680 107880 31840
rect 107720 31840 107880 32000
rect 107720 32000 107880 32160
rect 107720 32160 107880 32320
rect 107720 32320 107880 32480
rect 107720 32480 107880 32640
rect 107720 32640 107880 32800
rect 107720 32800 107880 32960
rect 107720 32960 107880 33120
rect 107720 35680 107880 35840
rect 107720 35840 107880 36000
rect 107720 36000 107880 36160
rect 107720 36160 107880 36320
rect 107720 36320 107880 36480
rect 107720 36480 107880 36640
rect 107720 36640 107880 36800
rect 107720 36800 107880 36960
rect 107720 36960 107880 37120
rect 107720 37120 107880 37280
rect 107720 37280 107880 37440
rect 107720 37440 107880 37600
rect 107720 37600 107880 37760
rect 107720 37760 107880 37920
rect 107720 37920 107880 38080
rect 107720 38080 107880 38240
rect 107720 38240 107880 38400
rect 107720 38400 107880 38560
rect 107720 38560 107880 38720
rect 107720 38720 107880 38880
rect 107720 38880 107880 39040
rect 107720 39040 107880 39200
rect 107720 39200 107880 39360
rect 107720 39360 107880 39520
rect 107720 39520 107880 39680
rect 107720 39680 107880 39840
rect 107720 39840 107880 40000
rect 107720 40000 107880 40160
rect 107720 40160 107880 40320
rect 107720 40320 107880 40480
rect 107720 40480 107880 40640
rect 107720 40640 107880 40800
rect 107720 40800 107880 40960
rect 107720 40960 107880 41120
rect 107720 41120 107880 41280
rect 107720 41280 107880 41440
rect 107720 41440 107880 41600
rect 107720 41600 107880 41760
rect 107720 41760 107880 41920
rect 107720 41920 107880 42080
rect 107720 42080 107880 42240
rect 107720 42240 107880 42400
rect 107720 42400 107880 42560
rect 107720 42560 107880 42720
rect 107720 42720 107880 42880
rect 107720 42880 107880 43040
rect 107720 43040 107880 43200
rect 107720 43200 107880 43360
rect 107720 43360 107880 43520
rect 107720 43520 107880 43680
rect 107720 43680 107880 43840
rect 107720 43840 107880 44000
rect 107720 44000 107880 44160
rect 107720 47520 107880 47680
rect 107720 47680 107880 47840
rect 107720 47840 107880 48000
rect 107720 48000 107880 48160
rect 107720 48160 107880 48320
rect 107720 48320 107880 48480
rect 107720 48480 107880 48640
rect 107720 48640 107880 48800
rect 107720 48800 107880 48960
rect 107720 48960 107880 49120
rect 107720 49120 107880 49280
rect 107720 49280 107880 49440
rect 107720 49440 107880 49600
rect 107720 49600 107880 49760
rect 107720 49760 107880 49920
rect 107720 49920 107880 50080
rect 107720 50080 107880 50240
rect 107720 50240 107880 50400
rect 107720 50400 107880 50560
rect 107720 50560 107880 50720
rect 107720 50720 107880 50880
rect 107720 50880 107880 51040
rect 107720 51040 107880 51200
rect 107720 51200 107880 51360
rect 107720 51360 107880 51520
rect 107720 51520 107880 51680
rect 107880 28000 108040 28160
rect 107880 28160 108040 28320
rect 107880 28320 108040 28480
rect 107880 28480 108040 28640
rect 107880 28640 108040 28800
rect 107880 28800 108040 28960
rect 107880 28960 108040 29120
rect 107880 29120 108040 29280
rect 107880 29280 108040 29440
rect 107880 29440 108040 29600
rect 107880 29600 108040 29760
rect 107880 29760 108040 29920
rect 107880 29920 108040 30080
rect 107880 30080 108040 30240
rect 107880 30240 108040 30400
rect 107880 30400 108040 30560
rect 107880 30560 108040 30720
rect 107880 30720 108040 30880
rect 107880 30880 108040 31040
rect 107880 31040 108040 31200
rect 107880 31200 108040 31360
rect 107880 31360 108040 31520
rect 107880 31520 108040 31680
rect 107880 31680 108040 31840
rect 107880 31840 108040 32000
rect 107880 32000 108040 32160
rect 107880 32160 108040 32320
rect 107880 32320 108040 32480
rect 107880 32480 108040 32640
rect 107880 32640 108040 32800
rect 107880 32800 108040 32960
rect 107880 32960 108040 33120
rect 107880 33120 108040 33280
rect 107880 33280 108040 33440
rect 107880 33440 108040 33600
rect 107880 34880 108040 35040
rect 107880 35040 108040 35200
rect 107880 35200 108040 35360
rect 107880 35360 108040 35520
rect 107880 35520 108040 35680
rect 107880 35680 108040 35840
rect 107880 35840 108040 36000
rect 107880 36000 108040 36160
rect 107880 36160 108040 36320
rect 107880 36320 108040 36480
rect 107880 36480 108040 36640
rect 107880 36640 108040 36800
rect 107880 36800 108040 36960
rect 107880 36960 108040 37120
rect 107880 37120 108040 37280
rect 107880 37280 108040 37440
rect 107880 37440 108040 37600
rect 107880 37600 108040 37760
rect 107880 37760 108040 37920
rect 107880 37920 108040 38080
rect 107880 38080 108040 38240
rect 107880 38240 108040 38400
rect 107880 38400 108040 38560
rect 107880 38560 108040 38720
rect 107880 38720 108040 38880
rect 107880 38880 108040 39040
rect 107880 39040 108040 39200
rect 107880 39200 108040 39360
rect 107880 39360 108040 39520
rect 107880 39520 108040 39680
rect 107880 39680 108040 39840
rect 107880 39840 108040 40000
rect 107880 40000 108040 40160
rect 107880 40160 108040 40320
rect 107880 40320 108040 40480
rect 107880 40480 108040 40640
rect 107880 40640 108040 40800
rect 107880 40800 108040 40960
rect 107880 40960 108040 41120
rect 107880 41120 108040 41280
rect 107880 41280 108040 41440
rect 107880 41440 108040 41600
rect 107880 41600 108040 41760
rect 107880 41760 108040 41920
rect 107880 41920 108040 42080
rect 107880 42080 108040 42240
rect 107880 42240 108040 42400
rect 107880 42400 108040 42560
rect 107880 42560 108040 42720
rect 107880 42720 108040 42880
rect 107880 42880 108040 43040
rect 107880 43040 108040 43200
rect 107880 43200 108040 43360
rect 107880 43360 108040 43520
rect 107880 47840 108040 48000
rect 107880 48000 108040 48160
rect 107880 48160 108040 48320
rect 107880 48320 108040 48480
rect 107880 48480 108040 48640
rect 107880 48640 108040 48800
rect 107880 48800 108040 48960
rect 107880 48960 108040 49120
rect 107880 49120 108040 49280
rect 107880 49280 108040 49440
rect 107880 49440 108040 49600
rect 107880 49600 108040 49760
rect 107880 49760 108040 49920
rect 107880 49920 108040 50080
rect 107880 50080 108040 50240
rect 107880 50240 108040 50400
rect 107880 50400 108040 50560
rect 107880 50560 108040 50720
rect 107880 50720 108040 50880
rect 107880 50880 108040 51040
rect 107880 51040 108040 51200
rect 107880 51200 108040 51360
rect 107880 51360 108040 51520
rect 108040 27840 108200 28000
rect 108040 28000 108200 28160
rect 108040 28160 108200 28320
rect 108040 28320 108200 28480
rect 108040 28480 108200 28640
rect 108040 28640 108200 28800
rect 108040 28800 108200 28960
rect 108040 28960 108200 29120
rect 108040 29120 108200 29280
rect 108040 29280 108200 29440
rect 108040 29440 108200 29600
rect 108040 29600 108200 29760
rect 108040 29760 108200 29920
rect 108040 29920 108200 30080
rect 108040 30080 108200 30240
rect 108040 30240 108200 30400
rect 108040 30400 108200 30560
rect 108040 30560 108200 30720
rect 108040 30720 108200 30880
rect 108040 30880 108200 31040
rect 108040 31040 108200 31200
rect 108040 31200 108200 31360
rect 108040 31360 108200 31520
rect 108040 31520 108200 31680
rect 108040 31680 108200 31840
rect 108040 31840 108200 32000
rect 108040 32000 108200 32160
rect 108040 32160 108200 32320
rect 108040 32320 108200 32480
rect 108040 32480 108200 32640
rect 108040 32640 108200 32800
rect 108040 32800 108200 32960
rect 108040 32960 108200 33120
rect 108040 33120 108200 33280
rect 108040 33280 108200 33440
rect 108040 33440 108200 33600
rect 108040 33600 108200 33760
rect 108040 33760 108200 33920
rect 108040 33920 108200 34080
rect 108040 34080 108200 34240
rect 108040 34240 108200 34400
rect 108040 34400 108200 34560
rect 108040 34560 108200 34720
rect 108040 34720 108200 34880
rect 108040 34880 108200 35040
rect 108040 35040 108200 35200
rect 108040 35200 108200 35360
rect 108040 35360 108200 35520
rect 108040 35520 108200 35680
rect 108040 35680 108200 35840
rect 108040 35840 108200 36000
rect 108040 36000 108200 36160
rect 108040 36160 108200 36320
rect 108040 36320 108200 36480
rect 108040 36480 108200 36640
rect 108040 36640 108200 36800
rect 108040 36800 108200 36960
rect 108040 36960 108200 37120
rect 108040 37120 108200 37280
rect 108040 37280 108200 37440
rect 108040 37440 108200 37600
rect 108040 37600 108200 37760
rect 108040 37760 108200 37920
rect 108040 37920 108200 38080
rect 108040 38080 108200 38240
rect 108040 38240 108200 38400
rect 108040 38400 108200 38560
rect 108040 38560 108200 38720
rect 108040 38720 108200 38880
rect 108040 38880 108200 39040
rect 108040 39040 108200 39200
rect 108040 39200 108200 39360
rect 108040 39360 108200 39520
rect 108040 39520 108200 39680
rect 108040 39680 108200 39840
rect 108040 39840 108200 40000
rect 108040 40000 108200 40160
rect 108040 40160 108200 40320
rect 108040 40320 108200 40480
rect 108040 40480 108200 40640
rect 108040 40640 108200 40800
rect 108040 40800 108200 40960
rect 108040 40960 108200 41120
rect 108040 41120 108200 41280
rect 108040 41280 108200 41440
rect 108040 41440 108200 41600
rect 108040 41600 108200 41760
rect 108040 41760 108200 41920
rect 108040 41920 108200 42080
rect 108040 42080 108200 42240
rect 108040 42240 108200 42400
rect 108040 42400 108200 42560
rect 108040 42560 108200 42720
rect 108040 42720 108200 42880
rect 108040 42880 108200 43040
rect 108040 48160 108200 48320
rect 108040 48320 108200 48480
rect 108040 48480 108200 48640
rect 108040 48640 108200 48800
rect 108040 48800 108200 48960
rect 108040 48960 108200 49120
rect 108040 49120 108200 49280
rect 108040 49280 108200 49440
rect 108040 49440 108200 49600
rect 108040 49600 108200 49760
rect 108040 49760 108200 49920
rect 108040 49920 108200 50080
rect 108040 50080 108200 50240
rect 108040 50240 108200 50400
rect 108040 50400 108200 50560
rect 108040 50560 108200 50720
rect 108040 50720 108200 50880
rect 108040 50880 108200 51040
rect 108200 27680 108360 27840
rect 108200 27840 108360 28000
rect 108200 28000 108360 28160
rect 108200 28160 108360 28320
rect 108200 28320 108360 28480
rect 108200 28480 108360 28640
rect 108200 28640 108360 28800
rect 108200 28800 108360 28960
rect 108200 28960 108360 29120
rect 108200 29120 108360 29280
rect 108200 29280 108360 29440
rect 108200 29440 108360 29600
rect 108200 29600 108360 29760
rect 108200 29760 108360 29920
rect 108200 29920 108360 30080
rect 108200 30080 108360 30240
rect 108200 30240 108360 30400
rect 108200 30400 108360 30560
rect 108200 30560 108360 30720
rect 108200 30720 108360 30880
rect 108200 30880 108360 31040
rect 108200 31040 108360 31200
rect 108200 31200 108360 31360
rect 108200 31360 108360 31520
rect 108200 31520 108360 31680
rect 108200 31680 108360 31840
rect 108200 31840 108360 32000
rect 108200 32000 108360 32160
rect 108200 32160 108360 32320
rect 108200 32320 108360 32480
rect 108200 32480 108360 32640
rect 108200 32640 108360 32800
rect 108200 32800 108360 32960
rect 108200 32960 108360 33120
rect 108200 33120 108360 33280
rect 108200 33280 108360 33440
rect 108200 33440 108360 33600
rect 108200 33600 108360 33760
rect 108200 33760 108360 33920
rect 108200 33920 108360 34080
rect 108200 34080 108360 34240
rect 108200 34240 108360 34400
rect 108200 34400 108360 34560
rect 108200 34560 108360 34720
rect 108200 34720 108360 34880
rect 108200 34880 108360 35040
rect 108200 35040 108360 35200
rect 108200 35200 108360 35360
rect 108200 35360 108360 35520
rect 108200 35520 108360 35680
rect 108200 35680 108360 35840
rect 108200 35840 108360 36000
rect 108200 36000 108360 36160
rect 108200 36160 108360 36320
rect 108200 36320 108360 36480
rect 108200 36480 108360 36640
rect 108200 36640 108360 36800
rect 108200 36800 108360 36960
rect 108200 36960 108360 37120
rect 108200 37120 108360 37280
rect 108200 37280 108360 37440
rect 108200 37440 108360 37600
rect 108200 37600 108360 37760
rect 108200 37760 108360 37920
rect 108200 37920 108360 38080
rect 108200 38080 108360 38240
rect 108200 38240 108360 38400
rect 108200 38400 108360 38560
rect 108200 38560 108360 38720
rect 108200 38720 108360 38880
rect 108200 38880 108360 39040
rect 108200 39040 108360 39200
rect 108200 39200 108360 39360
rect 108200 39360 108360 39520
rect 108200 39520 108360 39680
rect 108200 39680 108360 39840
rect 108200 39840 108360 40000
rect 108200 40000 108360 40160
rect 108200 40160 108360 40320
rect 108200 40320 108360 40480
rect 108200 40480 108360 40640
rect 108200 40640 108360 40800
rect 108200 40800 108360 40960
rect 108200 40960 108360 41120
rect 108200 41120 108360 41280
rect 108200 41280 108360 41440
rect 108200 41440 108360 41600
rect 108200 41600 108360 41760
rect 108200 41760 108360 41920
rect 108200 41920 108360 42080
rect 108200 42080 108360 42240
rect 108200 42240 108360 42400
rect 108200 42400 108360 42560
rect 108200 48640 108360 48800
rect 108200 48800 108360 48960
rect 108200 48960 108360 49120
rect 108200 49120 108360 49280
rect 108200 49280 108360 49440
rect 108200 49440 108360 49600
rect 108200 49600 108360 49760
rect 108200 49760 108360 49920
rect 108200 49920 108360 50080
rect 108200 50080 108360 50240
rect 108200 50240 108360 50400
rect 108200 50400 108360 50560
rect 108360 27520 108520 27680
rect 108360 27680 108520 27840
rect 108360 27840 108520 28000
rect 108360 28000 108520 28160
rect 108360 28160 108520 28320
rect 108360 28320 108520 28480
rect 108360 28480 108520 28640
rect 108360 28640 108520 28800
rect 108360 28800 108520 28960
rect 108360 28960 108520 29120
rect 108360 29120 108520 29280
rect 108360 29280 108520 29440
rect 108360 29440 108520 29600
rect 108360 29600 108520 29760
rect 108360 29760 108520 29920
rect 108360 29920 108520 30080
rect 108360 30080 108520 30240
rect 108360 30240 108520 30400
rect 108360 30400 108520 30560
rect 108360 30560 108520 30720
rect 108360 30720 108520 30880
rect 108360 30880 108520 31040
rect 108360 31040 108520 31200
rect 108360 31200 108520 31360
rect 108360 31360 108520 31520
rect 108360 31520 108520 31680
rect 108360 31680 108520 31840
rect 108360 31840 108520 32000
rect 108360 32000 108520 32160
rect 108360 32160 108520 32320
rect 108360 32320 108520 32480
rect 108360 32480 108520 32640
rect 108360 32640 108520 32800
rect 108360 32800 108520 32960
rect 108360 32960 108520 33120
rect 108360 33120 108520 33280
rect 108360 33280 108520 33440
rect 108360 33440 108520 33600
rect 108360 33600 108520 33760
rect 108360 33760 108520 33920
rect 108360 33920 108520 34080
rect 108360 34080 108520 34240
rect 108360 34240 108520 34400
rect 108360 34400 108520 34560
rect 108360 34560 108520 34720
rect 108360 34720 108520 34880
rect 108360 34880 108520 35040
rect 108360 35040 108520 35200
rect 108360 35200 108520 35360
rect 108360 35360 108520 35520
rect 108360 35520 108520 35680
rect 108360 35680 108520 35840
rect 108360 35840 108520 36000
rect 108360 36000 108520 36160
rect 108360 36160 108520 36320
rect 108360 36320 108520 36480
rect 108360 36480 108520 36640
rect 108360 36640 108520 36800
rect 108360 36800 108520 36960
rect 108360 36960 108520 37120
rect 108360 37120 108520 37280
rect 108360 37280 108520 37440
rect 108360 37440 108520 37600
rect 108360 37600 108520 37760
rect 108360 37760 108520 37920
rect 108360 37920 108520 38080
rect 108360 38080 108520 38240
rect 108360 38240 108520 38400
rect 108360 38400 108520 38560
rect 108360 38560 108520 38720
rect 108360 38720 108520 38880
rect 108360 38880 108520 39040
rect 108360 39040 108520 39200
rect 108360 39200 108520 39360
rect 108360 39360 108520 39520
rect 108360 39520 108520 39680
rect 108360 39680 108520 39840
rect 108360 39840 108520 40000
rect 108360 40000 108520 40160
rect 108360 40160 108520 40320
rect 108360 40320 108520 40480
rect 108360 40480 108520 40640
rect 108360 40640 108520 40800
rect 108360 40800 108520 40960
rect 108360 40960 108520 41120
rect 108360 41120 108520 41280
rect 108360 41280 108520 41440
rect 108360 41440 108520 41600
rect 108360 41600 108520 41760
rect 108360 41760 108520 41920
rect 108360 41920 108520 42080
rect 108520 27360 108680 27520
rect 108520 27520 108680 27680
rect 108520 27680 108680 27840
rect 108520 27840 108680 28000
rect 108520 28000 108680 28160
rect 108520 28160 108680 28320
rect 108520 28320 108680 28480
rect 108520 28480 108680 28640
rect 108520 28640 108680 28800
rect 108520 28800 108680 28960
rect 108520 28960 108680 29120
rect 108520 29120 108680 29280
rect 108520 29280 108680 29440
rect 108520 29440 108680 29600
rect 108520 29600 108680 29760
rect 108520 29760 108680 29920
rect 108520 29920 108680 30080
rect 108520 30080 108680 30240
rect 108520 30240 108680 30400
rect 108520 30400 108680 30560
rect 108520 30560 108680 30720
rect 108520 30720 108680 30880
rect 108520 30880 108680 31040
rect 108520 31040 108680 31200
rect 108520 31200 108680 31360
rect 108520 31360 108680 31520
rect 108520 31520 108680 31680
rect 108520 31680 108680 31840
rect 108520 31840 108680 32000
rect 108520 32000 108680 32160
rect 108520 32160 108680 32320
rect 108520 32320 108680 32480
rect 108520 32480 108680 32640
rect 108520 32640 108680 32800
rect 108520 32800 108680 32960
rect 108520 32960 108680 33120
rect 108520 33120 108680 33280
rect 108520 33280 108680 33440
rect 108520 33440 108680 33600
rect 108520 33600 108680 33760
rect 108520 33760 108680 33920
rect 108520 33920 108680 34080
rect 108520 34080 108680 34240
rect 108520 34240 108680 34400
rect 108520 34400 108680 34560
rect 108520 34560 108680 34720
rect 108520 34720 108680 34880
rect 108520 34880 108680 35040
rect 108520 35040 108680 35200
rect 108520 35200 108680 35360
rect 108520 35360 108680 35520
rect 108520 35520 108680 35680
rect 108520 35680 108680 35840
rect 108520 35840 108680 36000
rect 108520 36000 108680 36160
rect 108520 36160 108680 36320
rect 108520 36320 108680 36480
rect 108520 36480 108680 36640
rect 108520 36640 108680 36800
rect 108520 36800 108680 36960
rect 108520 36960 108680 37120
rect 108520 37120 108680 37280
rect 108520 37280 108680 37440
rect 108520 37440 108680 37600
rect 108520 37600 108680 37760
rect 108520 37760 108680 37920
rect 108520 37920 108680 38080
rect 108520 38080 108680 38240
rect 108520 38240 108680 38400
rect 108520 38400 108680 38560
rect 108520 38560 108680 38720
rect 108520 38720 108680 38880
rect 108520 38880 108680 39040
rect 108520 39040 108680 39200
rect 108520 39200 108680 39360
rect 108520 39360 108680 39520
rect 108520 39520 108680 39680
rect 108520 39680 108680 39840
rect 108520 39840 108680 40000
rect 108520 40000 108680 40160
rect 108520 40160 108680 40320
rect 108520 40320 108680 40480
rect 108520 40480 108680 40640
rect 108520 40640 108680 40800
rect 108520 40800 108680 40960
rect 108520 40960 108680 41120
rect 108520 41120 108680 41280
rect 108520 41280 108680 41440
rect 108520 41440 108680 41600
rect 108680 27200 108840 27360
rect 108680 27360 108840 27520
rect 108680 27520 108840 27680
rect 108680 27680 108840 27840
rect 108680 27840 108840 28000
rect 108680 28000 108840 28160
rect 108680 28160 108840 28320
rect 108680 28320 108840 28480
rect 108680 28480 108840 28640
rect 108680 28640 108840 28800
rect 108680 28800 108840 28960
rect 108680 28960 108840 29120
rect 108680 29120 108840 29280
rect 108680 29280 108840 29440
rect 108680 29440 108840 29600
rect 108680 29600 108840 29760
rect 108680 29760 108840 29920
rect 108680 29920 108840 30080
rect 108680 30080 108840 30240
rect 108680 30240 108840 30400
rect 108680 30400 108840 30560
rect 108680 30560 108840 30720
rect 108680 30720 108840 30880
rect 108680 30880 108840 31040
rect 108680 31040 108840 31200
rect 108680 31200 108840 31360
rect 108680 31360 108840 31520
rect 108680 31520 108840 31680
rect 108680 31680 108840 31840
rect 108680 31840 108840 32000
rect 108680 32000 108840 32160
rect 108680 32160 108840 32320
rect 108680 32320 108840 32480
rect 108680 32480 108840 32640
rect 108680 32640 108840 32800
rect 108680 32800 108840 32960
rect 108680 32960 108840 33120
rect 108680 33120 108840 33280
rect 108680 33280 108840 33440
rect 108680 33440 108840 33600
rect 108680 33600 108840 33760
rect 108680 33760 108840 33920
rect 108680 33920 108840 34080
rect 108680 34080 108840 34240
rect 108680 34240 108840 34400
rect 108680 34400 108840 34560
rect 108680 34560 108840 34720
rect 108680 34720 108840 34880
rect 108680 34880 108840 35040
rect 108680 35040 108840 35200
rect 108680 35200 108840 35360
rect 108680 35360 108840 35520
rect 108680 35520 108840 35680
rect 108680 35680 108840 35840
rect 108680 35840 108840 36000
rect 108680 36000 108840 36160
rect 108680 36160 108840 36320
rect 108680 36320 108840 36480
rect 108680 36480 108840 36640
rect 108680 36640 108840 36800
rect 108680 36800 108840 36960
rect 108680 36960 108840 37120
rect 108680 37120 108840 37280
rect 108680 37280 108840 37440
rect 108680 37440 108840 37600
rect 108680 37600 108840 37760
rect 108680 37760 108840 37920
rect 108680 37920 108840 38080
rect 108680 38080 108840 38240
rect 108680 38240 108840 38400
rect 108680 38400 108840 38560
rect 108680 38560 108840 38720
rect 108680 38720 108840 38880
rect 108680 38880 108840 39040
rect 108680 39040 108840 39200
rect 108680 39200 108840 39360
rect 108680 39360 108840 39520
rect 108680 39520 108840 39680
rect 108680 39680 108840 39840
rect 108680 39840 108840 40000
rect 108680 40000 108840 40160
rect 108680 40160 108840 40320
rect 108680 40320 108840 40480
rect 108680 40480 108840 40640
rect 108680 40640 108840 40800
rect 108680 40800 108840 40960
rect 108680 40960 108840 41120
rect 108840 27200 109000 27360
rect 108840 27360 109000 27520
rect 108840 27520 109000 27680
rect 108840 27680 109000 27840
rect 108840 27840 109000 28000
rect 108840 28000 109000 28160
rect 108840 28160 109000 28320
rect 108840 28320 109000 28480
rect 108840 28480 109000 28640
rect 108840 28640 109000 28800
rect 108840 28800 109000 28960
rect 108840 28960 109000 29120
rect 108840 29120 109000 29280
rect 108840 29280 109000 29440
rect 108840 29440 109000 29600
rect 108840 29600 109000 29760
rect 108840 29760 109000 29920
rect 108840 29920 109000 30080
rect 108840 30080 109000 30240
rect 108840 30240 109000 30400
rect 108840 30400 109000 30560
rect 108840 30560 109000 30720
rect 108840 30720 109000 30880
rect 108840 30880 109000 31040
rect 108840 31040 109000 31200
rect 108840 31200 109000 31360
rect 108840 31360 109000 31520
rect 108840 31520 109000 31680
rect 108840 31680 109000 31840
rect 108840 31840 109000 32000
rect 108840 32000 109000 32160
rect 108840 32160 109000 32320
rect 108840 32320 109000 32480
rect 108840 32480 109000 32640
rect 108840 32640 109000 32800
rect 108840 32800 109000 32960
rect 108840 32960 109000 33120
rect 108840 33120 109000 33280
rect 108840 33280 109000 33440
rect 108840 33440 109000 33600
rect 108840 33600 109000 33760
rect 108840 33760 109000 33920
rect 108840 33920 109000 34080
rect 108840 34080 109000 34240
rect 108840 34240 109000 34400
rect 108840 34400 109000 34560
rect 108840 34560 109000 34720
rect 108840 34720 109000 34880
rect 108840 34880 109000 35040
rect 108840 35040 109000 35200
rect 108840 35200 109000 35360
rect 108840 35360 109000 35520
rect 108840 35520 109000 35680
rect 108840 35680 109000 35840
rect 108840 35840 109000 36000
rect 108840 36000 109000 36160
rect 108840 36160 109000 36320
rect 108840 36320 109000 36480
rect 108840 36480 109000 36640
rect 108840 36640 109000 36800
rect 108840 36800 109000 36960
rect 108840 36960 109000 37120
rect 108840 37120 109000 37280
rect 108840 37280 109000 37440
rect 108840 37440 109000 37600
rect 108840 37600 109000 37760
rect 108840 37760 109000 37920
rect 108840 37920 109000 38080
rect 108840 38080 109000 38240
rect 108840 38240 109000 38400
rect 108840 38400 109000 38560
rect 108840 38560 109000 38720
rect 108840 38720 109000 38880
rect 108840 38880 109000 39040
rect 108840 39040 109000 39200
rect 108840 39200 109000 39360
rect 108840 39360 109000 39520
rect 108840 39520 109000 39680
rect 108840 39680 109000 39840
rect 108840 39840 109000 40000
rect 108840 40000 109000 40160
rect 108840 40160 109000 40320
rect 108840 40320 109000 40480
rect 108840 40480 109000 40640
rect 109000 27040 109160 27200
rect 109000 27200 109160 27360
rect 109000 27360 109160 27520
rect 109000 27520 109160 27680
rect 109000 27680 109160 27840
rect 109000 27840 109160 28000
rect 109000 28000 109160 28160
rect 109000 28160 109160 28320
rect 109000 28320 109160 28480
rect 109000 28480 109160 28640
rect 109000 28640 109160 28800
rect 109000 28800 109160 28960
rect 109000 28960 109160 29120
rect 109000 29120 109160 29280
rect 109000 29280 109160 29440
rect 109000 29440 109160 29600
rect 109000 29600 109160 29760
rect 109000 29760 109160 29920
rect 109000 29920 109160 30080
rect 109000 30080 109160 30240
rect 109000 30240 109160 30400
rect 109000 30400 109160 30560
rect 109000 30560 109160 30720
rect 109000 30720 109160 30880
rect 109000 30880 109160 31040
rect 109000 31040 109160 31200
rect 109000 31200 109160 31360
rect 109000 31360 109160 31520
rect 109000 31520 109160 31680
rect 109000 31680 109160 31840
rect 109000 31840 109160 32000
rect 109000 32000 109160 32160
rect 109000 32160 109160 32320
rect 109000 32320 109160 32480
rect 109000 32480 109160 32640
rect 109000 32640 109160 32800
rect 109000 32800 109160 32960
rect 109000 32960 109160 33120
rect 109000 33120 109160 33280
rect 109000 33280 109160 33440
rect 109000 33440 109160 33600
rect 109000 33600 109160 33760
rect 109000 33760 109160 33920
rect 109000 33920 109160 34080
rect 109000 34080 109160 34240
rect 109000 34240 109160 34400
rect 109000 34400 109160 34560
rect 109000 34560 109160 34720
rect 109000 34720 109160 34880
rect 109000 34880 109160 35040
rect 109000 35040 109160 35200
rect 109000 35200 109160 35360
rect 109000 35360 109160 35520
rect 109000 35520 109160 35680
rect 109000 35680 109160 35840
rect 109000 35840 109160 36000
rect 109000 36000 109160 36160
rect 109000 36160 109160 36320
rect 109000 36320 109160 36480
rect 109000 36480 109160 36640
rect 109000 36640 109160 36800
rect 109000 36800 109160 36960
rect 109000 36960 109160 37120
rect 109000 37120 109160 37280
rect 109000 37280 109160 37440
rect 109000 37440 109160 37600
rect 109000 37600 109160 37760
rect 109000 37760 109160 37920
rect 109000 37920 109160 38080
rect 109000 38080 109160 38240
rect 109000 38240 109160 38400
rect 109000 38400 109160 38560
rect 109000 38560 109160 38720
rect 109000 38720 109160 38880
rect 109000 38880 109160 39040
rect 109000 39040 109160 39200
rect 109000 39200 109160 39360
rect 109000 39360 109160 39520
rect 109000 39520 109160 39680
rect 109000 39680 109160 39840
rect 109000 39840 109160 40000
rect 109000 40000 109160 40160
rect 109160 27040 109320 27200
rect 109160 27200 109320 27360
rect 109160 27360 109320 27520
rect 109160 27520 109320 27680
rect 109160 27680 109320 27840
rect 109160 27840 109320 28000
rect 109160 28000 109320 28160
rect 109160 28160 109320 28320
rect 109160 28320 109320 28480
rect 109160 28480 109320 28640
rect 109160 28640 109320 28800
rect 109160 28800 109320 28960
rect 109160 28960 109320 29120
rect 109160 29120 109320 29280
rect 109160 29280 109320 29440
rect 109160 29440 109320 29600
rect 109160 29600 109320 29760
rect 109160 29760 109320 29920
rect 109160 29920 109320 30080
rect 109160 30080 109320 30240
rect 109160 30240 109320 30400
rect 109160 30400 109320 30560
rect 109160 30560 109320 30720
rect 109160 30720 109320 30880
rect 109160 30880 109320 31040
rect 109160 31040 109320 31200
rect 109160 31200 109320 31360
rect 109160 31360 109320 31520
rect 109160 31520 109320 31680
rect 109160 31680 109320 31840
rect 109160 31840 109320 32000
rect 109160 32000 109320 32160
rect 109160 32160 109320 32320
rect 109160 32320 109320 32480
rect 109160 32480 109320 32640
rect 109160 32640 109320 32800
rect 109160 32800 109320 32960
rect 109160 32960 109320 33120
rect 109160 33120 109320 33280
rect 109160 33280 109320 33440
rect 109160 33440 109320 33600
rect 109160 33600 109320 33760
rect 109160 33760 109320 33920
rect 109160 33920 109320 34080
rect 109160 34080 109320 34240
rect 109160 34240 109320 34400
rect 109160 34400 109320 34560
rect 109160 34560 109320 34720
rect 109160 34720 109320 34880
rect 109160 34880 109320 35040
rect 109160 35040 109320 35200
rect 109160 35200 109320 35360
rect 109160 35360 109320 35520
rect 109160 35520 109320 35680
rect 109160 35680 109320 35840
rect 109160 35840 109320 36000
rect 109160 36000 109320 36160
rect 109160 36160 109320 36320
rect 109160 36320 109320 36480
rect 109160 36480 109320 36640
rect 109160 36640 109320 36800
rect 109160 36800 109320 36960
rect 109160 36960 109320 37120
rect 109160 37120 109320 37280
rect 109160 37280 109320 37440
rect 109160 37440 109320 37600
rect 109160 37600 109320 37760
rect 109160 37760 109320 37920
rect 109160 37920 109320 38080
rect 109160 38080 109320 38240
rect 109160 38240 109320 38400
rect 109160 38400 109320 38560
rect 109160 38560 109320 38720
rect 109160 38720 109320 38880
rect 109160 38880 109320 39040
rect 109160 39040 109320 39200
rect 109160 39200 109320 39360
rect 109160 39360 109320 39520
rect 109160 39520 109320 39680
rect 109320 27040 109480 27200
rect 109320 27200 109480 27360
rect 109320 27360 109480 27520
rect 109320 27520 109480 27680
rect 109320 27680 109480 27840
rect 109320 27840 109480 28000
rect 109320 28000 109480 28160
rect 109320 28160 109480 28320
rect 109320 28320 109480 28480
rect 109320 28480 109480 28640
rect 109320 28640 109480 28800
rect 109320 28800 109480 28960
rect 109320 28960 109480 29120
rect 109320 29120 109480 29280
rect 109320 29280 109480 29440
rect 109320 29440 109480 29600
rect 109320 29600 109480 29760
rect 109320 29760 109480 29920
rect 109320 29920 109480 30080
rect 109320 30080 109480 30240
rect 109320 30240 109480 30400
rect 109320 30400 109480 30560
rect 109320 30560 109480 30720
rect 109320 30720 109480 30880
rect 109320 30880 109480 31040
rect 109320 31040 109480 31200
rect 109320 31200 109480 31360
rect 109320 31360 109480 31520
rect 109320 31520 109480 31680
rect 109320 31680 109480 31840
rect 109320 31840 109480 32000
rect 109320 32000 109480 32160
rect 109320 32160 109480 32320
rect 109320 32320 109480 32480
rect 109320 32480 109480 32640
rect 109320 32640 109480 32800
rect 109320 32800 109480 32960
rect 109320 32960 109480 33120
rect 109320 33120 109480 33280
rect 109320 33280 109480 33440
rect 109320 33440 109480 33600
rect 109320 33600 109480 33760
rect 109320 33760 109480 33920
rect 109320 33920 109480 34080
rect 109320 34080 109480 34240
rect 109320 34240 109480 34400
rect 109320 34400 109480 34560
rect 109320 34560 109480 34720
rect 109320 34720 109480 34880
rect 109320 34880 109480 35040
rect 109320 35040 109480 35200
rect 109320 35200 109480 35360
rect 109320 35360 109480 35520
rect 109320 35520 109480 35680
rect 109320 35680 109480 35840
rect 109320 35840 109480 36000
rect 109320 36000 109480 36160
rect 109320 36160 109480 36320
rect 109320 36320 109480 36480
rect 109320 36480 109480 36640
rect 109320 36640 109480 36800
rect 109320 36800 109480 36960
rect 109320 36960 109480 37120
rect 109320 37120 109480 37280
rect 109320 37280 109480 37440
rect 109320 37440 109480 37600
rect 109320 37600 109480 37760
rect 109320 37760 109480 37920
rect 109320 37920 109480 38080
rect 109320 38080 109480 38240
rect 109320 38240 109480 38400
rect 109320 38400 109480 38560
rect 109320 38560 109480 38720
rect 109320 38720 109480 38880
rect 109320 38880 109480 39040
rect 109320 39040 109480 39200
rect 109320 39200 109480 39360
rect 109480 26880 109640 27040
rect 109480 27040 109640 27200
rect 109480 27200 109640 27360
rect 109480 27360 109640 27520
rect 109480 27520 109640 27680
rect 109480 27680 109640 27840
rect 109480 27840 109640 28000
rect 109480 28000 109640 28160
rect 109480 28160 109640 28320
rect 109480 28320 109640 28480
rect 109480 28480 109640 28640
rect 109480 28640 109640 28800
rect 109480 28800 109640 28960
rect 109480 28960 109640 29120
rect 109480 29120 109640 29280
rect 109480 29280 109640 29440
rect 109480 29440 109640 29600
rect 109480 29600 109640 29760
rect 109480 29760 109640 29920
rect 109480 29920 109640 30080
rect 109480 30080 109640 30240
rect 109480 30240 109640 30400
rect 109480 30400 109640 30560
rect 109480 30560 109640 30720
rect 109480 30720 109640 30880
rect 109480 30880 109640 31040
rect 109480 31040 109640 31200
rect 109480 31200 109640 31360
rect 109480 31360 109640 31520
rect 109480 31520 109640 31680
rect 109480 31680 109640 31840
rect 109480 31840 109640 32000
rect 109480 32000 109640 32160
rect 109480 32160 109640 32320
rect 109480 32320 109640 32480
rect 109480 32480 109640 32640
rect 109480 32640 109640 32800
rect 109480 32800 109640 32960
rect 109480 32960 109640 33120
rect 109480 33120 109640 33280
rect 109480 33280 109640 33440
rect 109480 33440 109640 33600
rect 109480 33600 109640 33760
rect 109480 33760 109640 33920
rect 109480 33920 109640 34080
rect 109480 34080 109640 34240
rect 109480 34240 109640 34400
rect 109480 34400 109640 34560
rect 109480 34560 109640 34720
rect 109480 34720 109640 34880
rect 109480 34880 109640 35040
rect 109480 35040 109640 35200
rect 109480 35200 109640 35360
rect 109480 35360 109640 35520
rect 109480 35520 109640 35680
rect 109480 35680 109640 35840
rect 109480 35840 109640 36000
rect 109480 36000 109640 36160
rect 109480 36160 109640 36320
rect 109480 36320 109640 36480
rect 109480 36480 109640 36640
rect 109480 36640 109640 36800
rect 109480 36800 109640 36960
rect 109480 36960 109640 37120
rect 109480 37120 109640 37280
rect 109480 37280 109640 37440
rect 109480 37440 109640 37600
rect 109480 37600 109640 37760
rect 109480 37760 109640 37920
rect 109480 37920 109640 38080
rect 109480 38080 109640 38240
rect 109480 38240 109640 38400
rect 109480 38400 109640 38560
rect 109480 38560 109640 38720
rect 109480 38720 109640 38880
rect 109640 26880 109800 27040
rect 109640 27040 109800 27200
rect 109640 27200 109800 27360
rect 109640 27360 109800 27520
rect 109640 27520 109800 27680
rect 109640 27680 109800 27840
rect 109640 27840 109800 28000
rect 109640 28000 109800 28160
rect 109640 28160 109800 28320
rect 109640 28320 109800 28480
rect 109640 28480 109800 28640
rect 109640 28640 109800 28800
rect 109640 28800 109800 28960
rect 109640 28960 109800 29120
rect 109640 29120 109800 29280
rect 109640 29280 109800 29440
rect 109640 29440 109800 29600
rect 109640 29600 109800 29760
rect 109640 29760 109800 29920
rect 109640 29920 109800 30080
rect 109640 30080 109800 30240
rect 109640 30240 109800 30400
rect 109640 30880 109800 31040
rect 109640 31040 109800 31200
rect 109640 31200 109800 31360
rect 109640 31360 109800 31520
rect 109640 31520 109800 31680
rect 109640 31680 109800 31840
rect 109640 31840 109800 32000
rect 109640 32000 109800 32160
rect 109640 32160 109800 32320
rect 109640 32320 109800 32480
rect 109640 32480 109800 32640
rect 109640 32640 109800 32800
rect 109640 32800 109800 32960
rect 109640 32960 109800 33120
rect 109640 33120 109800 33280
rect 109640 33280 109800 33440
rect 109640 33440 109800 33600
rect 109640 33600 109800 33760
rect 109640 33760 109800 33920
rect 109640 33920 109800 34080
rect 109640 34080 109800 34240
rect 109640 34240 109800 34400
rect 109640 34400 109800 34560
rect 109640 34560 109800 34720
rect 109640 34720 109800 34880
rect 109640 34880 109800 35040
rect 109640 35040 109800 35200
rect 109640 35200 109800 35360
rect 109640 35360 109800 35520
rect 109640 35520 109800 35680
rect 109640 35680 109800 35840
rect 109640 35840 109800 36000
rect 109640 36000 109800 36160
rect 109640 36160 109800 36320
rect 109640 36320 109800 36480
rect 109640 36480 109800 36640
rect 109640 36640 109800 36800
rect 109640 36800 109800 36960
rect 109640 36960 109800 37120
rect 109640 37120 109800 37280
rect 109640 37280 109800 37440
rect 109640 37440 109800 37600
rect 109640 37600 109800 37760
rect 109640 37760 109800 37920
rect 109640 37920 109800 38080
rect 109640 38080 109800 38240
rect 109640 38240 109800 38400
rect 109800 26880 109960 27040
rect 109800 27040 109960 27200
rect 109800 27200 109960 27360
rect 109800 27360 109960 27520
rect 109800 27520 109960 27680
rect 109800 27680 109960 27840
rect 109800 27840 109960 28000
rect 109800 28000 109960 28160
rect 109800 28160 109960 28320
rect 109800 28320 109960 28480
rect 109800 28480 109960 28640
rect 109800 28640 109960 28800
rect 109800 28800 109960 28960
rect 109800 28960 109960 29120
rect 109800 29120 109960 29280
rect 109800 29280 109960 29440
rect 109800 29440 109960 29600
rect 109800 29600 109960 29760
rect 109800 29760 109960 29920
rect 109800 31360 109960 31520
rect 109800 31520 109960 31680
rect 109800 31680 109960 31840
rect 109800 31840 109960 32000
rect 109800 32000 109960 32160
rect 109800 32160 109960 32320
rect 109800 32320 109960 32480
rect 109800 32480 109960 32640
rect 109800 32640 109960 32800
rect 109800 32800 109960 32960
rect 109800 32960 109960 33120
rect 109800 33120 109960 33280
rect 109800 33280 109960 33440
rect 109800 33440 109960 33600
rect 109800 33600 109960 33760
rect 109800 33760 109960 33920
rect 109800 33920 109960 34080
rect 109800 34080 109960 34240
rect 109800 34240 109960 34400
rect 109800 34400 109960 34560
rect 109800 34560 109960 34720
rect 109800 34720 109960 34880
rect 109800 34880 109960 35040
rect 109800 35040 109960 35200
rect 109800 35200 109960 35360
rect 109800 35360 109960 35520
rect 109800 35520 109960 35680
rect 109800 35680 109960 35840
rect 109800 35840 109960 36000
rect 109800 36000 109960 36160
rect 109800 36160 109960 36320
rect 109800 36320 109960 36480
rect 109800 36480 109960 36640
rect 109800 36640 109960 36800
rect 109800 36800 109960 36960
rect 109800 36960 109960 37120
rect 109800 37120 109960 37280
rect 109800 37280 109960 37440
rect 109800 37440 109960 37600
rect 109800 37600 109960 37760
rect 109800 37760 109960 37920
rect 109960 26880 110120 27040
rect 109960 27040 110120 27200
rect 109960 27200 110120 27360
rect 109960 27360 110120 27520
rect 109960 27520 110120 27680
rect 109960 27680 110120 27840
rect 109960 27840 110120 28000
rect 109960 28000 110120 28160
rect 109960 28160 110120 28320
rect 109960 28320 110120 28480
rect 109960 28480 110120 28640
rect 109960 28640 110120 28800
rect 109960 28800 110120 28960
rect 109960 28960 110120 29120
rect 109960 29120 110120 29280
rect 109960 29280 110120 29440
rect 109960 29440 110120 29600
rect 109960 29600 110120 29760
rect 109960 31680 110120 31840
rect 109960 31840 110120 32000
rect 109960 32000 110120 32160
rect 109960 32160 110120 32320
rect 109960 32320 110120 32480
rect 109960 32480 110120 32640
rect 109960 32640 110120 32800
rect 109960 32800 110120 32960
rect 109960 32960 110120 33120
rect 109960 33120 110120 33280
rect 109960 33280 110120 33440
rect 109960 33440 110120 33600
rect 109960 33600 110120 33760
rect 109960 33760 110120 33920
rect 109960 33920 110120 34080
rect 109960 34080 110120 34240
rect 109960 34240 110120 34400
rect 109960 34400 110120 34560
rect 109960 34560 110120 34720
rect 109960 34720 110120 34880
rect 109960 34880 110120 35040
rect 109960 35040 110120 35200
rect 109960 35200 110120 35360
rect 109960 35360 110120 35520
rect 109960 35520 110120 35680
rect 109960 35680 110120 35840
rect 109960 35840 110120 36000
rect 109960 36000 110120 36160
rect 109960 36160 110120 36320
rect 109960 36320 110120 36480
rect 109960 36480 110120 36640
rect 109960 36640 110120 36800
rect 109960 36800 110120 36960
rect 109960 36960 110120 37120
rect 109960 37120 110120 37280
rect 109960 37280 110120 37440
rect 109960 37440 110120 37600
rect 110120 26720 110280 26880
rect 110120 26880 110280 27040
rect 110120 27040 110280 27200
rect 110120 27200 110280 27360
rect 110120 27360 110280 27520
rect 110120 27520 110280 27680
rect 110120 27680 110280 27840
rect 110120 27840 110280 28000
rect 110120 28000 110280 28160
rect 110120 28160 110280 28320
rect 110120 28320 110280 28480
rect 110120 28480 110280 28640
rect 110120 28640 110280 28800
rect 110120 28800 110280 28960
rect 110120 28960 110280 29120
rect 110120 29120 110280 29280
rect 110120 29280 110280 29440
rect 110120 29440 110280 29600
rect 110120 31840 110280 32000
rect 110120 32000 110280 32160
rect 110120 32160 110280 32320
rect 110120 32320 110280 32480
rect 110120 32480 110280 32640
rect 110120 32640 110280 32800
rect 110120 32800 110280 32960
rect 110120 32960 110280 33120
rect 110120 33120 110280 33280
rect 110120 33280 110280 33440
rect 110120 33440 110280 33600
rect 110120 33600 110280 33760
rect 110120 33760 110280 33920
rect 110120 33920 110280 34080
rect 110120 34080 110280 34240
rect 110120 34240 110280 34400
rect 110120 34400 110280 34560
rect 110120 34560 110280 34720
rect 110120 34720 110280 34880
rect 110120 34880 110280 35040
rect 110120 35040 110280 35200
rect 110120 35200 110280 35360
rect 110120 35360 110280 35520
rect 110120 35520 110280 35680
rect 110120 35680 110280 35840
rect 110120 35840 110280 36000
rect 110120 36000 110280 36160
rect 110120 36160 110280 36320
rect 110120 36320 110280 36480
rect 110120 36480 110280 36640
rect 110120 36640 110280 36800
rect 110120 36800 110280 36960
rect 110120 36960 110280 37120
rect 110280 26720 110440 26880
rect 110280 26880 110440 27040
rect 110280 27040 110440 27200
rect 110280 27200 110440 27360
rect 110280 27360 110440 27520
rect 110280 27520 110440 27680
rect 110280 27680 110440 27840
rect 110280 27840 110440 28000
rect 110280 28000 110440 28160
rect 110280 28160 110440 28320
rect 110280 28320 110440 28480
rect 110280 28480 110440 28640
rect 110280 28640 110440 28800
rect 110280 28800 110440 28960
rect 110280 28960 110440 29120
rect 110280 29120 110440 29280
rect 110280 29280 110440 29440
rect 110280 31840 110440 32000
rect 110280 32000 110440 32160
rect 110280 32160 110440 32320
rect 110280 32320 110440 32480
rect 110280 32480 110440 32640
rect 110280 32640 110440 32800
rect 110280 32800 110440 32960
rect 110280 32960 110440 33120
rect 110280 33120 110440 33280
rect 110280 33280 110440 33440
rect 110280 33440 110440 33600
rect 110280 33600 110440 33760
rect 110280 33760 110440 33920
rect 110280 33920 110440 34080
rect 110280 34080 110440 34240
rect 110280 34240 110440 34400
rect 110280 34400 110440 34560
rect 110280 34560 110440 34720
rect 110280 34720 110440 34880
rect 110280 34880 110440 35040
rect 110280 35040 110440 35200
rect 110280 35200 110440 35360
rect 110280 35360 110440 35520
rect 110280 35520 110440 35680
rect 110280 35680 110440 35840
rect 110280 35840 110440 36000
rect 110280 36000 110440 36160
rect 110280 36160 110440 36320
rect 110280 36320 110440 36480
rect 110280 36480 110440 36640
rect 110280 36640 110440 36800
rect 110440 26720 110600 26880
rect 110440 26880 110600 27040
rect 110440 27040 110600 27200
rect 110440 27200 110600 27360
rect 110440 27360 110600 27520
rect 110440 27520 110600 27680
rect 110440 27680 110600 27840
rect 110440 27840 110600 28000
rect 110440 28000 110600 28160
rect 110440 28160 110600 28320
rect 110440 28320 110600 28480
rect 110440 28480 110600 28640
rect 110440 28640 110600 28800
rect 110440 28800 110600 28960
rect 110440 28960 110600 29120
rect 110440 29120 110600 29280
rect 110440 29280 110600 29440
rect 110440 31840 110600 32000
rect 110440 32000 110600 32160
rect 110440 32160 110600 32320
rect 110440 32320 110600 32480
rect 110440 32480 110600 32640
rect 110440 32640 110600 32800
rect 110440 32800 110600 32960
rect 110440 32960 110600 33120
rect 110440 33120 110600 33280
rect 110440 33280 110600 33440
rect 110440 33440 110600 33600
rect 110440 33600 110600 33760
rect 110440 33760 110600 33920
rect 110440 33920 110600 34080
rect 110440 34080 110600 34240
rect 110440 34240 110600 34400
rect 110440 34400 110600 34560
rect 110440 34560 110600 34720
rect 110440 34720 110600 34880
rect 110440 34880 110600 35040
rect 110440 35040 110600 35200
rect 110440 35200 110600 35360
rect 110440 35360 110600 35520
rect 110440 35520 110600 35680
rect 110440 35680 110600 35840
rect 110440 35840 110600 36000
rect 110440 36000 110600 36160
rect 110440 36160 110600 36320
rect 110600 26720 110760 26880
rect 110600 26880 110760 27040
rect 110600 27040 110760 27200
rect 110600 27200 110760 27360
rect 110600 27360 110760 27520
rect 110600 27520 110760 27680
rect 110600 27680 110760 27840
rect 110600 27840 110760 28000
rect 110600 28000 110760 28160
rect 110600 28160 110760 28320
rect 110600 28320 110760 28480
rect 110600 28480 110760 28640
rect 110600 28640 110760 28800
rect 110600 28800 110760 28960
rect 110600 28960 110760 29120
rect 110600 29120 110760 29280
rect 110600 29280 110760 29440
rect 110600 31840 110760 32000
rect 110600 32000 110760 32160
rect 110600 32160 110760 32320
rect 110600 32320 110760 32480
rect 110600 32480 110760 32640
rect 110600 32640 110760 32800
rect 110600 32800 110760 32960
rect 110600 32960 110760 33120
rect 110600 33120 110760 33280
rect 110600 33280 110760 33440
rect 110600 33440 110760 33600
rect 110600 33600 110760 33760
rect 110600 33760 110760 33920
rect 110600 33920 110760 34080
rect 110600 34080 110760 34240
rect 110600 34240 110760 34400
rect 110600 34400 110760 34560
rect 110600 34560 110760 34720
rect 110600 34720 110760 34880
rect 110600 34880 110760 35040
rect 110600 35040 110760 35200
rect 110600 35200 110760 35360
rect 110600 35360 110760 35520
rect 110600 35520 110760 35680
rect 110600 35680 110760 35840
rect 110600 35840 110760 36000
rect 110760 26720 110920 26880
rect 110760 26880 110920 27040
rect 110760 27040 110920 27200
rect 110760 27200 110920 27360
rect 110760 27360 110920 27520
rect 110760 27520 110920 27680
rect 110760 27680 110920 27840
rect 110760 27840 110920 28000
rect 110760 28000 110920 28160
rect 110760 28160 110920 28320
rect 110760 28320 110920 28480
rect 110760 28480 110920 28640
rect 110760 28640 110920 28800
rect 110760 28800 110920 28960
rect 110760 28960 110920 29120
rect 110760 29120 110920 29280
rect 110760 31840 110920 32000
rect 110760 32000 110920 32160
rect 110760 32160 110920 32320
rect 110760 32320 110920 32480
rect 110760 32480 110920 32640
rect 110760 32640 110920 32800
rect 110760 32800 110920 32960
rect 110760 32960 110920 33120
rect 110760 33120 110920 33280
rect 110760 33280 110920 33440
rect 110760 33440 110920 33600
rect 110760 33600 110920 33760
rect 110760 33760 110920 33920
rect 110760 33920 110920 34080
rect 110760 34080 110920 34240
rect 110760 34240 110920 34400
rect 110760 34400 110920 34560
rect 110760 34560 110920 34720
rect 110760 34720 110920 34880
rect 110760 34880 110920 35040
rect 110760 35040 110920 35200
rect 110760 35200 110920 35360
rect 110760 35360 110920 35520
rect 110760 35520 110920 35680
rect 110920 26720 111080 26880
rect 110920 26880 111080 27040
rect 110920 27040 111080 27200
rect 110920 27200 111080 27360
rect 110920 27360 111080 27520
rect 110920 27520 111080 27680
rect 110920 27680 111080 27840
rect 110920 27840 111080 28000
rect 110920 28000 111080 28160
rect 110920 28160 111080 28320
rect 110920 28320 111080 28480
rect 110920 28480 111080 28640
rect 110920 28640 111080 28800
rect 110920 28800 111080 28960
rect 110920 28960 111080 29120
rect 110920 29120 111080 29280
rect 110920 29280 111080 29440
rect 110920 31840 111080 32000
rect 110920 32000 111080 32160
rect 110920 32160 111080 32320
rect 110920 32320 111080 32480
rect 110920 32480 111080 32640
rect 110920 32640 111080 32800
rect 110920 32800 111080 32960
rect 110920 32960 111080 33120
rect 110920 33120 111080 33280
rect 110920 33280 111080 33440
rect 110920 33440 111080 33600
rect 110920 33600 111080 33760
rect 110920 33760 111080 33920
rect 110920 33920 111080 34080
rect 110920 34080 111080 34240
rect 110920 34240 111080 34400
rect 110920 34400 111080 34560
rect 110920 34560 111080 34720
rect 110920 34720 111080 34880
rect 110920 34880 111080 35040
rect 110920 35040 111080 35200
rect 110920 35200 111080 35360
rect 110920 35360 111080 35520
rect 111080 26880 111240 27040
rect 111080 27040 111240 27200
rect 111080 27200 111240 27360
rect 111080 27360 111240 27520
rect 111080 27520 111240 27680
rect 111080 27680 111240 27840
rect 111080 27840 111240 28000
rect 111080 28000 111240 28160
rect 111080 28160 111240 28320
rect 111080 28320 111240 28480
rect 111080 28480 111240 28640
rect 111080 28640 111240 28800
rect 111080 28800 111240 28960
rect 111080 28960 111240 29120
rect 111080 29120 111240 29280
rect 111080 29280 111240 29440
rect 111080 31680 111240 31840
rect 111080 31840 111240 32000
rect 111080 32000 111240 32160
rect 111080 32160 111240 32320
rect 111080 32320 111240 32480
rect 111080 32480 111240 32640
rect 111080 32640 111240 32800
rect 111080 32800 111240 32960
rect 111080 32960 111240 33120
rect 111080 33120 111240 33280
rect 111080 33280 111240 33440
rect 111080 33440 111240 33600
rect 111080 33600 111240 33760
rect 111080 33760 111240 33920
rect 111080 33920 111240 34080
rect 111080 34080 111240 34240
rect 111080 34240 111240 34400
rect 111080 34400 111240 34560
rect 111080 34560 111240 34720
rect 111080 34720 111240 34880
rect 111080 34880 111240 35040
rect 111080 35040 111240 35200
rect 111240 26880 111400 27040
rect 111240 27040 111400 27200
rect 111240 27200 111400 27360
rect 111240 27360 111400 27520
rect 111240 27520 111400 27680
rect 111240 27680 111400 27840
rect 111240 27840 111400 28000
rect 111240 28000 111400 28160
rect 111240 28160 111400 28320
rect 111240 28320 111400 28480
rect 111240 28480 111400 28640
rect 111240 28640 111400 28800
rect 111240 28800 111400 28960
rect 111240 28960 111400 29120
rect 111240 29120 111400 29280
rect 111240 29280 111400 29440
rect 111240 31680 111400 31840
rect 111240 31840 111400 32000
rect 111240 32000 111400 32160
rect 111240 32160 111400 32320
rect 111240 32320 111400 32480
rect 111240 32480 111400 32640
rect 111240 32640 111400 32800
rect 111240 32800 111400 32960
rect 111240 32960 111400 33120
rect 111240 33120 111400 33280
rect 111240 33280 111400 33440
rect 111240 33440 111400 33600
rect 111240 33600 111400 33760
rect 111240 33760 111400 33920
rect 111240 33920 111400 34080
rect 111240 34080 111400 34240
rect 111240 34240 111400 34400
rect 111240 34400 111400 34560
rect 111240 34560 111400 34720
rect 111240 34720 111400 34880
rect 111240 34880 111400 35040
rect 111240 35040 111400 35200
rect 111240 35200 111400 35360
rect 111400 26880 111560 27040
rect 111400 27040 111560 27200
rect 111400 27200 111560 27360
rect 111400 27360 111560 27520
rect 111400 27520 111560 27680
rect 111400 27680 111560 27840
rect 111400 27840 111560 28000
rect 111400 28000 111560 28160
rect 111400 28160 111560 28320
rect 111400 28320 111560 28480
rect 111400 28480 111560 28640
rect 111400 28640 111560 28800
rect 111400 28800 111560 28960
rect 111400 28960 111560 29120
rect 111400 29120 111560 29280
rect 111400 29280 111560 29440
rect 111400 31520 111560 31680
rect 111400 31680 111560 31840
rect 111400 31840 111560 32000
rect 111400 32000 111560 32160
rect 111400 32160 111560 32320
rect 111400 32320 111560 32480
rect 111400 32480 111560 32640
rect 111400 32640 111560 32800
rect 111400 32800 111560 32960
rect 111400 32960 111560 33120
rect 111400 33120 111560 33280
rect 111400 33280 111560 33440
rect 111400 33440 111560 33600
rect 111400 33600 111560 33760
rect 111400 33760 111560 33920
rect 111400 33920 111560 34080
rect 111400 34080 111560 34240
rect 111400 34240 111560 34400
rect 111400 34400 111560 34560
rect 111400 34560 111560 34720
rect 111400 34720 111560 34880
rect 111400 34880 111560 35040
rect 111400 35040 111560 35200
rect 111400 35200 111560 35360
rect 111400 35360 111560 35520
rect 111400 35520 111560 35680
rect 111560 26880 111720 27040
rect 111560 27040 111720 27200
rect 111560 27200 111720 27360
rect 111560 27360 111720 27520
rect 111560 27520 111720 27680
rect 111560 27680 111720 27840
rect 111560 27840 111720 28000
rect 111560 28000 111720 28160
rect 111560 28160 111720 28320
rect 111560 28320 111720 28480
rect 111560 28480 111720 28640
rect 111560 28640 111720 28800
rect 111560 28800 111720 28960
rect 111560 28960 111720 29120
rect 111560 29120 111720 29280
rect 111560 29280 111720 29440
rect 111560 29440 111720 29600
rect 111560 31520 111720 31680
rect 111560 31680 111720 31840
rect 111560 31840 111720 32000
rect 111560 32000 111720 32160
rect 111560 32160 111720 32320
rect 111560 32320 111720 32480
rect 111560 32480 111720 32640
rect 111560 32640 111720 32800
rect 111560 32800 111720 32960
rect 111560 32960 111720 33120
rect 111560 33120 111720 33280
rect 111560 33280 111720 33440
rect 111560 33440 111720 33600
rect 111560 33600 111720 33760
rect 111560 33760 111720 33920
rect 111560 33920 111720 34080
rect 111560 34080 111720 34240
rect 111560 34240 111720 34400
rect 111560 34400 111720 34560
rect 111560 34560 111720 34720
rect 111560 34720 111720 34880
rect 111560 34880 111720 35040
rect 111560 35040 111720 35200
rect 111560 35200 111720 35360
rect 111560 35360 111720 35520
rect 111560 35520 111720 35680
rect 111560 35680 111720 35840
rect 111560 35840 111720 36000
rect 111560 36000 111720 36160
rect 111720 26880 111880 27040
rect 111720 27040 111880 27200
rect 111720 27200 111880 27360
rect 111720 27360 111880 27520
rect 111720 27520 111880 27680
rect 111720 27680 111880 27840
rect 111720 27840 111880 28000
rect 111720 28000 111880 28160
rect 111720 28160 111880 28320
rect 111720 28320 111880 28480
rect 111720 28480 111880 28640
rect 111720 28640 111880 28800
rect 111720 28800 111880 28960
rect 111720 28960 111880 29120
rect 111720 29120 111880 29280
rect 111720 29280 111880 29440
rect 111720 29440 111880 29600
rect 111720 29600 111880 29760
rect 111720 31360 111880 31520
rect 111720 31520 111880 31680
rect 111720 31680 111880 31840
rect 111720 31840 111880 32000
rect 111720 32000 111880 32160
rect 111720 32160 111880 32320
rect 111720 32320 111880 32480
rect 111720 32480 111880 32640
rect 111720 32640 111880 32800
rect 111720 32800 111880 32960
rect 111720 32960 111880 33120
rect 111720 33120 111880 33280
rect 111720 33280 111880 33440
rect 111720 33440 111880 33600
rect 111720 33600 111880 33760
rect 111720 33760 111880 33920
rect 111720 33920 111880 34080
rect 111720 34080 111880 34240
rect 111720 34240 111880 34400
rect 111720 34400 111880 34560
rect 111720 34560 111880 34720
rect 111720 34720 111880 34880
rect 111720 34880 111880 35040
rect 111720 35040 111880 35200
rect 111720 35200 111880 35360
rect 111720 35360 111880 35520
rect 111720 35520 111880 35680
rect 111720 35680 111880 35840
rect 111720 35840 111880 36000
rect 111720 36000 111880 36160
rect 111720 36160 111880 36320
rect 111720 36320 111880 36480
rect 111720 36480 111880 36640
rect 111880 27040 112040 27200
rect 111880 27200 112040 27360
rect 111880 27360 112040 27520
rect 111880 27520 112040 27680
rect 111880 27680 112040 27840
rect 111880 27840 112040 28000
rect 111880 28000 112040 28160
rect 111880 28160 112040 28320
rect 111880 28320 112040 28480
rect 111880 28480 112040 28640
rect 111880 28640 112040 28800
rect 111880 28800 112040 28960
rect 111880 28960 112040 29120
rect 111880 29120 112040 29280
rect 111880 29280 112040 29440
rect 111880 29440 112040 29600
rect 111880 29600 112040 29760
rect 111880 29760 112040 29920
rect 111880 31200 112040 31360
rect 111880 31360 112040 31520
rect 111880 31520 112040 31680
rect 111880 31680 112040 31840
rect 111880 31840 112040 32000
rect 111880 32000 112040 32160
rect 111880 32160 112040 32320
rect 111880 32320 112040 32480
rect 111880 32480 112040 32640
rect 111880 32640 112040 32800
rect 111880 32800 112040 32960
rect 111880 32960 112040 33120
rect 111880 33120 112040 33280
rect 111880 33280 112040 33440
rect 111880 33440 112040 33600
rect 111880 33600 112040 33760
rect 111880 33760 112040 33920
rect 111880 33920 112040 34080
rect 111880 34080 112040 34240
rect 111880 34240 112040 34400
rect 111880 34400 112040 34560
rect 111880 34560 112040 34720
rect 111880 34720 112040 34880
rect 111880 34880 112040 35040
rect 111880 35040 112040 35200
rect 111880 35200 112040 35360
rect 111880 35360 112040 35520
rect 111880 35520 112040 35680
rect 111880 35680 112040 35840
rect 111880 35840 112040 36000
rect 111880 36000 112040 36160
rect 111880 36160 112040 36320
rect 111880 36320 112040 36480
rect 111880 36480 112040 36640
rect 111880 36640 112040 36800
rect 111880 36800 112040 36960
rect 111880 36960 112040 37120
rect 112040 27040 112200 27200
rect 112040 27200 112200 27360
rect 112040 27360 112200 27520
rect 112040 27520 112200 27680
rect 112040 27680 112200 27840
rect 112040 27840 112200 28000
rect 112040 28000 112200 28160
rect 112040 28160 112200 28320
rect 112040 28320 112200 28480
rect 112040 28480 112200 28640
rect 112040 28640 112200 28800
rect 112040 28800 112200 28960
rect 112040 28960 112200 29120
rect 112040 29120 112200 29280
rect 112040 29280 112200 29440
rect 112040 29440 112200 29600
rect 112040 29600 112200 29760
rect 112040 29760 112200 29920
rect 112040 29920 112200 30080
rect 112040 31040 112200 31200
rect 112040 31200 112200 31360
rect 112040 31360 112200 31520
rect 112040 31520 112200 31680
rect 112040 31680 112200 31840
rect 112040 31840 112200 32000
rect 112040 32000 112200 32160
rect 112040 32160 112200 32320
rect 112040 32320 112200 32480
rect 112040 32480 112200 32640
rect 112040 32640 112200 32800
rect 112040 32800 112200 32960
rect 112040 32960 112200 33120
rect 112040 33120 112200 33280
rect 112040 33280 112200 33440
rect 112040 33440 112200 33600
rect 112040 33600 112200 33760
rect 112040 33760 112200 33920
rect 112040 33920 112200 34080
rect 112040 34080 112200 34240
rect 112040 34240 112200 34400
rect 112040 34400 112200 34560
rect 112040 34560 112200 34720
rect 112040 34720 112200 34880
rect 112040 34880 112200 35040
rect 112040 35040 112200 35200
rect 112040 35200 112200 35360
rect 112040 35360 112200 35520
rect 112040 35520 112200 35680
rect 112040 35680 112200 35840
rect 112040 35840 112200 36000
rect 112040 36000 112200 36160
rect 112040 36160 112200 36320
rect 112040 36320 112200 36480
rect 112040 36480 112200 36640
rect 112040 36640 112200 36800
rect 112040 36800 112200 36960
rect 112040 36960 112200 37120
rect 112040 37120 112200 37280
rect 112040 37280 112200 37440
rect 112200 27040 112360 27200
rect 112200 27200 112360 27360
rect 112200 27360 112360 27520
rect 112200 27520 112360 27680
rect 112200 27680 112360 27840
rect 112200 27840 112360 28000
rect 112200 28000 112360 28160
rect 112200 28160 112360 28320
rect 112200 28320 112360 28480
rect 112200 28480 112360 28640
rect 112200 28640 112360 28800
rect 112200 28800 112360 28960
rect 112200 28960 112360 29120
rect 112200 29120 112360 29280
rect 112200 29280 112360 29440
rect 112200 29440 112360 29600
rect 112200 29600 112360 29760
rect 112200 29760 112360 29920
rect 112200 29920 112360 30080
rect 112200 30080 112360 30240
rect 112200 30240 112360 30400
rect 112200 30400 112360 30560
rect 112200 30560 112360 30720
rect 112200 30720 112360 30880
rect 112200 30880 112360 31040
rect 112200 31040 112360 31200
rect 112200 31200 112360 31360
rect 112200 31360 112360 31520
rect 112200 31520 112360 31680
rect 112200 31680 112360 31840
rect 112200 31840 112360 32000
rect 112200 32000 112360 32160
rect 112200 32160 112360 32320
rect 112200 32320 112360 32480
rect 112200 32480 112360 32640
rect 112200 32640 112360 32800
rect 112200 32800 112360 32960
rect 112200 32960 112360 33120
rect 112200 33120 112360 33280
rect 112200 33280 112360 33440
rect 112200 33440 112360 33600
rect 112200 33600 112360 33760
rect 112200 33760 112360 33920
rect 112200 33920 112360 34080
rect 112200 34080 112360 34240
rect 112200 34240 112360 34400
rect 112200 34400 112360 34560
rect 112200 34560 112360 34720
rect 112200 34720 112360 34880
rect 112200 34880 112360 35040
rect 112200 35040 112360 35200
rect 112200 35200 112360 35360
rect 112200 35360 112360 35520
rect 112200 35520 112360 35680
rect 112200 35680 112360 35840
rect 112200 35840 112360 36000
rect 112200 36000 112360 36160
rect 112200 36160 112360 36320
rect 112200 36320 112360 36480
rect 112200 36480 112360 36640
rect 112200 36640 112360 36800
rect 112200 36800 112360 36960
rect 112200 36960 112360 37120
rect 112200 37120 112360 37280
rect 112200 37280 112360 37440
rect 112200 37440 112360 37600
rect 112200 37600 112360 37760
rect 112200 37760 112360 37920
rect 112360 27200 112520 27360
rect 112360 27360 112520 27520
rect 112360 27520 112520 27680
rect 112360 27680 112520 27840
rect 112360 27840 112520 28000
rect 112360 28000 112520 28160
rect 112360 28160 112520 28320
rect 112360 28320 112520 28480
rect 112360 28480 112520 28640
rect 112360 28640 112520 28800
rect 112360 28800 112520 28960
rect 112360 28960 112520 29120
rect 112360 29120 112520 29280
rect 112360 29280 112520 29440
rect 112360 29440 112520 29600
rect 112360 29600 112520 29760
rect 112360 29760 112520 29920
rect 112360 29920 112520 30080
rect 112360 30080 112520 30240
rect 112360 30240 112520 30400
rect 112360 30400 112520 30560
rect 112360 30560 112520 30720
rect 112360 30720 112520 30880
rect 112360 30880 112520 31040
rect 112360 31040 112520 31200
rect 112360 31200 112520 31360
rect 112360 31360 112520 31520
rect 112360 31520 112520 31680
rect 112360 31680 112520 31840
rect 112360 31840 112520 32000
rect 112360 32000 112520 32160
rect 112360 32160 112520 32320
rect 112360 32320 112520 32480
rect 112360 32480 112520 32640
rect 112360 32640 112520 32800
rect 112360 32800 112520 32960
rect 112360 32960 112520 33120
rect 112360 33120 112520 33280
rect 112360 33280 112520 33440
rect 112360 33440 112520 33600
rect 112360 33600 112520 33760
rect 112360 33760 112520 33920
rect 112360 33920 112520 34080
rect 112360 34080 112520 34240
rect 112360 34240 112520 34400
rect 112360 34400 112520 34560
rect 112360 34560 112520 34720
rect 112360 34720 112520 34880
rect 112360 34880 112520 35040
rect 112360 35040 112520 35200
rect 112360 35200 112520 35360
rect 112360 35360 112520 35520
rect 112360 35520 112520 35680
rect 112360 35680 112520 35840
rect 112360 35840 112520 36000
rect 112360 36000 112520 36160
rect 112360 36160 112520 36320
rect 112360 36320 112520 36480
rect 112360 36480 112520 36640
rect 112360 36640 112520 36800
rect 112360 36800 112520 36960
rect 112360 36960 112520 37120
rect 112360 37120 112520 37280
rect 112360 37280 112520 37440
rect 112360 37440 112520 37600
rect 112360 37600 112520 37760
rect 112360 37760 112520 37920
rect 112360 37920 112520 38080
rect 112360 38080 112520 38240
rect 112360 38240 112520 38400
rect 112520 27200 112680 27360
rect 112520 27360 112680 27520
rect 112520 27520 112680 27680
rect 112520 27680 112680 27840
rect 112520 27840 112680 28000
rect 112520 28000 112680 28160
rect 112520 28160 112680 28320
rect 112520 28320 112680 28480
rect 112520 28480 112680 28640
rect 112520 28640 112680 28800
rect 112520 28800 112680 28960
rect 112520 28960 112680 29120
rect 112520 29120 112680 29280
rect 112520 29280 112680 29440
rect 112520 29440 112680 29600
rect 112520 29600 112680 29760
rect 112520 29760 112680 29920
rect 112520 29920 112680 30080
rect 112520 30080 112680 30240
rect 112520 30240 112680 30400
rect 112520 30400 112680 30560
rect 112520 30560 112680 30720
rect 112520 30720 112680 30880
rect 112520 30880 112680 31040
rect 112520 31040 112680 31200
rect 112520 31200 112680 31360
rect 112520 31360 112680 31520
rect 112520 31520 112680 31680
rect 112520 31680 112680 31840
rect 112520 31840 112680 32000
rect 112520 32000 112680 32160
rect 112520 32160 112680 32320
rect 112520 32320 112680 32480
rect 112520 32480 112680 32640
rect 112520 32640 112680 32800
rect 112520 32800 112680 32960
rect 112520 32960 112680 33120
rect 112520 33120 112680 33280
rect 112520 33280 112680 33440
rect 112520 33440 112680 33600
rect 112520 33600 112680 33760
rect 112520 33760 112680 33920
rect 112520 33920 112680 34080
rect 112520 34080 112680 34240
rect 112520 34240 112680 34400
rect 112520 34400 112680 34560
rect 112520 34560 112680 34720
rect 112520 34720 112680 34880
rect 112520 34880 112680 35040
rect 112520 35040 112680 35200
rect 112520 35200 112680 35360
rect 112520 35360 112680 35520
rect 112520 35520 112680 35680
rect 112520 35680 112680 35840
rect 112520 35840 112680 36000
rect 112520 36000 112680 36160
rect 112520 36160 112680 36320
rect 112520 36320 112680 36480
rect 112520 36480 112680 36640
rect 112520 36640 112680 36800
rect 112520 36800 112680 36960
rect 112520 36960 112680 37120
rect 112520 37120 112680 37280
rect 112520 37280 112680 37440
rect 112520 37440 112680 37600
rect 112520 37600 112680 37760
rect 112520 37760 112680 37920
rect 112520 37920 112680 38080
rect 112520 38080 112680 38240
rect 112520 38240 112680 38400
rect 112520 38400 112680 38560
rect 112520 38560 112680 38720
rect 112520 38720 112680 38880
rect 112680 27360 112840 27520
rect 112680 27520 112840 27680
rect 112680 27680 112840 27840
rect 112680 27840 112840 28000
rect 112680 28000 112840 28160
rect 112680 28160 112840 28320
rect 112680 28320 112840 28480
rect 112680 28480 112840 28640
rect 112680 28640 112840 28800
rect 112680 28800 112840 28960
rect 112680 28960 112840 29120
rect 112680 29120 112840 29280
rect 112680 29280 112840 29440
rect 112680 29440 112840 29600
rect 112680 29600 112840 29760
rect 112680 29760 112840 29920
rect 112680 29920 112840 30080
rect 112680 30080 112840 30240
rect 112680 30240 112840 30400
rect 112680 30400 112840 30560
rect 112680 30560 112840 30720
rect 112680 30720 112840 30880
rect 112680 30880 112840 31040
rect 112680 31040 112840 31200
rect 112680 31200 112840 31360
rect 112680 31360 112840 31520
rect 112680 31520 112840 31680
rect 112680 31680 112840 31840
rect 112680 31840 112840 32000
rect 112680 32000 112840 32160
rect 112680 32160 112840 32320
rect 112680 32320 112840 32480
rect 112680 32480 112840 32640
rect 112680 32640 112840 32800
rect 112680 32800 112840 32960
rect 112680 32960 112840 33120
rect 112680 33120 112840 33280
rect 112680 33280 112840 33440
rect 112680 33440 112840 33600
rect 112680 33600 112840 33760
rect 112680 33760 112840 33920
rect 112680 33920 112840 34080
rect 112680 34080 112840 34240
rect 112680 34240 112840 34400
rect 112680 34400 112840 34560
rect 112680 34560 112840 34720
rect 112680 34720 112840 34880
rect 112680 34880 112840 35040
rect 112680 35040 112840 35200
rect 112680 35200 112840 35360
rect 112680 35360 112840 35520
rect 112680 35520 112840 35680
rect 112680 35680 112840 35840
rect 112680 35840 112840 36000
rect 112680 36000 112840 36160
rect 112680 36160 112840 36320
rect 112680 36320 112840 36480
rect 112680 36480 112840 36640
rect 112680 36640 112840 36800
rect 112680 36800 112840 36960
rect 112680 36960 112840 37120
rect 112680 37120 112840 37280
rect 112680 37280 112840 37440
rect 112680 37440 112840 37600
rect 112680 37600 112840 37760
rect 112680 37760 112840 37920
rect 112680 37920 112840 38080
rect 112680 38080 112840 38240
rect 112680 38240 112840 38400
rect 112680 38400 112840 38560
rect 112680 38560 112840 38720
rect 112680 38720 112840 38880
rect 112680 38880 112840 39040
rect 112680 39040 112840 39200
rect 112840 27360 113000 27520
rect 112840 27520 113000 27680
rect 112840 27680 113000 27840
rect 112840 27840 113000 28000
rect 112840 28000 113000 28160
rect 112840 28160 113000 28320
rect 112840 28320 113000 28480
rect 112840 28480 113000 28640
rect 112840 28640 113000 28800
rect 112840 28800 113000 28960
rect 112840 28960 113000 29120
rect 112840 29120 113000 29280
rect 112840 29280 113000 29440
rect 112840 29440 113000 29600
rect 112840 29600 113000 29760
rect 112840 29760 113000 29920
rect 112840 29920 113000 30080
rect 112840 30080 113000 30240
rect 112840 30240 113000 30400
rect 112840 30400 113000 30560
rect 112840 30560 113000 30720
rect 112840 30720 113000 30880
rect 112840 30880 113000 31040
rect 112840 31040 113000 31200
rect 112840 31200 113000 31360
rect 112840 31360 113000 31520
rect 112840 31520 113000 31680
rect 112840 31680 113000 31840
rect 112840 31840 113000 32000
rect 112840 32000 113000 32160
rect 112840 32160 113000 32320
rect 112840 32320 113000 32480
rect 112840 32480 113000 32640
rect 112840 32640 113000 32800
rect 112840 32800 113000 32960
rect 112840 32960 113000 33120
rect 112840 33120 113000 33280
rect 112840 33280 113000 33440
rect 112840 33440 113000 33600
rect 112840 33600 113000 33760
rect 112840 33760 113000 33920
rect 112840 33920 113000 34080
rect 112840 34080 113000 34240
rect 112840 34240 113000 34400
rect 112840 34400 113000 34560
rect 112840 34560 113000 34720
rect 112840 34720 113000 34880
rect 112840 34880 113000 35040
rect 112840 35040 113000 35200
rect 112840 35200 113000 35360
rect 112840 35360 113000 35520
rect 112840 35520 113000 35680
rect 112840 35680 113000 35840
rect 112840 35840 113000 36000
rect 112840 36000 113000 36160
rect 112840 36160 113000 36320
rect 112840 36320 113000 36480
rect 112840 36480 113000 36640
rect 112840 36640 113000 36800
rect 112840 36800 113000 36960
rect 112840 36960 113000 37120
rect 112840 37120 113000 37280
rect 112840 37280 113000 37440
rect 112840 37440 113000 37600
rect 112840 37600 113000 37760
rect 112840 37760 113000 37920
rect 112840 37920 113000 38080
rect 112840 38080 113000 38240
rect 112840 38240 113000 38400
rect 112840 38400 113000 38560
rect 112840 38560 113000 38720
rect 112840 38720 113000 38880
rect 112840 38880 113000 39040
rect 112840 39040 113000 39200
rect 112840 39200 113000 39360
rect 112840 39360 113000 39520
rect 112840 39520 113000 39680
rect 113000 27520 113160 27680
rect 113000 27680 113160 27840
rect 113000 27840 113160 28000
rect 113000 28000 113160 28160
rect 113000 28160 113160 28320
rect 113000 28320 113160 28480
rect 113000 28480 113160 28640
rect 113000 28640 113160 28800
rect 113000 28800 113160 28960
rect 113000 28960 113160 29120
rect 113000 29120 113160 29280
rect 113000 29280 113160 29440
rect 113000 29440 113160 29600
rect 113000 29600 113160 29760
rect 113000 29760 113160 29920
rect 113000 29920 113160 30080
rect 113000 30080 113160 30240
rect 113000 30240 113160 30400
rect 113000 30400 113160 30560
rect 113000 30560 113160 30720
rect 113000 30720 113160 30880
rect 113000 30880 113160 31040
rect 113000 31040 113160 31200
rect 113000 31200 113160 31360
rect 113000 31360 113160 31520
rect 113000 31520 113160 31680
rect 113000 31680 113160 31840
rect 113000 31840 113160 32000
rect 113000 32000 113160 32160
rect 113000 32160 113160 32320
rect 113000 32320 113160 32480
rect 113000 32480 113160 32640
rect 113000 32640 113160 32800
rect 113000 32800 113160 32960
rect 113000 32960 113160 33120
rect 113000 33120 113160 33280
rect 113000 33280 113160 33440
rect 113000 33440 113160 33600
rect 113000 33600 113160 33760
rect 113000 33760 113160 33920
rect 113000 33920 113160 34080
rect 113000 34080 113160 34240
rect 113000 34240 113160 34400
rect 113000 34400 113160 34560
rect 113000 34560 113160 34720
rect 113000 34720 113160 34880
rect 113000 34880 113160 35040
rect 113000 35040 113160 35200
rect 113000 35200 113160 35360
rect 113000 35360 113160 35520
rect 113000 35520 113160 35680
rect 113000 35680 113160 35840
rect 113000 35840 113160 36000
rect 113000 36000 113160 36160
rect 113000 36160 113160 36320
rect 113000 36320 113160 36480
rect 113000 36480 113160 36640
rect 113000 36640 113160 36800
rect 113000 36800 113160 36960
rect 113000 36960 113160 37120
rect 113000 37120 113160 37280
rect 113000 37280 113160 37440
rect 113000 37440 113160 37600
rect 113000 37600 113160 37760
rect 113000 37760 113160 37920
rect 113000 37920 113160 38080
rect 113000 38080 113160 38240
rect 113000 38240 113160 38400
rect 113000 38400 113160 38560
rect 113000 38560 113160 38720
rect 113000 38720 113160 38880
rect 113000 38880 113160 39040
rect 113000 39040 113160 39200
rect 113000 39200 113160 39360
rect 113000 39360 113160 39520
rect 113000 39520 113160 39680
rect 113000 39680 113160 39840
rect 113000 39840 113160 40000
rect 113000 40000 113160 40160
rect 113160 27520 113320 27680
rect 113160 27680 113320 27840
rect 113160 27840 113320 28000
rect 113160 28000 113320 28160
rect 113160 28160 113320 28320
rect 113160 28320 113320 28480
rect 113160 28480 113320 28640
rect 113160 28640 113320 28800
rect 113160 28800 113320 28960
rect 113160 28960 113320 29120
rect 113160 29120 113320 29280
rect 113160 29280 113320 29440
rect 113160 29440 113320 29600
rect 113160 29600 113320 29760
rect 113160 29760 113320 29920
rect 113160 29920 113320 30080
rect 113160 30080 113320 30240
rect 113160 30240 113320 30400
rect 113160 30400 113320 30560
rect 113160 30560 113320 30720
rect 113160 30720 113320 30880
rect 113160 30880 113320 31040
rect 113160 31040 113320 31200
rect 113160 31200 113320 31360
rect 113160 31360 113320 31520
rect 113160 31520 113320 31680
rect 113160 31680 113320 31840
rect 113160 31840 113320 32000
rect 113160 32000 113320 32160
rect 113160 32160 113320 32320
rect 113160 32320 113320 32480
rect 113160 32480 113320 32640
rect 113160 32640 113320 32800
rect 113160 32800 113320 32960
rect 113160 32960 113320 33120
rect 113160 33120 113320 33280
rect 113160 33280 113320 33440
rect 113160 33440 113320 33600
rect 113160 33600 113320 33760
rect 113160 33760 113320 33920
rect 113160 33920 113320 34080
rect 113160 34080 113320 34240
rect 113160 34240 113320 34400
rect 113160 34400 113320 34560
rect 113160 34560 113320 34720
rect 113160 34720 113320 34880
rect 113160 34880 113320 35040
rect 113160 35040 113320 35200
rect 113160 35200 113320 35360
rect 113160 35360 113320 35520
rect 113160 35520 113320 35680
rect 113160 35680 113320 35840
rect 113160 35840 113320 36000
rect 113160 36000 113320 36160
rect 113160 36160 113320 36320
rect 113160 36320 113320 36480
rect 113160 36480 113320 36640
rect 113160 36640 113320 36800
rect 113160 36800 113320 36960
rect 113160 36960 113320 37120
rect 113160 37120 113320 37280
rect 113160 37280 113320 37440
rect 113160 37440 113320 37600
rect 113160 37600 113320 37760
rect 113160 37760 113320 37920
rect 113160 37920 113320 38080
rect 113160 38080 113320 38240
rect 113160 38240 113320 38400
rect 113160 38400 113320 38560
rect 113160 38560 113320 38720
rect 113160 38720 113320 38880
rect 113160 38880 113320 39040
rect 113160 39040 113320 39200
rect 113160 39200 113320 39360
rect 113160 39360 113320 39520
rect 113160 39520 113320 39680
rect 113160 39680 113320 39840
rect 113160 39840 113320 40000
rect 113160 40000 113320 40160
rect 113160 40160 113320 40320
rect 113160 40320 113320 40480
rect 113160 40480 113320 40640
rect 113320 27680 113480 27840
rect 113320 27840 113480 28000
rect 113320 28000 113480 28160
rect 113320 28160 113480 28320
rect 113320 28320 113480 28480
rect 113320 28480 113480 28640
rect 113320 28640 113480 28800
rect 113320 28800 113480 28960
rect 113320 28960 113480 29120
rect 113320 29120 113480 29280
rect 113320 29280 113480 29440
rect 113320 29440 113480 29600
rect 113320 29600 113480 29760
rect 113320 29760 113480 29920
rect 113320 29920 113480 30080
rect 113320 30080 113480 30240
rect 113320 30240 113480 30400
rect 113320 30400 113480 30560
rect 113320 30560 113480 30720
rect 113320 30720 113480 30880
rect 113320 30880 113480 31040
rect 113320 31040 113480 31200
rect 113320 31200 113480 31360
rect 113320 31360 113480 31520
rect 113320 31520 113480 31680
rect 113320 31680 113480 31840
rect 113320 31840 113480 32000
rect 113320 32000 113480 32160
rect 113320 32160 113480 32320
rect 113320 32320 113480 32480
rect 113320 32480 113480 32640
rect 113320 32640 113480 32800
rect 113320 32800 113480 32960
rect 113320 32960 113480 33120
rect 113320 33120 113480 33280
rect 113320 33280 113480 33440
rect 113320 33440 113480 33600
rect 113320 33600 113480 33760
rect 113320 33760 113480 33920
rect 113320 33920 113480 34080
rect 113320 34080 113480 34240
rect 113320 34240 113480 34400
rect 113320 34400 113480 34560
rect 113320 34560 113480 34720
rect 113320 34720 113480 34880
rect 113320 34880 113480 35040
rect 113320 35040 113480 35200
rect 113320 35200 113480 35360
rect 113320 35360 113480 35520
rect 113320 35520 113480 35680
rect 113320 35680 113480 35840
rect 113320 35840 113480 36000
rect 113320 36000 113480 36160
rect 113320 36160 113480 36320
rect 113320 36320 113480 36480
rect 113320 36480 113480 36640
rect 113320 36640 113480 36800
rect 113320 36800 113480 36960
rect 113320 36960 113480 37120
rect 113320 37120 113480 37280
rect 113320 37280 113480 37440
rect 113320 37440 113480 37600
rect 113320 37600 113480 37760
rect 113320 37760 113480 37920
rect 113320 37920 113480 38080
rect 113320 38080 113480 38240
rect 113320 38240 113480 38400
rect 113320 38400 113480 38560
rect 113320 38560 113480 38720
rect 113320 38720 113480 38880
rect 113320 38880 113480 39040
rect 113320 39040 113480 39200
rect 113320 39200 113480 39360
rect 113320 39360 113480 39520
rect 113320 39520 113480 39680
rect 113320 39680 113480 39840
rect 113320 39840 113480 40000
rect 113320 40000 113480 40160
rect 113320 40160 113480 40320
rect 113320 40320 113480 40480
rect 113320 40480 113480 40640
rect 113320 40640 113480 40800
rect 113320 40800 113480 40960
rect 113320 40960 113480 41120
rect 113480 27840 113640 28000
rect 113480 28000 113640 28160
rect 113480 28160 113640 28320
rect 113480 28320 113640 28480
rect 113480 28480 113640 28640
rect 113480 28640 113640 28800
rect 113480 28800 113640 28960
rect 113480 28960 113640 29120
rect 113480 29120 113640 29280
rect 113480 29280 113640 29440
rect 113480 29440 113640 29600
rect 113480 29600 113640 29760
rect 113480 29760 113640 29920
rect 113480 29920 113640 30080
rect 113480 30080 113640 30240
rect 113480 30240 113640 30400
rect 113480 30400 113640 30560
rect 113480 30560 113640 30720
rect 113480 30720 113640 30880
rect 113480 30880 113640 31040
rect 113480 31040 113640 31200
rect 113480 31200 113640 31360
rect 113480 31360 113640 31520
rect 113480 31520 113640 31680
rect 113480 31680 113640 31840
rect 113480 31840 113640 32000
rect 113480 32000 113640 32160
rect 113480 32160 113640 32320
rect 113480 32320 113640 32480
rect 113480 32480 113640 32640
rect 113480 32640 113640 32800
rect 113480 32800 113640 32960
rect 113480 32960 113640 33120
rect 113480 33120 113640 33280
rect 113480 33280 113640 33440
rect 113480 33440 113640 33600
rect 113480 33600 113640 33760
rect 113480 33760 113640 33920
rect 113480 33920 113640 34080
rect 113480 34080 113640 34240
rect 113480 34240 113640 34400
rect 113480 34400 113640 34560
rect 113480 34560 113640 34720
rect 113480 34720 113640 34880
rect 113480 34880 113640 35040
rect 113480 35040 113640 35200
rect 113480 35200 113640 35360
rect 113480 35360 113640 35520
rect 113480 35520 113640 35680
rect 113480 35680 113640 35840
rect 113480 35840 113640 36000
rect 113480 36000 113640 36160
rect 113480 36160 113640 36320
rect 113480 36320 113640 36480
rect 113480 36480 113640 36640
rect 113480 36640 113640 36800
rect 113480 36800 113640 36960
rect 113480 36960 113640 37120
rect 113480 37120 113640 37280
rect 113480 37280 113640 37440
rect 113480 37440 113640 37600
rect 113480 37600 113640 37760
rect 113480 37760 113640 37920
rect 113480 37920 113640 38080
rect 113480 38080 113640 38240
rect 113480 38240 113640 38400
rect 113480 38400 113640 38560
rect 113480 38560 113640 38720
rect 113480 38720 113640 38880
rect 113480 38880 113640 39040
rect 113480 39040 113640 39200
rect 113480 39200 113640 39360
rect 113480 39360 113640 39520
rect 113480 39520 113640 39680
rect 113480 39680 113640 39840
rect 113480 39840 113640 40000
rect 113480 40000 113640 40160
rect 113480 40160 113640 40320
rect 113480 40320 113640 40480
rect 113480 40480 113640 40640
rect 113480 40640 113640 40800
rect 113480 40800 113640 40960
rect 113480 40960 113640 41120
rect 113480 41120 113640 41280
rect 113480 41280 113640 41440
rect 113480 41440 113640 41600
rect 113640 28000 113800 28160
rect 113640 28160 113800 28320
rect 113640 28320 113800 28480
rect 113640 28480 113800 28640
rect 113640 28640 113800 28800
rect 113640 28800 113800 28960
rect 113640 28960 113800 29120
rect 113640 29120 113800 29280
rect 113640 29280 113800 29440
rect 113640 29440 113800 29600
rect 113640 29600 113800 29760
rect 113640 29760 113800 29920
rect 113640 29920 113800 30080
rect 113640 30080 113800 30240
rect 113640 30240 113800 30400
rect 113640 30400 113800 30560
rect 113640 30560 113800 30720
rect 113640 30720 113800 30880
rect 113640 30880 113800 31040
rect 113640 31040 113800 31200
rect 113640 31200 113800 31360
rect 113640 31360 113800 31520
rect 113640 31520 113800 31680
rect 113640 31680 113800 31840
rect 113640 31840 113800 32000
rect 113640 32000 113800 32160
rect 113640 32160 113800 32320
rect 113640 32320 113800 32480
rect 113640 32480 113800 32640
rect 113640 32640 113800 32800
rect 113640 32800 113800 32960
rect 113640 32960 113800 33120
rect 113640 33120 113800 33280
rect 113640 33280 113800 33440
rect 113640 33920 113800 34080
rect 113640 34080 113800 34240
rect 113640 34240 113800 34400
rect 113640 34400 113800 34560
rect 113640 34560 113800 34720
rect 113640 34720 113800 34880
rect 113640 34880 113800 35040
rect 113640 35040 113800 35200
rect 113640 35200 113800 35360
rect 113640 35360 113800 35520
rect 113640 35520 113800 35680
rect 113640 35680 113800 35840
rect 113640 35840 113800 36000
rect 113640 36000 113800 36160
rect 113640 36160 113800 36320
rect 113640 36320 113800 36480
rect 113640 36480 113800 36640
rect 113640 36640 113800 36800
rect 113640 36800 113800 36960
rect 113640 36960 113800 37120
rect 113640 37120 113800 37280
rect 113640 37280 113800 37440
rect 113640 37440 113800 37600
rect 113640 37600 113800 37760
rect 113640 37760 113800 37920
rect 113640 37920 113800 38080
rect 113640 38080 113800 38240
rect 113640 38240 113800 38400
rect 113640 38400 113800 38560
rect 113640 38560 113800 38720
rect 113640 38720 113800 38880
rect 113640 38880 113800 39040
rect 113640 39040 113800 39200
rect 113640 39200 113800 39360
rect 113640 39360 113800 39520
rect 113640 39520 113800 39680
rect 113640 39680 113800 39840
rect 113640 39840 113800 40000
rect 113640 40000 113800 40160
rect 113640 40160 113800 40320
rect 113640 40320 113800 40480
rect 113640 40480 113800 40640
rect 113640 40640 113800 40800
rect 113640 40800 113800 40960
rect 113640 40960 113800 41120
rect 113640 41120 113800 41280
rect 113640 41280 113800 41440
rect 113640 41440 113800 41600
rect 113640 41600 113800 41760
rect 113640 41760 113800 41920
rect 113640 41920 113800 42080
rect 113800 28160 113960 28320
rect 113800 28320 113960 28480
rect 113800 28480 113960 28640
rect 113800 28640 113960 28800
rect 113800 28800 113960 28960
rect 113800 28960 113960 29120
rect 113800 29120 113960 29280
rect 113800 29280 113960 29440
rect 113800 29440 113960 29600
rect 113800 29600 113960 29760
rect 113800 29760 113960 29920
rect 113800 29920 113960 30080
rect 113800 30080 113960 30240
rect 113800 30240 113960 30400
rect 113800 30400 113960 30560
rect 113800 30560 113960 30720
rect 113800 30720 113960 30880
rect 113800 30880 113960 31040
rect 113800 31040 113960 31200
rect 113800 31200 113960 31360
rect 113800 31360 113960 31520
rect 113800 31520 113960 31680
rect 113800 31680 113960 31840
rect 113800 31840 113960 32000
rect 113800 32000 113960 32160
rect 113800 32160 113960 32320
rect 113800 32320 113960 32480
rect 113800 32480 113960 32640
rect 113800 32640 113960 32800
rect 113800 32800 113960 32960
rect 113800 32960 113960 33120
rect 113800 33120 113960 33280
rect 113800 34400 113960 34560
rect 113800 34560 113960 34720
rect 113800 34720 113960 34880
rect 113800 34880 113960 35040
rect 113800 35040 113960 35200
rect 113800 35200 113960 35360
rect 113800 35360 113960 35520
rect 113800 35520 113960 35680
rect 113800 35680 113960 35840
rect 113800 35840 113960 36000
rect 113800 36000 113960 36160
rect 113800 36160 113960 36320
rect 113800 36320 113960 36480
rect 113800 36480 113960 36640
rect 113800 36640 113960 36800
rect 113800 36800 113960 36960
rect 113800 36960 113960 37120
rect 113800 37120 113960 37280
rect 113800 37280 113960 37440
rect 113800 37440 113960 37600
rect 113800 37600 113960 37760
rect 113800 37760 113960 37920
rect 113800 37920 113960 38080
rect 113800 38080 113960 38240
rect 113800 38240 113960 38400
rect 113800 38400 113960 38560
rect 113800 38560 113960 38720
rect 113800 38720 113960 38880
rect 113800 38880 113960 39040
rect 113800 39040 113960 39200
rect 113800 39200 113960 39360
rect 113800 39360 113960 39520
rect 113800 39520 113960 39680
rect 113800 39680 113960 39840
rect 113800 39840 113960 40000
rect 113800 40000 113960 40160
rect 113800 40160 113960 40320
rect 113800 40320 113960 40480
rect 113800 40480 113960 40640
rect 113800 40640 113960 40800
rect 113800 40800 113960 40960
rect 113800 40960 113960 41120
rect 113800 41120 113960 41280
rect 113800 41280 113960 41440
rect 113800 41440 113960 41600
rect 113800 41600 113960 41760
rect 113800 41760 113960 41920
rect 113800 41920 113960 42080
rect 113800 42080 113960 42240
rect 113800 42240 113960 42400
rect 113960 28320 114120 28480
rect 113960 28480 114120 28640
rect 113960 28640 114120 28800
rect 113960 28800 114120 28960
rect 113960 28960 114120 29120
rect 113960 29120 114120 29280
rect 113960 29280 114120 29440
rect 113960 29440 114120 29600
rect 113960 29600 114120 29760
rect 113960 29760 114120 29920
rect 113960 29920 114120 30080
rect 113960 30080 114120 30240
rect 113960 30240 114120 30400
rect 113960 30400 114120 30560
rect 113960 30560 114120 30720
rect 113960 30720 114120 30880
rect 113960 30880 114120 31040
rect 113960 31040 114120 31200
rect 113960 31200 114120 31360
rect 113960 31360 114120 31520
rect 113960 31520 114120 31680
rect 113960 31680 114120 31840
rect 113960 31840 114120 32000
rect 113960 32000 114120 32160
rect 113960 32160 114120 32320
rect 113960 32320 114120 32480
rect 113960 32480 114120 32640
rect 113960 32640 114120 32800
rect 113960 32800 114120 32960
rect 113960 32960 114120 33120
rect 113960 34880 114120 35040
rect 113960 35040 114120 35200
rect 113960 35200 114120 35360
rect 113960 35360 114120 35520
rect 113960 35520 114120 35680
rect 113960 35680 114120 35840
rect 113960 35840 114120 36000
rect 113960 36000 114120 36160
rect 113960 36160 114120 36320
rect 113960 36320 114120 36480
rect 113960 36480 114120 36640
rect 113960 36640 114120 36800
rect 113960 36800 114120 36960
rect 113960 36960 114120 37120
rect 113960 37120 114120 37280
rect 113960 37280 114120 37440
rect 113960 37440 114120 37600
rect 113960 37600 114120 37760
rect 113960 37760 114120 37920
rect 113960 37920 114120 38080
rect 113960 38080 114120 38240
rect 113960 38240 114120 38400
rect 113960 38400 114120 38560
rect 113960 38560 114120 38720
rect 113960 38720 114120 38880
rect 113960 38880 114120 39040
rect 113960 39040 114120 39200
rect 113960 39200 114120 39360
rect 113960 39360 114120 39520
rect 113960 39520 114120 39680
rect 113960 39680 114120 39840
rect 113960 39840 114120 40000
rect 113960 40000 114120 40160
rect 113960 40160 114120 40320
rect 113960 40320 114120 40480
rect 113960 40480 114120 40640
rect 113960 40640 114120 40800
rect 113960 40800 114120 40960
rect 113960 40960 114120 41120
rect 113960 41120 114120 41280
rect 113960 41280 114120 41440
rect 113960 41440 114120 41600
rect 113960 41600 114120 41760
rect 113960 41760 114120 41920
rect 113960 41920 114120 42080
rect 113960 42080 114120 42240
rect 113960 42240 114120 42400
rect 113960 42400 114120 42560
rect 113960 42560 114120 42720
rect 113960 42720 114120 42880
rect 114120 28480 114280 28640
rect 114120 28640 114280 28800
rect 114120 28800 114280 28960
rect 114120 28960 114280 29120
rect 114120 29120 114280 29280
rect 114120 29280 114280 29440
rect 114120 29440 114280 29600
rect 114120 29600 114280 29760
rect 114120 29760 114280 29920
rect 114120 29920 114280 30080
rect 114120 30080 114280 30240
rect 114120 30240 114280 30400
rect 114120 30400 114280 30560
rect 114120 30560 114280 30720
rect 114120 30720 114280 30880
rect 114120 30880 114280 31040
rect 114120 31040 114280 31200
rect 114120 31200 114280 31360
rect 114120 31360 114280 31520
rect 114120 31520 114280 31680
rect 114120 31680 114280 31840
rect 114120 31840 114280 32000
rect 114120 32000 114280 32160
rect 114120 32160 114280 32320
rect 114120 32320 114280 32480
rect 114120 32480 114280 32640
rect 114120 32640 114280 32800
rect 114120 35360 114280 35520
rect 114120 35520 114280 35680
rect 114120 35680 114280 35840
rect 114120 35840 114280 36000
rect 114120 36000 114280 36160
rect 114120 36160 114280 36320
rect 114120 36320 114280 36480
rect 114120 36480 114280 36640
rect 114120 36640 114280 36800
rect 114120 36800 114280 36960
rect 114120 36960 114280 37120
rect 114120 37120 114280 37280
rect 114120 37280 114280 37440
rect 114120 37440 114280 37600
rect 114120 37600 114280 37760
rect 114120 37760 114280 37920
rect 114120 37920 114280 38080
rect 114120 38080 114280 38240
rect 114120 38240 114280 38400
rect 114120 38400 114280 38560
rect 114120 38560 114280 38720
rect 114120 38720 114280 38880
rect 114120 38880 114280 39040
rect 114120 39040 114280 39200
rect 114120 39200 114280 39360
rect 114120 39360 114280 39520
rect 114120 39520 114280 39680
rect 114120 39680 114280 39840
rect 114120 39840 114280 40000
rect 114120 40000 114280 40160
rect 114120 40160 114280 40320
rect 114120 40320 114280 40480
rect 114120 40480 114280 40640
rect 114120 40640 114280 40800
rect 114120 40800 114280 40960
rect 114120 40960 114280 41120
rect 114120 41120 114280 41280
rect 114120 41280 114280 41440
rect 114120 41440 114280 41600
rect 114120 41600 114280 41760
rect 114120 41760 114280 41920
rect 114120 41920 114280 42080
rect 114120 42080 114280 42240
rect 114120 42240 114280 42400
rect 114120 42400 114280 42560
rect 114120 42560 114280 42720
rect 114120 42720 114280 42880
rect 114120 42880 114280 43040
rect 114120 43040 114280 43200
rect 114120 43200 114280 43360
rect 114280 28800 114440 28960
rect 114280 28960 114440 29120
rect 114280 29120 114440 29280
rect 114280 29280 114440 29440
rect 114280 29440 114440 29600
rect 114280 29600 114440 29760
rect 114280 29760 114440 29920
rect 114280 29920 114440 30080
rect 114280 30080 114440 30240
rect 114280 30240 114440 30400
rect 114280 30400 114440 30560
rect 114280 30560 114440 30720
rect 114280 30720 114440 30880
rect 114280 30880 114440 31040
rect 114280 31040 114440 31200
rect 114280 31200 114440 31360
rect 114280 31360 114440 31520
rect 114280 31520 114440 31680
rect 114280 31680 114440 31840
rect 114280 31840 114440 32000
rect 114280 32000 114440 32160
rect 114280 32160 114440 32320
rect 114280 32320 114440 32480
rect 114280 32480 114440 32640
rect 114280 35840 114440 36000
rect 114280 36000 114440 36160
rect 114280 36160 114440 36320
rect 114280 36320 114440 36480
rect 114280 36480 114440 36640
rect 114280 36640 114440 36800
rect 114280 36800 114440 36960
rect 114280 36960 114440 37120
rect 114280 37120 114440 37280
rect 114280 37280 114440 37440
rect 114280 37440 114440 37600
rect 114280 37600 114440 37760
rect 114280 37760 114440 37920
rect 114280 37920 114440 38080
rect 114280 38080 114440 38240
rect 114280 38240 114440 38400
rect 114280 38400 114440 38560
rect 114280 38560 114440 38720
rect 114280 38720 114440 38880
rect 114280 38880 114440 39040
rect 114280 39040 114440 39200
rect 114280 39200 114440 39360
rect 114280 39360 114440 39520
rect 114280 39520 114440 39680
rect 114280 39680 114440 39840
rect 114280 39840 114440 40000
rect 114280 40000 114440 40160
rect 114280 40160 114440 40320
rect 114280 40320 114440 40480
rect 114280 40480 114440 40640
rect 114280 40640 114440 40800
rect 114280 40800 114440 40960
rect 114280 40960 114440 41120
rect 114280 41120 114440 41280
rect 114280 41280 114440 41440
rect 114280 41440 114440 41600
rect 114280 41600 114440 41760
rect 114280 41760 114440 41920
rect 114280 41920 114440 42080
rect 114280 42080 114440 42240
rect 114280 42240 114440 42400
rect 114280 42400 114440 42560
rect 114280 42560 114440 42720
rect 114280 42720 114440 42880
rect 114280 42880 114440 43040
rect 114280 43040 114440 43200
rect 114280 43200 114440 43360
rect 114280 43360 114440 43520
rect 114280 43520 114440 43680
rect 114280 43680 114440 43840
rect 114440 29120 114600 29280
rect 114440 29280 114600 29440
rect 114440 29440 114600 29600
rect 114440 29600 114600 29760
rect 114440 29760 114600 29920
rect 114440 29920 114600 30080
rect 114440 30080 114600 30240
rect 114440 30240 114600 30400
rect 114440 30400 114600 30560
rect 114440 30560 114600 30720
rect 114440 30720 114600 30880
rect 114440 30880 114600 31040
rect 114440 31040 114600 31200
rect 114440 31200 114600 31360
rect 114440 31360 114600 31520
rect 114440 31520 114600 31680
rect 114440 31680 114600 31840
rect 114440 31840 114600 32000
rect 114440 32000 114600 32160
rect 114440 32160 114600 32320
rect 114440 36160 114600 36320
rect 114440 36320 114600 36480
rect 114440 36480 114600 36640
rect 114440 36640 114600 36800
rect 114440 36800 114600 36960
rect 114440 36960 114600 37120
rect 114440 37120 114600 37280
rect 114440 37280 114600 37440
rect 114440 37440 114600 37600
rect 114440 37600 114600 37760
rect 114440 37760 114600 37920
rect 114440 37920 114600 38080
rect 114440 38080 114600 38240
rect 114440 38240 114600 38400
rect 114440 38400 114600 38560
rect 114440 38560 114600 38720
rect 114440 38720 114600 38880
rect 114440 38880 114600 39040
rect 114440 39040 114600 39200
rect 114440 39200 114600 39360
rect 114440 39360 114600 39520
rect 114440 39520 114600 39680
rect 114440 39680 114600 39840
rect 114440 39840 114600 40000
rect 114440 40000 114600 40160
rect 114440 40160 114600 40320
rect 114440 40320 114600 40480
rect 114440 40480 114600 40640
rect 114440 40640 114600 40800
rect 114440 40800 114600 40960
rect 114440 40960 114600 41120
rect 114440 41120 114600 41280
rect 114440 41280 114600 41440
rect 114440 41440 114600 41600
rect 114440 41600 114600 41760
rect 114440 41760 114600 41920
rect 114440 41920 114600 42080
rect 114440 42080 114600 42240
rect 114440 42240 114600 42400
rect 114440 42400 114600 42560
rect 114440 42560 114600 42720
rect 114440 42720 114600 42880
rect 114440 42880 114600 43040
rect 114440 43040 114600 43200
rect 114440 43200 114600 43360
rect 114440 43360 114600 43520
rect 114440 43520 114600 43680
rect 114440 43680 114600 43840
rect 114440 43840 114600 44000
rect 114440 44000 114600 44160
rect 114440 44160 114600 44320
rect 114600 29600 114760 29760
rect 114600 29760 114760 29920
rect 114600 29920 114760 30080
rect 114600 30080 114760 30240
rect 114600 30240 114760 30400
rect 114600 30400 114760 30560
rect 114600 30560 114760 30720
rect 114600 30720 114760 30880
rect 114600 30880 114760 31040
rect 114600 31040 114760 31200
rect 114600 31200 114760 31360
rect 114600 31360 114760 31520
rect 114600 31520 114760 31680
rect 114600 31680 114760 31840
rect 114600 36640 114760 36800
rect 114600 36800 114760 36960
rect 114600 36960 114760 37120
rect 114600 37120 114760 37280
rect 114600 37280 114760 37440
rect 114600 37440 114760 37600
rect 114600 37600 114760 37760
rect 114600 37760 114760 37920
rect 114600 37920 114760 38080
rect 114600 38080 114760 38240
rect 114600 38240 114760 38400
rect 114600 38400 114760 38560
rect 114600 38560 114760 38720
rect 114600 38720 114760 38880
rect 114600 38880 114760 39040
rect 114600 39040 114760 39200
rect 114600 39200 114760 39360
rect 114600 39360 114760 39520
rect 114600 39520 114760 39680
rect 114600 39680 114760 39840
rect 114600 39840 114760 40000
rect 114600 40000 114760 40160
rect 114600 40160 114760 40320
rect 114600 40320 114760 40480
rect 114600 40480 114760 40640
rect 114600 40640 114760 40800
rect 114600 40800 114760 40960
rect 114600 40960 114760 41120
rect 114600 41120 114760 41280
rect 114600 41280 114760 41440
rect 114600 41440 114760 41600
rect 114600 41600 114760 41760
rect 114600 41760 114760 41920
rect 114600 41920 114760 42080
rect 114600 42080 114760 42240
rect 114600 42240 114760 42400
rect 114600 42400 114760 42560
rect 114600 42560 114760 42720
rect 114600 42720 114760 42880
rect 114600 42880 114760 43040
rect 114600 43040 114760 43200
rect 114600 43200 114760 43360
rect 114600 43360 114760 43520
rect 114600 43520 114760 43680
rect 114600 43680 114760 43840
rect 114600 43840 114760 44000
rect 114600 44000 114760 44160
rect 114600 44160 114760 44320
rect 114600 44320 114760 44480
rect 114600 44480 114760 44640
rect 114600 44640 114760 44800
rect 114600 50400 114760 50560
rect 114600 50560 114760 50720
rect 114600 50720 114760 50880
rect 114600 50880 114760 51040
rect 114600 51040 114760 51200
rect 114600 51200 114760 51360
rect 114600 51360 114760 51520
rect 114600 51520 114760 51680
rect 114600 51680 114760 51840
rect 114600 51840 114760 52000
rect 114600 52000 114760 52160
rect 114600 52160 114760 52320
rect 114760 30400 114920 30560
rect 114760 30560 114920 30720
rect 114760 30720 114920 30880
rect 114760 30880 114920 31040
rect 114760 31040 114920 31200
rect 114760 31200 114920 31360
rect 114760 37120 114920 37280
rect 114760 37280 114920 37440
rect 114760 37440 114920 37600
rect 114760 37600 114920 37760
rect 114760 37760 114920 37920
rect 114760 37920 114920 38080
rect 114760 38080 114920 38240
rect 114760 38240 114920 38400
rect 114760 38400 114920 38560
rect 114760 38560 114920 38720
rect 114760 38720 114920 38880
rect 114760 38880 114920 39040
rect 114760 39040 114920 39200
rect 114760 39200 114920 39360
rect 114760 39360 114920 39520
rect 114760 39520 114920 39680
rect 114760 39680 114920 39840
rect 114760 39840 114920 40000
rect 114760 40000 114920 40160
rect 114760 40160 114920 40320
rect 114760 40320 114920 40480
rect 114760 40480 114920 40640
rect 114760 40640 114920 40800
rect 114760 40800 114920 40960
rect 114760 40960 114920 41120
rect 114760 41120 114920 41280
rect 114760 41280 114920 41440
rect 114760 41440 114920 41600
rect 114760 41600 114920 41760
rect 114760 41760 114920 41920
rect 114760 41920 114920 42080
rect 114760 42080 114920 42240
rect 114760 42240 114920 42400
rect 114760 42400 114920 42560
rect 114760 42560 114920 42720
rect 114760 42720 114920 42880
rect 114760 42880 114920 43040
rect 114760 43040 114920 43200
rect 114760 43200 114920 43360
rect 114760 43360 114920 43520
rect 114760 43520 114920 43680
rect 114760 43680 114920 43840
rect 114760 43840 114920 44000
rect 114760 44000 114920 44160
rect 114760 44160 114920 44320
rect 114760 44320 114920 44480
rect 114760 44480 114920 44640
rect 114760 44640 114920 44800
rect 114760 44800 114920 44960
rect 114760 44960 114920 45120
rect 114760 45120 114920 45280
rect 114760 45280 114920 45440
rect 114760 49920 114920 50080
rect 114760 50080 114920 50240
rect 114760 50240 114920 50400
rect 114760 50400 114920 50560
rect 114760 50560 114920 50720
rect 114760 50720 114920 50880
rect 114760 50880 114920 51040
rect 114760 51040 114920 51200
rect 114760 51200 114920 51360
rect 114760 51360 114920 51520
rect 114760 51520 114920 51680
rect 114760 51680 114920 51840
rect 114760 51840 114920 52000
rect 114760 52000 114920 52160
rect 114760 52160 114920 52320
rect 114760 52320 114920 52480
rect 114760 52480 114920 52640
rect 114760 52640 114920 52800
rect 114920 37600 115080 37760
rect 114920 37760 115080 37920
rect 114920 37920 115080 38080
rect 114920 38080 115080 38240
rect 114920 38240 115080 38400
rect 114920 38400 115080 38560
rect 114920 38560 115080 38720
rect 114920 38720 115080 38880
rect 114920 38880 115080 39040
rect 114920 39040 115080 39200
rect 114920 39200 115080 39360
rect 114920 39360 115080 39520
rect 114920 39520 115080 39680
rect 114920 39680 115080 39840
rect 114920 39840 115080 40000
rect 114920 40000 115080 40160
rect 114920 40160 115080 40320
rect 114920 40320 115080 40480
rect 114920 40480 115080 40640
rect 114920 40640 115080 40800
rect 114920 40800 115080 40960
rect 114920 40960 115080 41120
rect 114920 41120 115080 41280
rect 114920 41280 115080 41440
rect 114920 41440 115080 41600
rect 114920 41600 115080 41760
rect 114920 41760 115080 41920
rect 114920 41920 115080 42080
rect 114920 42080 115080 42240
rect 114920 42240 115080 42400
rect 114920 42400 115080 42560
rect 114920 42560 115080 42720
rect 114920 42720 115080 42880
rect 114920 42880 115080 43040
rect 114920 43040 115080 43200
rect 114920 43200 115080 43360
rect 114920 43360 115080 43520
rect 114920 43520 115080 43680
rect 114920 43680 115080 43840
rect 114920 43840 115080 44000
rect 114920 44000 115080 44160
rect 114920 44160 115080 44320
rect 114920 44320 115080 44480
rect 114920 44480 115080 44640
rect 114920 44640 115080 44800
rect 114920 44800 115080 44960
rect 114920 44960 115080 45120
rect 114920 45120 115080 45280
rect 114920 45280 115080 45440
rect 114920 45440 115080 45600
rect 114920 45600 115080 45760
rect 114920 45760 115080 45920
rect 114920 49440 115080 49600
rect 114920 49600 115080 49760
rect 114920 49760 115080 49920
rect 114920 49920 115080 50080
rect 114920 50080 115080 50240
rect 114920 50240 115080 50400
rect 114920 50400 115080 50560
rect 114920 50560 115080 50720
rect 114920 50720 115080 50880
rect 114920 50880 115080 51040
rect 114920 51040 115080 51200
rect 114920 51200 115080 51360
rect 114920 51360 115080 51520
rect 114920 51520 115080 51680
rect 114920 51680 115080 51840
rect 114920 51840 115080 52000
rect 114920 52000 115080 52160
rect 114920 52160 115080 52320
rect 114920 52320 115080 52480
rect 114920 52480 115080 52640
rect 114920 52640 115080 52800
rect 114920 52800 115080 52960
rect 114920 52960 115080 53120
rect 115080 37920 115240 38080
rect 115080 38080 115240 38240
rect 115080 38240 115240 38400
rect 115080 38400 115240 38560
rect 115080 38560 115240 38720
rect 115080 38720 115240 38880
rect 115080 38880 115240 39040
rect 115080 39040 115240 39200
rect 115080 39200 115240 39360
rect 115080 39360 115240 39520
rect 115080 39520 115240 39680
rect 115080 39680 115240 39840
rect 115080 39840 115240 40000
rect 115080 40000 115240 40160
rect 115080 40160 115240 40320
rect 115080 40320 115240 40480
rect 115080 40480 115240 40640
rect 115080 40640 115240 40800
rect 115080 40800 115240 40960
rect 115080 40960 115240 41120
rect 115080 41120 115240 41280
rect 115080 41280 115240 41440
rect 115080 41440 115240 41600
rect 115080 41600 115240 41760
rect 115080 41760 115240 41920
rect 115080 41920 115240 42080
rect 115080 42080 115240 42240
rect 115080 42240 115240 42400
rect 115080 42400 115240 42560
rect 115080 42560 115240 42720
rect 115080 42720 115240 42880
rect 115080 42880 115240 43040
rect 115080 43040 115240 43200
rect 115080 43200 115240 43360
rect 115080 43360 115240 43520
rect 115080 43520 115240 43680
rect 115080 43680 115240 43840
rect 115080 43840 115240 44000
rect 115080 44000 115240 44160
rect 115080 44160 115240 44320
rect 115080 44320 115240 44480
rect 115080 44480 115240 44640
rect 115080 44640 115240 44800
rect 115080 44800 115240 44960
rect 115080 44960 115240 45120
rect 115080 45120 115240 45280
rect 115080 45280 115240 45440
rect 115080 45440 115240 45600
rect 115080 45600 115240 45760
rect 115080 45760 115240 45920
rect 115080 45920 115240 46080
rect 115080 46080 115240 46240
rect 115080 46240 115240 46400
rect 115080 46400 115240 46560
rect 115080 49120 115240 49280
rect 115080 49280 115240 49440
rect 115080 49440 115240 49600
rect 115080 49600 115240 49760
rect 115080 49760 115240 49920
rect 115080 49920 115240 50080
rect 115080 50080 115240 50240
rect 115080 50240 115240 50400
rect 115080 50400 115240 50560
rect 115080 50560 115240 50720
rect 115080 50720 115240 50880
rect 115080 50880 115240 51040
rect 115080 51040 115240 51200
rect 115080 51200 115240 51360
rect 115080 51360 115240 51520
rect 115080 51520 115240 51680
rect 115080 51680 115240 51840
rect 115080 51840 115240 52000
rect 115080 52000 115240 52160
rect 115080 52160 115240 52320
rect 115080 52320 115240 52480
rect 115080 52480 115240 52640
rect 115080 52640 115240 52800
rect 115080 52800 115240 52960
rect 115080 52960 115240 53120
rect 115080 53120 115240 53280
rect 115080 53280 115240 53440
rect 115240 38400 115400 38560
rect 115240 38560 115400 38720
rect 115240 38720 115400 38880
rect 115240 38880 115400 39040
rect 115240 39040 115400 39200
rect 115240 39200 115400 39360
rect 115240 39360 115400 39520
rect 115240 39520 115400 39680
rect 115240 39680 115400 39840
rect 115240 39840 115400 40000
rect 115240 40000 115400 40160
rect 115240 40160 115400 40320
rect 115240 40320 115400 40480
rect 115240 40480 115400 40640
rect 115240 40640 115400 40800
rect 115240 40800 115400 40960
rect 115240 40960 115400 41120
rect 115240 41120 115400 41280
rect 115240 41280 115400 41440
rect 115240 41440 115400 41600
rect 115240 41600 115400 41760
rect 115240 41760 115400 41920
rect 115240 41920 115400 42080
rect 115240 42080 115400 42240
rect 115240 42240 115400 42400
rect 115240 42400 115400 42560
rect 115240 42560 115400 42720
rect 115240 42720 115400 42880
rect 115240 42880 115400 43040
rect 115240 43040 115400 43200
rect 115240 43200 115400 43360
rect 115240 43360 115400 43520
rect 115240 43520 115400 43680
rect 115240 43680 115400 43840
rect 115240 43840 115400 44000
rect 115240 44000 115400 44160
rect 115240 44160 115400 44320
rect 115240 44320 115400 44480
rect 115240 44480 115400 44640
rect 115240 44640 115400 44800
rect 115240 44800 115400 44960
rect 115240 44960 115400 45120
rect 115240 45120 115400 45280
rect 115240 45280 115400 45440
rect 115240 45440 115400 45600
rect 115240 45600 115400 45760
rect 115240 45760 115400 45920
rect 115240 45920 115400 46080
rect 115240 46080 115400 46240
rect 115240 46240 115400 46400
rect 115240 46400 115400 46560
rect 115240 46560 115400 46720
rect 115240 46720 115400 46880
rect 115240 46880 115400 47040
rect 115240 47040 115400 47200
rect 115240 48640 115400 48800
rect 115240 48800 115400 48960
rect 115240 48960 115400 49120
rect 115240 49120 115400 49280
rect 115240 49280 115400 49440
rect 115240 49440 115400 49600
rect 115240 49600 115400 49760
rect 115240 49760 115400 49920
rect 115240 49920 115400 50080
rect 115240 50080 115400 50240
rect 115240 50240 115400 50400
rect 115240 50400 115400 50560
rect 115240 50560 115400 50720
rect 115240 50720 115400 50880
rect 115240 50880 115400 51040
rect 115240 51040 115400 51200
rect 115240 51200 115400 51360
rect 115240 51360 115400 51520
rect 115240 51520 115400 51680
rect 115240 51680 115400 51840
rect 115240 51840 115400 52000
rect 115240 52000 115400 52160
rect 115240 52160 115400 52320
rect 115240 52320 115400 52480
rect 115240 52480 115400 52640
rect 115240 52640 115400 52800
rect 115240 52800 115400 52960
rect 115240 52960 115400 53120
rect 115240 53120 115400 53280
rect 115240 53280 115400 53440
rect 115240 53440 115400 53600
rect 115400 38880 115560 39040
rect 115400 39040 115560 39200
rect 115400 39200 115560 39360
rect 115400 39360 115560 39520
rect 115400 39520 115560 39680
rect 115400 39680 115560 39840
rect 115400 39840 115560 40000
rect 115400 40000 115560 40160
rect 115400 40160 115560 40320
rect 115400 40320 115560 40480
rect 115400 40480 115560 40640
rect 115400 40640 115560 40800
rect 115400 40800 115560 40960
rect 115400 40960 115560 41120
rect 115400 41120 115560 41280
rect 115400 41280 115560 41440
rect 115400 41440 115560 41600
rect 115400 41600 115560 41760
rect 115400 41760 115560 41920
rect 115400 41920 115560 42080
rect 115400 42080 115560 42240
rect 115400 42240 115560 42400
rect 115400 42400 115560 42560
rect 115400 42560 115560 42720
rect 115400 42720 115560 42880
rect 115400 42880 115560 43040
rect 115400 43040 115560 43200
rect 115400 43200 115560 43360
rect 115400 43360 115560 43520
rect 115400 43520 115560 43680
rect 115400 43680 115560 43840
rect 115400 43840 115560 44000
rect 115400 44000 115560 44160
rect 115400 44160 115560 44320
rect 115400 44320 115560 44480
rect 115400 44480 115560 44640
rect 115400 44640 115560 44800
rect 115400 44800 115560 44960
rect 115400 44960 115560 45120
rect 115400 45120 115560 45280
rect 115400 45280 115560 45440
rect 115400 45440 115560 45600
rect 115400 45600 115560 45760
rect 115400 45760 115560 45920
rect 115400 45920 115560 46080
rect 115400 46080 115560 46240
rect 115400 46240 115560 46400
rect 115400 46400 115560 46560
rect 115400 46560 115560 46720
rect 115400 46720 115560 46880
rect 115400 46880 115560 47040
rect 115400 47040 115560 47200
rect 115400 47200 115560 47360
rect 115400 47360 115560 47520
rect 115400 47520 115560 47680
rect 115400 47680 115560 47840
rect 115400 47840 115560 48000
rect 115400 48000 115560 48160
rect 115400 48160 115560 48320
rect 115400 48320 115560 48480
rect 115400 48480 115560 48640
rect 115400 48640 115560 48800
rect 115400 48800 115560 48960
rect 115400 48960 115560 49120
rect 115400 49120 115560 49280
rect 115400 49280 115560 49440
rect 115400 49440 115560 49600
rect 115400 49600 115560 49760
rect 115400 49760 115560 49920
rect 115400 49920 115560 50080
rect 115400 50080 115560 50240
rect 115400 50240 115560 50400
rect 115400 50400 115560 50560
rect 115400 50560 115560 50720
rect 115400 50720 115560 50880
rect 115400 50880 115560 51040
rect 115400 51040 115560 51200
rect 115400 51200 115560 51360
rect 115400 51360 115560 51520
rect 115400 51520 115560 51680
rect 115400 51680 115560 51840
rect 115400 51840 115560 52000
rect 115400 52000 115560 52160
rect 115400 52160 115560 52320
rect 115400 52320 115560 52480
rect 115400 52480 115560 52640
rect 115400 52640 115560 52800
rect 115400 52800 115560 52960
rect 115400 52960 115560 53120
rect 115400 53120 115560 53280
rect 115400 53280 115560 53440
rect 115400 53440 115560 53600
rect 115400 53600 115560 53760
rect 115400 53760 115560 53920
rect 115560 39360 115720 39520
rect 115560 39520 115720 39680
rect 115560 39680 115720 39840
rect 115560 39840 115720 40000
rect 115560 40000 115720 40160
rect 115560 40160 115720 40320
rect 115560 40320 115720 40480
rect 115560 40480 115720 40640
rect 115560 40640 115720 40800
rect 115560 40800 115720 40960
rect 115560 40960 115720 41120
rect 115560 41120 115720 41280
rect 115560 41280 115720 41440
rect 115560 41440 115720 41600
rect 115560 41600 115720 41760
rect 115560 41760 115720 41920
rect 115560 41920 115720 42080
rect 115560 42080 115720 42240
rect 115560 42240 115720 42400
rect 115560 42400 115720 42560
rect 115560 42560 115720 42720
rect 115560 42720 115720 42880
rect 115560 42880 115720 43040
rect 115560 43040 115720 43200
rect 115560 43200 115720 43360
rect 115560 43360 115720 43520
rect 115560 43520 115720 43680
rect 115560 43680 115720 43840
rect 115560 43840 115720 44000
rect 115560 44000 115720 44160
rect 115560 44160 115720 44320
rect 115560 44320 115720 44480
rect 115560 44480 115720 44640
rect 115560 44640 115720 44800
rect 115560 44800 115720 44960
rect 115560 44960 115720 45120
rect 115560 45120 115720 45280
rect 115560 45280 115720 45440
rect 115560 45440 115720 45600
rect 115560 45600 115720 45760
rect 115560 45760 115720 45920
rect 115560 45920 115720 46080
rect 115560 46080 115720 46240
rect 115560 46240 115720 46400
rect 115560 46400 115720 46560
rect 115560 46560 115720 46720
rect 115560 46720 115720 46880
rect 115560 46880 115720 47040
rect 115560 47040 115720 47200
rect 115560 47200 115720 47360
rect 115560 47360 115720 47520
rect 115560 47520 115720 47680
rect 115560 47680 115720 47840
rect 115560 47840 115720 48000
rect 115560 48000 115720 48160
rect 115560 48160 115720 48320
rect 115560 48320 115720 48480
rect 115560 48480 115720 48640
rect 115560 48640 115720 48800
rect 115560 48800 115720 48960
rect 115560 48960 115720 49120
rect 115560 49120 115720 49280
rect 115560 49280 115720 49440
rect 115560 49440 115720 49600
rect 115560 49600 115720 49760
rect 115560 49760 115720 49920
rect 115560 49920 115720 50080
rect 115560 50080 115720 50240
rect 115560 50240 115720 50400
rect 115560 50400 115720 50560
rect 115560 50560 115720 50720
rect 115560 50720 115720 50880
rect 115560 50880 115720 51040
rect 115560 51040 115720 51200
rect 115560 51200 115720 51360
rect 115560 51360 115720 51520
rect 115560 51520 115720 51680
rect 115560 51680 115720 51840
rect 115560 51840 115720 52000
rect 115560 52000 115720 52160
rect 115560 52160 115720 52320
rect 115560 52320 115720 52480
rect 115560 52480 115720 52640
rect 115560 52640 115720 52800
rect 115560 52800 115720 52960
rect 115560 52960 115720 53120
rect 115560 53120 115720 53280
rect 115560 53280 115720 53440
rect 115560 53440 115720 53600
rect 115560 53600 115720 53760
rect 115560 53760 115720 53920
rect 115560 53920 115720 54080
rect 115720 39840 115880 40000
rect 115720 40000 115880 40160
rect 115720 40160 115880 40320
rect 115720 40320 115880 40480
rect 115720 40480 115880 40640
rect 115720 40640 115880 40800
rect 115720 40800 115880 40960
rect 115720 40960 115880 41120
rect 115720 41120 115880 41280
rect 115720 41280 115880 41440
rect 115720 41440 115880 41600
rect 115720 41600 115880 41760
rect 115720 41760 115880 41920
rect 115720 41920 115880 42080
rect 115720 42080 115880 42240
rect 115720 42240 115880 42400
rect 115720 42400 115880 42560
rect 115720 42560 115880 42720
rect 115720 42720 115880 42880
rect 115720 42880 115880 43040
rect 115720 43040 115880 43200
rect 115720 43200 115880 43360
rect 115720 43360 115880 43520
rect 115720 43520 115880 43680
rect 115720 43680 115880 43840
rect 115720 43840 115880 44000
rect 115720 44000 115880 44160
rect 115720 44160 115880 44320
rect 115720 44320 115880 44480
rect 115720 44480 115880 44640
rect 115720 44640 115880 44800
rect 115720 44800 115880 44960
rect 115720 44960 115880 45120
rect 115720 45120 115880 45280
rect 115720 45280 115880 45440
rect 115720 45440 115880 45600
rect 115720 45600 115880 45760
rect 115720 45760 115880 45920
rect 115720 45920 115880 46080
rect 115720 46080 115880 46240
rect 115720 46240 115880 46400
rect 115720 46400 115880 46560
rect 115720 46560 115880 46720
rect 115720 46720 115880 46880
rect 115720 46880 115880 47040
rect 115720 47040 115880 47200
rect 115720 47200 115880 47360
rect 115720 47360 115880 47520
rect 115720 47520 115880 47680
rect 115720 47680 115880 47840
rect 115720 47840 115880 48000
rect 115720 48000 115880 48160
rect 115720 48160 115880 48320
rect 115720 48320 115880 48480
rect 115720 48480 115880 48640
rect 115720 48640 115880 48800
rect 115720 48800 115880 48960
rect 115720 48960 115880 49120
rect 115720 49120 115880 49280
rect 115720 49280 115880 49440
rect 115720 49440 115880 49600
rect 115720 49600 115880 49760
rect 115720 49760 115880 49920
rect 115720 49920 115880 50080
rect 115720 50080 115880 50240
rect 115720 50240 115880 50400
rect 115720 50400 115880 50560
rect 115720 50560 115880 50720
rect 115720 50720 115880 50880
rect 115720 50880 115880 51040
rect 115720 51040 115880 51200
rect 115720 51200 115880 51360
rect 115720 51360 115880 51520
rect 115720 51520 115880 51680
rect 115720 51680 115880 51840
rect 115720 51840 115880 52000
rect 115720 52000 115880 52160
rect 115720 52160 115880 52320
rect 115720 52320 115880 52480
rect 115720 52480 115880 52640
rect 115720 52640 115880 52800
rect 115720 52800 115880 52960
rect 115720 52960 115880 53120
rect 115720 53120 115880 53280
rect 115720 53280 115880 53440
rect 115720 53440 115880 53600
rect 115720 53600 115880 53760
rect 115720 53760 115880 53920
rect 115720 53920 115880 54080
rect 115720 54080 115880 54240
rect 115880 40160 116040 40320
rect 115880 40320 116040 40480
rect 115880 40480 116040 40640
rect 115880 40640 116040 40800
rect 115880 40800 116040 40960
rect 115880 40960 116040 41120
rect 115880 41120 116040 41280
rect 115880 41280 116040 41440
rect 115880 41440 116040 41600
rect 115880 41600 116040 41760
rect 115880 41760 116040 41920
rect 115880 41920 116040 42080
rect 115880 42080 116040 42240
rect 115880 42240 116040 42400
rect 115880 42400 116040 42560
rect 115880 42560 116040 42720
rect 115880 42720 116040 42880
rect 115880 42880 116040 43040
rect 115880 43040 116040 43200
rect 115880 43200 116040 43360
rect 115880 43360 116040 43520
rect 115880 43520 116040 43680
rect 115880 43680 116040 43840
rect 115880 43840 116040 44000
rect 115880 44000 116040 44160
rect 115880 44160 116040 44320
rect 115880 44320 116040 44480
rect 115880 44480 116040 44640
rect 115880 44640 116040 44800
rect 115880 44800 116040 44960
rect 115880 44960 116040 45120
rect 115880 45120 116040 45280
rect 115880 45280 116040 45440
rect 115880 45440 116040 45600
rect 115880 45600 116040 45760
rect 115880 45760 116040 45920
rect 115880 45920 116040 46080
rect 115880 46080 116040 46240
rect 115880 46240 116040 46400
rect 115880 46400 116040 46560
rect 115880 46560 116040 46720
rect 115880 46720 116040 46880
rect 115880 46880 116040 47040
rect 115880 47040 116040 47200
rect 115880 47200 116040 47360
rect 115880 47360 116040 47520
rect 115880 47520 116040 47680
rect 115880 47680 116040 47840
rect 115880 47840 116040 48000
rect 115880 48000 116040 48160
rect 115880 48160 116040 48320
rect 115880 48320 116040 48480
rect 115880 48480 116040 48640
rect 115880 48640 116040 48800
rect 115880 48800 116040 48960
rect 115880 48960 116040 49120
rect 115880 49120 116040 49280
rect 115880 49280 116040 49440
rect 115880 49440 116040 49600
rect 115880 49600 116040 49760
rect 115880 49760 116040 49920
rect 115880 49920 116040 50080
rect 115880 50080 116040 50240
rect 115880 50240 116040 50400
rect 115880 50400 116040 50560
rect 115880 50560 116040 50720
rect 115880 50720 116040 50880
rect 115880 50880 116040 51040
rect 115880 51040 116040 51200
rect 115880 51200 116040 51360
rect 115880 51360 116040 51520
rect 115880 51520 116040 51680
rect 115880 51680 116040 51840
rect 115880 51840 116040 52000
rect 115880 52000 116040 52160
rect 115880 52160 116040 52320
rect 115880 52320 116040 52480
rect 115880 52480 116040 52640
rect 115880 52640 116040 52800
rect 115880 52800 116040 52960
rect 115880 52960 116040 53120
rect 115880 53120 116040 53280
rect 115880 53280 116040 53440
rect 115880 53440 116040 53600
rect 115880 53600 116040 53760
rect 115880 53760 116040 53920
rect 115880 53920 116040 54080
rect 115880 54080 116040 54240
rect 115880 54240 116040 54400
rect 116040 40640 116200 40800
rect 116040 40800 116200 40960
rect 116040 40960 116200 41120
rect 116040 41120 116200 41280
rect 116040 41280 116200 41440
rect 116040 41440 116200 41600
rect 116040 41600 116200 41760
rect 116040 41760 116200 41920
rect 116040 41920 116200 42080
rect 116040 42080 116200 42240
rect 116040 42240 116200 42400
rect 116040 42400 116200 42560
rect 116040 42560 116200 42720
rect 116040 42720 116200 42880
rect 116040 42880 116200 43040
rect 116040 43040 116200 43200
rect 116040 43200 116200 43360
rect 116040 43360 116200 43520
rect 116040 43520 116200 43680
rect 116040 43680 116200 43840
rect 116040 43840 116200 44000
rect 116040 44000 116200 44160
rect 116040 44160 116200 44320
rect 116040 44320 116200 44480
rect 116040 44480 116200 44640
rect 116040 44640 116200 44800
rect 116040 44800 116200 44960
rect 116040 44960 116200 45120
rect 116040 45120 116200 45280
rect 116040 45280 116200 45440
rect 116040 45440 116200 45600
rect 116040 45600 116200 45760
rect 116040 45760 116200 45920
rect 116040 45920 116200 46080
rect 116040 46080 116200 46240
rect 116040 46240 116200 46400
rect 116040 46400 116200 46560
rect 116040 46560 116200 46720
rect 116040 46720 116200 46880
rect 116040 46880 116200 47040
rect 116040 47040 116200 47200
rect 116040 47200 116200 47360
rect 116040 47360 116200 47520
rect 116040 47520 116200 47680
rect 116040 47680 116200 47840
rect 116040 47840 116200 48000
rect 116040 48000 116200 48160
rect 116040 48160 116200 48320
rect 116040 48320 116200 48480
rect 116040 48480 116200 48640
rect 116040 48640 116200 48800
rect 116040 48800 116200 48960
rect 116040 48960 116200 49120
rect 116040 49120 116200 49280
rect 116040 49280 116200 49440
rect 116040 49440 116200 49600
rect 116040 49600 116200 49760
rect 116040 49760 116200 49920
rect 116040 49920 116200 50080
rect 116040 50080 116200 50240
rect 116040 50240 116200 50400
rect 116040 50400 116200 50560
rect 116040 50560 116200 50720
rect 116040 50720 116200 50880
rect 116040 50880 116200 51040
rect 116040 51040 116200 51200
rect 116040 51200 116200 51360
rect 116040 51360 116200 51520
rect 116040 51520 116200 51680
rect 116040 51680 116200 51840
rect 116040 51840 116200 52000
rect 116040 52000 116200 52160
rect 116040 52160 116200 52320
rect 116040 52320 116200 52480
rect 116040 52480 116200 52640
rect 116040 52640 116200 52800
rect 116040 52800 116200 52960
rect 116040 52960 116200 53120
rect 116040 53120 116200 53280
rect 116040 53280 116200 53440
rect 116040 53440 116200 53600
rect 116040 53600 116200 53760
rect 116040 53760 116200 53920
rect 116040 53920 116200 54080
rect 116040 54080 116200 54240
rect 116040 54240 116200 54400
rect 116200 41120 116360 41280
rect 116200 41280 116360 41440
rect 116200 41440 116360 41600
rect 116200 41600 116360 41760
rect 116200 41760 116360 41920
rect 116200 41920 116360 42080
rect 116200 42080 116360 42240
rect 116200 42240 116360 42400
rect 116200 42400 116360 42560
rect 116200 42560 116360 42720
rect 116200 42720 116360 42880
rect 116200 42880 116360 43040
rect 116200 43040 116360 43200
rect 116200 43200 116360 43360
rect 116200 43360 116360 43520
rect 116200 43520 116360 43680
rect 116200 43680 116360 43840
rect 116200 43840 116360 44000
rect 116200 44000 116360 44160
rect 116200 44160 116360 44320
rect 116200 44320 116360 44480
rect 116200 44480 116360 44640
rect 116200 44640 116360 44800
rect 116200 44800 116360 44960
rect 116200 44960 116360 45120
rect 116200 45120 116360 45280
rect 116200 45280 116360 45440
rect 116200 45440 116360 45600
rect 116200 45600 116360 45760
rect 116200 45760 116360 45920
rect 116200 45920 116360 46080
rect 116200 46080 116360 46240
rect 116200 46240 116360 46400
rect 116200 46400 116360 46560
rect 116200 46560 116360 46720
rect 116200 46720 116360 46880
rect 116200 46880 116360 47040
rect 116200 47040 116360 47200
rect 116200 47200 116360 47360
rect 116200 47360 116360 47520
rect 116200 47520 116360 47680
rect 116200 47680 116360 47840
rect 116200 47840 116360 48000
rect 116200 48000 116360 48160
rect 116200 48160 116360 48320
rect 116200 48320 116360 48480
rect 116200 48480 116360 48640
rect 116200 48640 116360 48800
rect 116200 48800 116360 48960
rect 116200 48960 116360 49120
rect 116200 49120 116360 49280
rect 116200 49280 116360 49440
rect 116200 49440 116360 49600
rect 116200 49600 116360 49760
rect 116200 49760 116360 49920
rect 116200 49920 116360 50080
rect 116200 50080 116360 50240
rect 116200 50240 116360 50400
rect 116200 50400 116360 50560
rect 116200 50560 116360 50720
rect 116200 50720 116360 50880
rect 116200 50880 116360 51040
rect 116200 51040 116360 51200
rect 116200 51200 116360 51360
rect 116200 51360 116360 51520
rect 116200 51520 116360 51680
rect 116200 51680 116360 51840
rect 116200 51840 116360 52000
rect 116200 52000 116360 52160
rect 116200 52160 116360 52320
rect 116200 52320 116360 52480
rect 116200 52480 116360 52640
rect 116200 52640 116360 52800
rect 116200 52800 116360 52960
rect 116200 52960 116360 53120
rect 116200 53120 116360 53280
rect 116200 53280 116360 53440
rect 116200 53440 116360 53600
rect 116200 53600 116360 53760
rect 116200 53760 116360 53920
rect 116200 53920 116360 54080
rect 116200 54080 116360 54240
rect 116200 54240 116360 54400
rect 116200 54400 116360 54560
rect 116360 41440 116520 41600
rect 116360 41600 116520 41760
rect 116360 41760 116520 41920
rect 116360 41920 116520 42080
rect 116360 42080 116520 42240
rect 116360 42240 116520 42400
rect 116360 42400 116520 42560
rect 116360 42560 116520 42720
rect 116360 42720 116520 42880
rect 116360 42880 116520 43040
rect 116360 43040 116520 43200
rect 116360 43200 116520 43360
rect 116360 43360 116520 43520
rect 116360 43520 116520 43680
rect 116360 43680 116520 43840
rect 116360 43840 116520 44000
rect 116360 44000 116520 44160
rect 116360 44160 116520 44320
rect 116360 44320 116520 44480
rect 116360 44480 116520 44640
rect 116360 44640 116520 44800
rect 116360 44800 116520 44960
rect 116360 44960 116520 45120
rect 116360 45120 116520 45280
rect 116360 45280 116520 45440
rect 116360 45440 116520 45600
rect 116360 45600 116520 45760
rect 116360 45760 116520 45920
rect 116360 45920 116520 46080
rect 116360 46080 116520 46240
rect 116360 46240 116520 46400
rect 116360 46400 116520 46560
rect 116360 46560 116520 46720
rect 116360 46720 116520 46880
rect 116360 46880 116520 47040
rect 116360 47040 116520 47200
rect 116360 47200 116520 47360
rect 116360 47360 116520 47520
rect 116360 47520 116520 47680
rect 116360 47680 116520 47840
rect 116360 47840 116520 48000
rect 116360 48000 116520 48160
rect 116360 48160 116520 48320
rect 116360 48320 116520 48480
rect 116360 48480 116520 48640
rect 116360 48640 116520 48800
rect 116360 48800 116520 48960
rect 116360 48960 116520 49120
rect 116360 49120 116520 49280
rect 116360 49280 116520 49440
rect 116360 49440 116520 49600
rect 116360 49600 116520 49760
rect 116360 49760 116520 49920
rect 116360 49920 116520 50080
rect 116360 50080 116520 50240
rect 116360 50240 116520 50400
rect 116360 50400 116520 50560
rect 116360 50560 116520 50720
rect 116360 50720 116520 50880
rect 116360 50880 116520 51040
rect 116360 51040 116520 51200
rect 116360 51200 116520 51360
rect 116360 51360 116520 51520
rect 116360 51520 116520 51680
rect 116360 51680 116520 51840
rect 116360 51840 116520 52000
rect 116360 52000 116520 52160
rect 116360 52160 116520 52320
rect 116360 52320 116520 52480
rect 116360 52480 116520 52640
rect 116360 52640 116520 52800
rect 116360 52800 116520 52960
rect 116360 52960 116520 53120
rect 116360 53120 116520 53280
rect 116360 53280 116520 53440
rect 116360 53440 116520 53600
rect 116360 53600 116520 53760
rect 116360 53760 116520 53920
rect 116360 53920 116520 54080
rect 116360 54080 116520 54240
rect 116360 54240 116520 54400
rect 116360 54400 116520 54560
rect 116360 54560 116520 54720
rect 116520 41920 116680 42080
rect 116520 42080 116680 42240
rect 116520 42240 116680 42400
rect 116520 42400 116680 42560
rect 116520 42560 116680 42720
rect 116520 42720 116680 42880
rect 116520 42880 116680 43040
rect 116520 43040 116680 43200
rect 116520 43200 116680 43360
rect 116520 43360 116680 43520
rect 116520 43520 116680 43680
rect 116520 43680 116680 43840
rect 116520 43840 116680 44000
rect 116520 44000 116680 44160
rect 116520 44160 116680 44320
rect 116520 44320 116680 44480
rect 116520 44480 116680 44640
rect 116520 44640 116680 44800
rect 116520 44800 116680 44960
rect 116520 44960 116680 45120
rect 116520 45120 116680 45280
rect 116520 45280 116680 45440
rect 116520 45440 116680 45600
rect 116520 45600 116680 45760
rect 116520 45760 116680 45920
rect 116520 45920 116680 46080
rect 116520 46080 116680 46240
rect 116520 46240 116680 46400
rect 116520 46400 116680 46560
rect 116520 46560 116680 46720
rect 116520 46720 116680 46880
rect 116520 46880 116680 47040
rect 116520 47040 116680 47200
rect 116520 47200 116680 47360
rect 116520 47360 116680 47520
rect 116520 47520 116680 47680
rect 116520 47680 116680 47840
rect 116520 47840 116680 48000
rect 116520 48000 116680 48160
rect 116520 48160 116680 48320
rect 116520 48320 116680 48480
rect 116520 48480 116680 48640
rect 116520 48640 116680 48800
rect 116520 48800 116680 48960
rect 116520 48960 116680 49120
rect 116520 49120 116680 49280
rect 116520 49280 116680 49440
rect 116520 49440 116680 49600
rect 116520 49600 116680 49760
rect 116520 49760 116680 49920
rect 116520 49920 116680 50080
rect 116520 50080 116680 50240
rect 116520 50240 116680 50400
rect 116520 50400 116680 50560
rect 116520 50560 116680 50720
rect 116520 50720 116680 50880
rect 116520 50880 116680 51040
rect 116520 51040 116680 51200
rect 116520 51200 116680 51360
rect 116520 51360 116680 51520
rect 116520 51520 116680 51680
rect 116520 51680 116680 51840
rect 116520 51840 116680 52000
rect 116520 52000 116680 52160
rect 116520 52160 116680 52320
rect 116520 52320 116680 52480
rect 116520 52480 116680 52640
rect 116520 52640 116680 52800
rect 116520 52800 116680 52960
rect 116520 52960 116680 53120
rect 116520 53120 116680 53280
rect 116520 53280 116680 53440
rect 116520 53440 116680 53600
rect 116520 53600 116680 53760
rect 116520 53760 116680 53920
rect 116520 53920 116680 54080
rect 116520 54080 116680 54240
rect 116520 54240 116680 54400
rect 116520 54400 116680 54560
rect 116520 54560 116680 54720
rect 116680 42400 116840 42560
rect 116680 42560 116840 42720
rect 116680 42720 116840 42880
rect 116680 42880 116840 43040
rect 116680 43040 116840 43200
rect 116680 43200 116840 43360
rect 116680 43360 116840 43520
rect 116680 43520 116840 43680
rect 116680 43680 116840 43840
rect 116680 43840 116840 44000
rect 116680 44000 116840 44160
rect 116680 44160 116840 44320
rect 116680 44320 116840 44480
rect 116680 44480 116840 44640
rect 116680 44640 116840 44800
rect 116680 44800 116840 44960
rect 116680 44960 116840 45120
rect 116680 45120 116840 45280
rect 116680 45280 116840 45440
rect 116680 45440 116840 45600
rect 116680 45600 116840 45760
rect 116680 45760 116840 45920
rect 116680 45920 116840 46080
rect 116680 46080 116840 46240
rect 116680 46240 116840 46400
rect 116680 46400 116840 46560
rect 116680 46560 116840 46720
rect 116680 46720 116840 46880
rect 116680 46880 116840 47040
rect 116680 47040 116840 47200
rect 116680 47200 116840 47360
rect 116680 47360 116840 47520
rect 116680 47520 116840 47680
rect 116680 47680 116840 47840
rect 116680 47840 116840 48000
rect 116680 48000 116840 48160
rect 116680 48160 116840 48320
rect 116680 48320 116840 48480
rect 116680 48480 116840 48640
rect 116680 48640 116840 48800
rect 116680 48800 116840 48960
rect 116680 48960 116840 49120
rect 116680 49120 116840 49280
rect 116680 49280 116840 49440
rect 116680 49440 116840 49600
rect 116680 49600 116840 49760
rect 116680 49760 116840 49920
rect 116680 49920 116840 50080
rect 116680 50080 116840 50240
rect 116680 50240 116840 50400
rect 116680 50400 116840 50560
rect 116680 50560 116840 50720
rect 116680 50720 116840 50880
rect 116680 50880 116840 51040
rect 116680 51040 116840 51200
rect 116680 51200 116840 51360
rect 116680 51360 116840 51520
rect 116680 51520 116840 51680
rect 116680 51680 116840 51840
rect 116680 51840 116840 52000
rect 116680 52000 116840 52160
rect 116680 52160 116840 52320
rect 116680 52320 116840 52480
rect 116680 52480 116840 52640
rect 116680 52640 116840 52800
rect 116680 52800 116840 52960
rect 116680 52960 116840 53120
rect 116680 53120 116840 53280
rect 116680 53280 116840 53440
rect 116680 53440 116840 53600
rect 116680 53600 116840 53760
rect 116680 53760 116840 53920
rect 116680 53920 116840 54080
rect 116680 54080 116840 54240
rect 116680 54240 116840 54400
rect 116680 54400 116840 54560
rect 116680 54560 116840 54720
rect 116680 54720 116840 54880
rect 116840 42720 117000 42880
rect 116840 42880 117000 43040
rect 116840 43040 117000 43200
rect 116840 43200 117000 43360
rect 116840 43360 117000 43520
rect 116840 43520 117000 43680
rect 116840 43680 117000 43840
rect 116840 43840 117000 44000
rect 116840 44000 117000 44160
rect 116840 44160 117000 44320
rect 116840 44320 117000 44480
rect 116840 44480 117000 44640
rect 116840 44640 117000 44800
rect 116840 44800 117000 44960
rect 116840 44960 117000 45120
rect 116840 45120 117000 45280
rect 116840 45280 117000 45440
rect 116840 45440 117000 45600
rect 116840 45600 117000 45760
rect 116840 45760 117000 45920
rect 116840 45920 117000 46080
rect 116840 46080 117000 46240
rect 116840 46240 117000 46400
rect 116840 46400 117000 46560
rect 116840 46560 117000 46720
rect 116840 46720 117000 46880
rect 116840 46880 117000 47040
rect 116840 47040 117000 47200
rect 116840 47200 117000 47360
rect 116840 47360 117000 47520
rect 116840 47520 117000 47680
rect 116840 47680 117000 47840
rect 116840 47840 117000 48000
rect 116840 48000 117000 48160
rect 116840 48160 117000 48320
rect 116840 48320 117000 48480
rect 116840 48480 117000 48640
rect 116840 48640 117000 48800
rect 116840 48800 117000 48960
rect 116840 48960 117000 49120
rect 116840 49120 117000 49280
rect 116840 49280 117000 49440
rect 116840 49440 117000 49600
rect 116840 49600 117000 49760
rect 116840 49760 117000 49920
rect 116840 49920 117000 50080
rect 116840 50080 117000 50240
rect 116840 50240 117000 50400
rect 116840 50400 117000 50560
rect 116840 50560 117000 50720
rect 116840 50720 117000 50880
rect 116840 50880 117000 51040
rect 116840 51040 117000 51200
rect 116840 51200 117000 51360
rect 116840 51360 117000 51520
rect 116840 51520 117000 51680
rect 116840 51680 117000 51840
rect 116840 51840 117000 52000
rect 116840 52000 117000 52160
rect 116840 52160 117000 52320
rect 116840 52320 117000 52480
rect 116840 52480 117000 52640
rect 116840 52640 117000 52800
rect 116840 52800 117000 52960
rect 116840 52960 117000 53120
rect 116840 53120 117000 53280
rect 116840 53280 117000 53440
rect 116840 53440 117000 53600
rect 116840 53600 117000 53760
rect 116840 53760 117000 53920
rect 116840 53920 117000 54080
rect 116840 54080 117000 54240
rect 116840 54240 117000 54400
rect 116840 54400 117000 54560
rect 116840 54560 117000 54720
rect 116840 54720 117000 54880
rect 117000 43200 117160 43360
rect 117000 43360 117160 43520
rect 117000 43520 117160 43680
rect 117000 43680 117160 43840
rect 117000 43840 117160 44000
rect 117000 44000 117160 44160
rect 117000 44160 117160 44320
rect 117000 44320 117160 44480
rect 117000 44480 117160 44640
rect 117000 44640 117160 44800
rect 117000 44800 117160 44960
rect 117000 44960 117160 45120
rect 117000 45120 117160 45280
rect 117000 45280 117160 45440
rect 117000 45440 117160 45600
rect 117000 45600 117160 45760
rect 117000 45760 117160 45920
rect 117000 45920 117160 46080
rect 117000 46080 117160 46240
rect 117000 46240 117160 46400
rect 117000 46400 117160 46560
rect 117000 46560 117160 46720
rect 117000 46720 117160 46880
rect 117000 46880 117160 47040
rect 117000 47040 117160 47200
rect 117000 47200 117160 47360
rect 117000 47360 117160 47520
rect 117000 47520 117160 47680
rect 117000 47680 117160 47840
rect 117000 47840 117160 48000
rect 117000 48000 117160 48160
rect 117000 48160 117160 48320
rect 117000 48320 117160 48480
rect 117000 48480 117160 48640
rect 117000 48640 117160 48800
rect 117000 48800 117160 48960
rect 117000 48960 117160 49120
rect 117000 49120 117160 49280
rect 117000 49280 117160 49440
rect 117000 49440 117160 49600
rect 117000 49600 117160 49760
rect 117000 49760 117160 49920
rect 117000 49920 117160 50080
rect 117000 50080 117160 50240
rect 117000 50240 117160 50400
rect 117000 50400 117160 50560
rect 117000 50560 117160 50720
rect 117000 50720 117160 50880
rect 117000 50880 117160 51040
rect 117000 51040 117160 51200
rect 117000 51200 117160 51360
rect 117000 51360 117160 51520
rect 117000 51520 117160 51680
rect 117000 51680 117160 51840
rect 117000 51840 117160 52000
rect 117000 52000 117160 52160
rect 117000 52160 117160 52320
rect 117000 52320 117160 52480
rect 117000 52480 117160 52640
rect 117000 52640 117160 52800
rect 117000 52800 117160 52960
rect 117000 52960 117160 53120
rect 117000 53120 117160 53280
rect 117000 53280 117160 53440
rect 117000 53440 117160 53600
rect 117000 53600 117160 53760
rect 117000 53760 117160 53920
rect 117000 53920 117160 54080
rect 117000 54080 117160 54240
rect 117000 54240 117160 54400
rect 117000 54400 117160 54560
rect 117000 54560 117160 54720
rect 117000 54720 117160 54880
rect 117160 43520 117320 43680
rect 117160 43680 117320 43840
rect 117160 43840 117320 44000
rect 117160 44000 117320 44160
rect 117160 44160 117320 44320
rect 117160 44320 117320 44480
rect 117160 44480 117320 44640
rect 117160 44640 117320 44800
rect 117160 44800 117320 44960
rect 117160 44960 117320 45120
rect 117160 45120 117320 45280
rect 117160 45280 117320 45440
rect 117160 45440 117320 45600
rect 117160 45600 117320 45760
rect 117160 45760 117320 45920
rect 117160 45920 117320 46080
rect 117160 46080 117320 46240
rect 117160 46240 117320 46400
rect 117160 46400 117320 46560
rect 117160 46560 117320 46720
rect 117160 46720 117320 46880
rect 117160 46880 117320 47040
rect 117160 47040 117320 47200
rect 117160 47200 117320 47360
rect 117160 47360 117320 47520
rect 117160 47520 117320 47680
rect 117160 47680 117320 47840
rect 117160 47840 117320 48000
rect 117160 48000 117320 48160
rect 117160 48160 117320 48320
rect 117160 48320 117320 48480
rect 117160 48480 117320 48640
rect 117160 48640 117320 48800
rect 117160 48800 117320 48960
rect 117160 48960 117320 49120
rect 117160 49120 117320 49280
rect 117160 49280 117320 49440
rect 117160 49440 117320 49600
rect 117160 49600 117320 49760
rect 117160 49760 117320 49920
rect 117160 49920 117320 50080
rect 117160 50080 117320 50240
rect 117160 50240 117320 50400
rect 117160 50400 117320 50560
rect 117160 50560 117320 50720
rect 117160 51680 117320 51840
rect 117160 51840 117320 52000
rect 117160 52000 117320 52160
rect 117160 52160 117320 52320
rect 117160 52320 117320 52480
rect 117160 52480 117320 52640
rect 117160 52640 117320 52800
rect 117160 52800 117320 52960
rect 117160 52960 117320 53120
rect 117160 53120 117320 53280
rect 117160 53280 117320 53440
rect 117160 53440 117320 53600
rect 117160 53600 117320 53760
rect 117160 53760 117320 53920
rect 117160 53920 117320 54080
rect 117160 54080 117320 54240
rect 117160 54240 117320 54400
rect 117160 54400 117320 54560
rect 117160 54560 117320 54720
rect 117160 54720 117320 54880
rect 117160 54880 117320 55040
rect 117320 44000 117480 44160
rect 117320 44160 117480 44320
rect 117320 44320 117480 44480
rect 117320 44480 117480 44640
rect 117320 44640 117480 44800
rect 117320 44800 117480 44960
rect 117320 44960 117480 45120
rect 117320 45120 117480 45280
rect 117320 45280 117480 45440
rect 117320 45440 117480 45600
rect 117320 45600 117480 45760
rect 117320 45760 117480 45920
rect 117320 45920 117480 46080
rect 117320 46080 117480 46240
rect 117320 46240 117480 46400
rect 117320 46400 117480 46560
rect 117320 46560 117480 46720
rect 117320 46720 117480 46880
rect 117320 46880 117480 47040
rect 117320 47040 117480 47200
rect 117320 47200 117480 47360
rect 117320 47360 117480 47520
rect 117320 47520 117480 47680
rect 117320 47680 117480 47840
rect 117320 47840 117480 48000
rect 117320 48000 117480 48160
rect 117320 48160 117480 48320
rect 117320 48320 117480 48480
rect 117320 48480 117480 48640
rect 117320 48640 117480 48800
rect 117320 48800 117480 48960
rect 117320 48960 117480 49120
rect 117320 49120 117480 49280
rect 117320 49280 117480 49440
rect 117320 49440 117480 49600
rect 117320 49600 117480 49760
rect 117320 49760 117480 49920
rect 117320 49920 117480 50080
rect 117320 50080 117480 50240
rect 117320 50240 117480 50400
rect 117320 51840 117480 52000
rect 117320 52000 117480 52160
rect 117320 52160 117480 52320
rect 117320 52320 117480 52480
rect 117320 52480 117480 52640
rect 117320 52640 117480 52800
rect 117320 52800 117480 52960
rect 117320 52960 117480 53120
rect 117320 53120 117480 53280
rect 117320 53280 117480 53440
rect 117320 53440 117480 53600
rect 117320 53600 117480 53760
rect 117320 53760 117480 53920
rect 117320 53920 117480 54080
rect 117320 54080 117480 54240
rect 117320 54240 117480 54400
rect 117320 54400 117480 54560
rect 117320 54560 117480 54720
rect 117320 54720 117480 54880
rect 117320 54880 117480 55040
rect 117480 44320 117640 44480
rect 117480 44480 117640 44640
rect 117480 44640 117640 44800
rect 117480 44800 117640 44960
rect 117480 44960 117640 45120
rect 117480 45120 117640 45280
rect 117480 45280 117640 45440
rect 117480 45440 117640 45600
rect 117480 45600 117640 45760
rect 117480 45760 117640 45920
rect 117480 45920 117640 46080
rect 117480 46080 117640 46240
rect 117480 46240 117640 46400
rect 117480 46400 117640 46560
rect 117480 46560 117640 46720
rect 117480 46720 117640 46880
rect 117480 46880 117640 47040
rect 117480 47040 117640 47200
rect 117480 47200 117640 47360
rect 117480 47360 117640 47520
rect 117480 47520 117640 47680
rect 117480 47680 117640 47840
rect 117480 47840 117640 48000
rect 117480 48000 117640 48160
rect 117480 48160 117640 48320
rect 117480 48320 117640 48480
rect 117480 48480 117640 48640
rect 117480 48640 117640 48800
rect 117480 48800 117640 48960
rect 117480 48960 117640 49120
rect 117480 49120 117640 49280
rect 117480 49280 117640 49440
rect 117480 49440 117640 49600
rect 117480 49600 117640 49760
rect 117480 49760 117640 49920
rect 117480 49920 117640 50080
rect 117480 50080 117640 50240
rect 117480 52000 117640 52160
rect 117480 52160 117640 52320
rect 117480 52320 117640 52480
rect 117480 52480 117640 52640
rect 117480 52640 117640 52800
rect 117480 52800 117640 52960
rect 117480 52960 117640 53120
rect 117480 53120 117640 53280
rect 117480 53280 117640 53440
rect 117480 53440 117640 53600
rect 117480 53600 117640 53760
rect 117480 53760 117640 53920
rect 117480 53920 117640 54080
rect 117480 54080 117640 54240
rect 117480 54240 117640 54400
rect 117480 54400 117640 54560
rect 117480 54560 117640 54720
rect 117480 54720 117640 54880
rect 117480 54880 117640 55040
rect 117640 44640 117800 44800
rect 117640 44800 117800 44960
rect 117640 44960 117800 45120
rect 117640 45120 117800 45280
rect 117640 45280 117800 45440
rect 117640 45440 117800 45600
rect 117640 45600 117800 45760
rect 117640 45760 117800 45920
rect 117640 45920 117800 46080
rect 117640 46080 117800 46240
rect 117640 46240 117800 46400
rect 117640 46400 117800 46560
rect 117640 46560 117800 46720
rect 117640 46720 117800 46880
rect 117640 46880 117800 47040
rect 117640 47040 117800 47200
rect 117640 47200 117800 47360
rect 117640 47360 117800 47520
rect 117640 47520 117800 47680
rect 117640 47680 117800 47840
rect 117640 47840 117800 48000
rect 117640 48000 117800 48160
rect 117640 48160 117800 48320
rect 117640 48320 117800 48480
rect 117640 48480 117800 48640
rect 117640 48640 117800 48800
rect 117640 48800 117800 48960
rect 117640 48960 117800 49120
rect 117640 49120 117800 49280
rect 117640 49280 117800 49440
rect 117640 49440 117800 49600
rect 117640 49600 117800 49760
rect 117640 49760 117800 49920
rect 117640 49920 117800 50080
rect 117640 50080 117800 50240
rect 117640 52000 117800 52160
rect 117640 52160 117800 52320
rect 117640 52320 117800 52480
rect 117640 52480 117800 52640
rect 117640 52640 117800 52800
rect 117640 52800 117800 52960
rect 117640 52960 117800 53120
rect 117640 53120 117800 53280
rect 117640 53280 117800 53440
rect 117640 53440 117800 53600
rect 117640 53600 117800 53760
rect 117640 53760 117800 53920
rect 117640 53920 117800 54080
rect 117640 54080 117800 54240
rect 117640 54240 117800 54400
rect 117640 54400 117800 54560
rect 117640 54560 117800 54720
rect 117640 54720 117800 54880
rect 117640 54880 117800 55040
rect 117800 45120 117960 45280
rect 117800 45280 117960 45440
rect 117800 45440 117960 45600
rect 117800 45600 117960 45760
rect 117800 45760 117960 45920
rect 117800 45920 117960 46080
rect 117800 46080 117960 46240
rect 117800 46240 117960 46400
rect 117800 46400 117960 46560
rect 117800 46560 117960 46720
rect 117800 46720 117960 46880
rect 117800 46880 117960 47040
rect 117800 47040 117960 47200
rect 117800 47200 117960 47360
rect 117800 47360 117960 47520
rect 117800 47520 117960 47680
rect 117800 47680 117960 47840
rect 117800 47840 117960 48000
rect 117800 48000 117960 48160
rect 117800 48160 117960 48320
rect 117800 48320 117960 48480
rect 117800 48480 117960 48640
rect 117800 48640 117960 48800
rect 117800 48800 117960 48960
rect 117800 48960 117960 49120
rect 117800 49120 117960 49280
rect 117800 49280 117960 49440
rect 117800 49440 117960 49600
rect 117800 49600 117960 49760
rect 117800 49760 117960 49920
rect 117800 49920 117960 50080
rect 117800 52160 117960 52320
rect 117800 52320 117960 52480
rect 117800 52480 117960 52640
rect 117800 52640 117960 52800
rect 117800 52800 117960 52960
rect 117800 52960 117960 53120
rect 117800 53120 117960 53280
rect 117800 53280 117960 53440
rect 117800 53440 117960 53600
rect 117800 53600 117960 53760
rect 117800 53760 117960 53920
rect 117800 53920 117960 54080
rect 117800 54080 117960 54240
rect 117800 54240 117960 54400
rect 117800 54400 117960 54560
rect 117800 54560 117960 54720
rect 117800 54720 117960 54880
rect 117800 54880 117960 55040
rect 117800 55040 117960 55200
rect 117960 45440 118120 45600
rect 117960 45600 118120 45760
rect 117960 45760 118120 45920
rect 117960 45920 118120 46080
rect 117960 46080 118120 46240
rect 117960 46240 118120 46400
rect 117960 46400 118120 46560
rect 117960 46560 118120 46720
rect 117960 46720 118120 46880
rect 117960 46880 118120 47040
rect 117960 47040 118120 47200
rect 117960 47200 118120 47360
rect 117960 47360 118120 47520
rect 117960 47520 118120 47680
rect 117960 47680 118120 47840
rect 117960 47840 118120 48000
rect 117960 48000 118120 48160
rect 117960 48160 118120 48320
rect 117960 48320 118120 48480
rect 117960 48480 118120 48640
rect 117960 48640 118120 48800
rect 117960 48800 118120 48960
rect 117960 48960 118120 49120
rect 117960 49120 118120 49280
rect 117960 49280 118120 49440
rect 117960 49440 118120 49600
rect 117960 49600 118120 49760
rect 117960 49760 118120 49920
rect 117960 49920 118120 50080
rect 117960 52160 118120 52320
rect 117960 52320 118120 52480
rect 117960 52480 118120 52640
rect 117960 52640 118120 52800
rect 117960 52800 118120 52960
rect 117960 52960 118120 53120
rect 117960 53120 118120 53280
rect 117960 53280 118120 53440
rect 117960 53440 118120 53600
rect 117960 53600 118120 53760
rect 117960 53760 118120 53920
rect 117960 53920 118120 54080
rect 117960 54080 118120 54240
rect 117960 54240 118120 54400
rect 117960 54400 118120 54560
rect 117960 54560 118120 54720
rect 117960 54720 118120 54880
rect 117960 54880 118120 55040
rect 117960 55040 118120 55200
rect 118120 45760 118280 45920
rect 118120 45920 118280 46080
rect 118120 46080 118280 46240
rect 118120 46240 118280 46400
rect 118120 46400 118280 46560
rect 118120 46560 118280 46720
rect 118120 46720 118280 46880
rect 118120 46880 118280 47040
rect 118120 47040 118280 47200
rect 118120 47200 118280 47360
rect 118120 47360 118280 47520
rect 118120 47520 118280 47680
rect 118120 47680 118280 47840
rect 118120 47840 118280 48000
rect 118120 48000 118280 48160
rect 118120 48160 118280 48320
rect 118120 48320 118280 48480
rect 118120 48480 118280 48640
rect 118120 48640 118280 48800
rect 118120 48800 118280 48960
rect 118120 48960 118280 49120
rect 118120 49120 118280 49280
rect 118120 49280 118280 49440
rect 118120 49440 118280 49600
rect 118120 49600 118280 49760
rect 118120 49760 118280 49920
rect 118120 52320 118280 52480
rect 118120 52480 118280 52640
rect 118120 52640 118280 52800
rect 118120 52800 118280 52960
rect 118120 52960 118280 53120
rect 118120 53120 118280 53280
rect 118120 53280 118280 53440
rect 118120 53440 118280 53600
rect 118120 53600 118280 53760
rect 118120 53760 118280 53920
rect 118120 53920 118280 54080
rect 118120 54080 118280 54240
rect 118120 54240 118280 54400
rect 118120 54400 118280 54560
rect 118120 54560 118280 54720
rect 118120 54720 118280 54880
rect 118120 54880 118280 55040
rect 118120 55040 118280 55200
rect 118280 46080 118440 46240
rect 118280 46240 118440 46400
rect 118280 46400 118440 46560
rect 118280 46560 118440 46720
rect 118280 46720 118440 46880
rect 118280 46880 118440 47040
rect 118280 47040 118440 47200
rect 118280 47200 118440 47360
rect 118280 47360 118440 47520
rect 118280 47520 118440 47680
rect 118280 47680 118440 47840
rect 118280 47840 118440 48000
rect 118280 48000 118440 48160
rect 118280 48160 118440 48320
rect 118280 48320 118440 48480
rect 118280 48480 118440 48640
rect 118280 48640 118440 48800
rect 118280 48800 118440 48960
rect 118280 48960 118440 49120
rect 118280 49120 118440 49280
rect 118280 49280 118440 49440
rect 118280 49440 118440 49600
rect 118280 49600 118440 49760
rect 118280 49760 118440 49920
rect 118280 52320 118440 52480
rect 118280 52480 118440 52640
rect 118280 52640 118440 52800
rect 118280 52800 118440 52960
rect 118280 52960 118440 53120
rect 118280 53120 118440 53280
rect 118280 53280 118440 53440
rect 118280 53440 118440 53600
rect 118280 53600 118440 53760
rect 118280 53760 118440 53920
rect 118280 53920 118440 54080
rect 118280 54080 118440 54240
rect 118280 54240 118440 54400
rect 118280 54400 118440 54560
rect 118280 54560 118440 54720
rect 118280 54720 118440 54880
rect 118280 54880 118440 55040
rect 118280 55040 118440 55200
rect 118440 46240 118600 46400
rect 118440 46400 118600 46560
rect 118440 46560 118600 46720
rect 118440 46720 118600 46880
rect 118440 46880 118600 47040
rect 118440 47040 118600 47200
rect 118440 47200 118600 47360
rect 118440 47360 118600 47520
rect 118440 47520 118600 47680
rect 118440 47680 118600 47840
rect 118440 47840 118600 48000
rect 118440 48000 118600 48160
rect 118440 48160 118600 48320
rect 118440 48320 118600 48480
rect 118440 48480 118600 48640
rect 118440 48640 118600 48800
rect 118440 48800 118600 48960
rect 118440 48960 118600 49120
rect 118440 49120 118600 49280
rect 118440 49280 118600 49440
rect 118440 49440 118600 49600
rect 118440 49600 118600 49760
rect 118440 49760 118600 49920
rect 118440 52320 118600 52480
rect 118440 52480 118600 52640
rect 118440 52640 118600 52800
rect 118440 52800 118600 52960
rect 118440 52960 118600 53120
rect 118440 53120 118600 53280
rect 118440 53280 118600 53440
rect 118440 53440 118600 53600
rect 118440 53600 118600 53760
rect 118440 53760 118600 53920
rect 118440 53920 118600 54080
rect 118440 54080 118600 54240
rect 118440 54240 118600 54400
rect 118440 54400 118600 54560
rect 118440 54560 118600 54720
rect 118440 54720 118600 54880
rect 118440 54880 118600 55040
rect 118440 55040 118600 55200
rect 118600 46560 118760 46720
rect 118600 46720 118760 46880
rect 118600 46880 118760 47040
rect 118600 47040 118760 47200
rect 118600 47200 118760 47360
rect 118600 47360 118760 47520
rect 118600 47520 118760 47680
rect 118600 47680 118760 47840
rect 118600 47840 118760 48000
rect 118600 48000 118760 48160
rect 118600 48160 118760 48320
rect 118600 48320 118760 48480
rect 118600 48480 118760 48640
rect 118600 48640 118760 48800
rect 118600 48800 118760 48960
rect 118600 48960 118760 49120
rect 118600 49120 118760 49280
rect 118600 49280 118760 49440
rect 118600 49440 118760 49600
rect 118600 49600 118760 49760
rect 118600 49760 118760 49920
rect 118600 52320 118760 52480
rect 118600 52480 118760 52640
rect 118600 52640 118760 52800
rect 118600 52800 118760 52960
rect 118600 52960 118760 53120
rect 118600 53120 118760 53280
rect 118600 53280 118760 53440
rect 118600 53440 118760 53600
rect 118600 53600 118760 53760
rect 118600 53760 118760 53920
rect 118600 53920 118760 54080
rect 118600 54080 118760 54240
rect 118600 54240 118760 54400
rect 118600 54400 118760 54560
rect 118600 54560 118760 54720
rect 118600 54720 118760 54880
rect 118600 54880 118760 55040
rect 118600 55040 118760 55200
rect 118760 46720 118920 46880
rect 118760 46880 118920 47040
rect 118760 47040 118920 47200
rect 118760 47200 118920 47360
rect 118760 47360 118920 47520
rect 118760 47520 118920 47680
rect 118760 47680 118920 47840
rect 118760 47840 118920 48000
rect 118760 48000 118920 48160
rect 118760 48160 118920 48320
rect 118760 48320 118920 48480
rect 118760 48480 118920 48640
rect 118760 48640 118920 48800
rect 118760 48800 118920 48960
rect 118760 48960 118920 49120
rect 118760 49120 118920 49280
rect 118760 49280 118920 49440
rect 118760 49440 118920 49600
rect 118760 49600 118920 49760
rect 118760 49760 118920 49920
rect 118760 52320 118920 52480
rect 118760 52480 118920 52640
rect 118760 52640 118920 52800
rect 118760 52800 118920 52960
rect 118760 52960 118920 53120
rect 118760 53120 118920 53280
rect 118760 53280 118920 53440
rect 118760 53440 118920 53600
rect 118760 53600 118920 53760
rect 118760 53760 118920 53920
rect 118760 53920 118920 54080
rect 118760 54080 118920 54240
rect 118760 54240 118920 54400
rect 118760 54400 118920 54560
rect 118760 54560 118920 54720
rect 118760 54720 118920 54880
rect 118760 54880 118920 55040
rect 118920 47040 119080 47200
rect 118920 47200 119080 47360
rect 118920 47360 119080 47520
rect 118920 47520 119080 47680
rect 118920 47680 119080 47840
rect 118920 47840 119080 48000
rect 118920 48000 119080 48160
rect 118920 48160 119080 48320
rect 118920 48320 119080 48480
rect 118920 48480 119080 48640
rect 118920 48640 119080 48800
rect 118920 48800 119080 48960
rect 118920 48960 119080 49120
rect 118920 49120 119080 49280
rect 118920 49280 119080 49440
rect 118920 49440 119080 49600
rect 118920 49600 119080 49760
rect 118920 49760 119080 49920
rect 118920 49920 119080 50080
rect 118920 52320 119080 52480
rect 118920 52480 119080 52640
rect 118920 52640 119080 52800
rect 118920 52800 119080 52960
rect 118920 52960 119080 53120
rect 118920 53120 119080 53280
rect 118920 53280 119080 53440
rect 118920 53440 119080 53600
rect 118920 53600 119080 53760
rect 118920 53760 119080 53920
rect 118920 53920 119080 54080
rect 118920 54080 119080 54240
rect 118920 54240 119080 54400
rect 118920 54400 119080 54560
rect 118920 54560 119080 54720
rect 118920 54720 119080 54880
rect 118920 54880 119080 55040
rect 119080 47200 119240 47360
rect 119080 47360 119240 47520
rect 119080 47520 119240 47680
rect 119080 47680 119240 47840
rect 119080 47840 119240 48000
rect 119080 48000 119240 48160
rect 119080 48160 119240 48320
rect 119080 48320 119240 48480
rect 119080 48480 119240 48640
rect 119080 48640 119240 48800
rect 119080 48800 119240 48960
rect 119080 48960 119240 49120
rect 119080 49120 119240 49280
rect 119080 49280 119240 49440
rect 119080 49440 119240 49600
rect 119080 49600 119240 49760
rect 119080 49760 119240 49920
rect 119080 49920 119240 50080
rect 119080 52320 119240 52480
rect 119080 52480 119240 52640
rect 119080 52640 119240 52800
rect 119080 52800 119240 52960
rect 119080 52960 119240 53120
rect 119080 53120 119240 53280
rect 119080 53280 119240 53440
rect 119080 53440 119240 53600
rect 119080 53600 119240 53760
rect 119080 53760 119240 53920
rect 119080 53920 119240 54080
rect 119080 54080 119240 54240
rect 119080 54240 119240 54400
rect 119080 54400 119240 54560
rect 119080 54560 119240 54720
rect 119080 54720 119240 54880
rect 119080 54880 119240 55040
rect 119240 47200 119400 47360
rect 119240 47360 119400 47520
rect 119240 47520 119400 47680
rect 119240 47680 119400 47840
rect 119240 47840 119400 48000
rect 119240 48000 119400 48160
rect 119240 48160 119400 48320
rect 119240 48320 119400 48480
rect 119240 48480 119400 48640
rect 119240 48640 119400 48800
rect 119240 48800 119400 48960
rect 119240 48960 119400 49120
rect 119240 49120 119400 49280
rect 119240 49280 119400 49440
rect 119240 49440 119400 49600
rect 119240 49600 119400 49760
rect 119240 49760 119400 49920
rect 119240 49920 119400 50080
rect 119240 50080 119400 50240
rect 119240 52160 119400 52320
rect 119240 52320 119400 52480
rect 119240 52480 119400 52640
rect 119240 52640 119400 52800
rect 119240 52800 119400 52960
rect 119240 52960 119400 53120
rect 119240 53120 119400 53280
rect 119240 53280 119400 53440
rect 119240 53440 119400 53600
rect 119240 53600 119400 53760
rect 119240 53760 119400 53920
rect 119240 53920 119400 54080
rect 119240 54080 119400 54240
rect 119240 54240 119400 54400
rect 119240 54400 119400 54560
rect 119240 54560 119400 54720
rect 119240 54720 119400 54880
rect 119240 54880 119400 55040
rect 119400 47360 119560 47520
rect 119400 47520 119560 47680
rect 119400 47680 119560 47840
rect 119400 47840 119560 48000
rect 119400 48000 119560 48160
rect 119400 48160 119560 48320
rect 119400 48320 119560 48480
rect 119400 48480 119560 48640
rect 119400 48640 119560 48800
rect 119400 48800 119560 48960
rect 119400 48960 119560 49120
rect 119400 49120 119560 49280
rect 119400 49280 119560 49440
rect 119400 49440 119560 49600
rect 119400 49600 119560 49760
rect 119400 49760 119560 49920
rect 119400 49920 119560 50080
rect 119400 50080 119560 50240
rect 119400 50240 119560 50400
rect 119400 52000 119560 52160
rect 119400 52160 119560 52320
rect 119400 52320 119560 52480
rect 119400 52480 119560 52640
rect 119400 52640 119560 52800
rect 119400 52800 119560 52960
rect 119400 52960 119560 53120
rect 119400 53120 119560 53280
rect 119400 53280 119560 53440
rect 119400 53440 119560 53600
rect 119400 53600 119560 53760
rect 119400 53760 119560 53920
rect 119400 53920 119560 54080
rect 119400 54080 119560 54240
rect 119400 54240 119560 54400
rect 119400 54400 119560 54560
rect 119400 54560 119560 54720
rect 119400 54720 119560 54880
rect 119400 54880 119560 55040
rect 119560 47520 119720 47680
rect 119560 47680 119720 47840
rect 119560 47840 119720 48000
rect 119560 48000 119720 48160
rect 119560 48160 119720 48320
rect 119560 48320 119720 48480
rect 119560 48480 119720 48640
rect 119560 48640 119720 48800
rect 119560 48800 119720 48960
rect 119560 48960 119720 49120
rect 119560 49120 119720 49280
rect 119560 49280 119720 49440
rect 119560 49440 119720 49600
rect 119560 49600 119720 49760
rect 119560 49760 119720 49920
rect 119560 49920 119720 50080
rect 119560 50080 119720 50240
rect 119560 50240 119720 50400
rect 119560 50400 119720 50560
rect 119560 50560 119720 50720
rect 119560 51520 119720 51680
rect 119560 51680 119720 51840
rect 119560 51840 119720 52000
rect 119560 52000 119720 52160
rect 119560 52160 119720 52320
rect 119560 52320 119720 52480
rect 119560 52480 119720 52640
rect 119560 52640 119720 52800
rect 119560 52800 119720 52960
rect 119560 52960 119720 53120
rect 119560 53120 119720 53280
rect 119560 53280 119720 53440
rect 119560 53440 119720 53600
rect 119560 53600 119720 53760
rect 119560 53760 119720 53920
rect 119560 53920 119720 54080
rect 119560 54080 119720 54240
rect 119560 54240 119720 54400
rect 119560 54400 119720 54560
rect 119560 54560 119720 54720
rect 119560 54720 119720 54880
rect 119720 47520 119880 47680
rect 119720 47680 119880 47840
rect 119720 47840 119880 48000
rect 119720 48000 119880 48160
rect 119720 48160 119880 48320
rect 119720 48320 119880 48480
rect 119720 48480 119880 48640
rect 119720 48640 119880 48800
rect 119720 48800 119880 48960
rect 119720 48960 119880 49120
rect 119720 49120 119880 49280
rect 119720 49280 119880 49440
rect 119720 49440 119880 49600
rect 119720 49600 119880 49760
rect 119720 49760 119880 49920
rect 119720 49920 119880 50080
rect 119720 50080 119880 50240
rect 119720 50240 119880 50400
rect 119720 50400 119880 50560
rect 119720 50560 119880 50720
rect 119720 50720 119880 50880
rect 119720 50880 119880 51040
rect 119720 51040 119880 51200
rect 119720 51200 119880 51360
rect 119720 51360 119880 51520
rect 119720 51520 119880 51680
rect 119720 51680 119880 51840
rect 119720 51840 119880 52000
rect 119720 52000 119880 52160
rect 119720 52160 119880 52320
rect 119720 52320 119880 52480
rect 119720 52480 119880 52640
rect 119720 52640 119880 52800
rect 119720 52800 119880 52960
rect 119720 52960 119880 53120
rect 119720 53120 119880 53280
rect 119720 53280 119880 53440
rect 119720 53440 119880 53600
rect 119720 53600 119880 53760
rect 119720 53760 119880 53920
rect 119720 53920 119880 54080
rect 119720 54080 119880 54240
rect 119720 54240 119880 54400
rect 119720 54400 119880 54560
rect 119720 54560 119880 54720
rect 119720 54720 119880 54880
rect 119880 47680 120040 47840
rect 119880 47840 120040 48000
rect 119880 48000 120040 48160
rect 119880 48160 120040 48320
rect 119880 48320 120040 48480
rect 119880 48480 120040 48640
rect 119880 48640 120040 48800
rect 119880 48800 120040 48960
rect 119880 48960 120040 49120
rect 119880 49120 120040 49280
rect 119880 49280 120040 49440
rect 119880 49440 120040 49600
rect 119880 49600 120040 49760
rect 119880 49760 120040 49920
rect 119880 49920 120040 50080
rect 119880 50080 120040 50240
rect 119880 50240 120040 50400
rect 119880 50400 120040 50560
rect 119880 50560 120040 50720
rect 119880 50720 120040 50880
rect 119880 50880 120040 51040
rect 119880 51040 120040 51200
rect 119880 51200 120040 51360
rect 119880 51360 120040 51520
rect 119880 51520 120040 51680
rect 119880 51680 120040 51840
rect 119880 51840 120040 52000
rect 119880 52000 120040 52160
rect 119880 52160 120040 52320
rect 119880 52320 120040 52480
rect 119880 52480 120040 52640
rect 119880 52640 120040 52800
rect 119880 52800 120040 52960
rect 119880 52960 120040 53120
rect 119880 53120 120040 53280
rect 119880 53280 120040 53440
rect 119880 53440 120040 53600
rect 119880 53600 120040 53760
rect 119880 53760 120040 53920
rect 119880 53920 120040 54080
rect 119880 54080 120040 54240
rect 119880 54240 120040 54400
rect 119880 54400 120040 54560
rect 119880 54560 120040 54720
rect 120040 47680 120200 47840
rect 120040 47840 120200 48000
rect 120040 48000 120200 48160
rect 120040 48160 120200 48320
rect 120040 48320 120200 48480
rect 120040 48480 120200 48640
rect 120040 48640 120200 48800
rect 120040 48800 120200 48960
rect 120040 48960 120200 49120
rect 120040 49120 120200 49280
rect 120040 49280 120200 49440
rect 120040 49440 120200 49600
rect 120040 49600 120200 49760
rect 120040 49760 120200 49920
rect 120040 49920 120200 50080
rect 120040 50080 120200 50240
rect 120040 50240 120200 50400
rect 120040 50400 120200 50560
rect 120040 50560 120200 50720
rect 120040 50720 120200 50880
rect 120040 50880 120200 51040
rect 120040 51040 120200 51200
rect 120040 51200 120200 51360
rect 120040 51360 120200 51520
rect 120040 51520 120200 51680
rect 120040 51680 120200 51840
rect 120040 51840 120200 52000
rect 120040 52000 120200 52160
rect 120040 52160 120200 52320
rect 120040 52320 120200 52480
rect 120040 52480 120200 52640
rect 120040 52640 120200 52800
rect 120040 52800 120200 52960
rect 120040 52960 120200 53120
rect 120040 53120 120200 53280
rect 120040 53280 120200 53440
rect 120040 53440 120200 53600
rect 120040 53600 120200 53760
rect 120040 53760 120200 53920
rect 120040 53920 120200 54080
rect 120040 54080 120200 54240
rect 120040 54240 120200 54400
rect 120040 54400 120200 54560
rect 120040 54560 120200 54720
rect 120200 47840 120360 48000
rect 120200 48000 120360 48160
rect 120200 48160 120360 48320
rect 120200 48320 120360 48480
rect 120200 48480 120360 48640
rect 120200 48640 120360 48800
rect 120200 48800 120360 48960
rect 120200 48960 120360 49120
rect 120200 49120 120360 49280
rect 120200 49280 120360 49440
rect 120200 49440 120360 49600
rect 120200 49600 120360 49760
rect 120200 49760 120360 49920
rect 120200 49920 120360 50080
rect 120200 50080 120360 50240
rect 120200 50240 120360 50400
rect 120200 50400 120360 50560
rect 120200 50560 120360 50720
rect 120200 50720 120360 50880
rect 120200 50880 120360 51040
rect 120200 51040 120360 51200
rect 120200 51200 120360 51360
rect 120200 51360 120360 51520
rect 120200 51520 120360 51680
rect 120200 51680 120360 51840
rect 120200 51840 120360 52000
rect 120200 52000 120360 52160
rect 120200 52160 120360 52320
rect 120200 52320 120360 52480
rect 120200 52480 120360 52640
rect 120200 52640 120360 52800
rect 120200 52800 120360 52960
rect 120200 52960 120360 53120
rect 120200 53120 120360 53280
rect 120200 53280 120360 53440
rect 120200 53440 120360 53600
rect 120200 53600 120360 53760
rect 120200 53760 120360 53920
rect 120200 53920 120360 54080
rect 120200 54080 120360 54240
rect 120200 54240 120360 54400
rect 120200 54400 120360 54560
rect 120360 47840 120520 48000
rect 120360 48000 120520 48160
rect 120360 48160 120520 48320
rect 120360 48320 120520 48480
rect 120360 48480 120520 48640
rect 120360 48640 120520 48800
rect 120360 48800 120520 48960
rect 120360 48960 120520 49120
rect 120360 49120 120520 49280
rect 120360 49280 120520 49440
rect 120360 49440 120520 49600
rect 120360 49600 120520 49760
rect 120360 49760 120520 49920
rect 120360 49920 120520 50080
rect 120360 50080 120520 50240
rect 120360 50240 120520 50400
rect 120360 50400 120520 50560
rect 120360 50560 120520 50720
rect 120360 50720 120520 50880
rect 120360 50880 120520 51040
rect 120360 51040 120520 51200
rect 120360 51200 120520 51360
rect 120360 51360 120520 51520
rect 120360 51520 120520 51680
rect 120360 51680 120520 51840
rect 120360 51840 120520 52000
rect 120360 52000 120520 52160
rect 120360 52160 120520 52320
rect 120360 52320 120520 52480
rect 120360 52480 120520 52640
rect 120360 52640 120520 52800
rect 120360 52800 120520 52960
rect 120360 52960 120520 53120
rect 120360 53120 120520 53280
rect 120360 53280 120520 53440
rect 120360 53440 120520 53600
rect 120360 53600 120520 53760
rect 120360 53760 120520 53920
rect 120360 53920 120520 54080
rect 120360 54080 120520 54240
rect 120360 54240 120520 54400
rect 120360 54400 120520 54560
rect 120520 48000 120680 48160
rect 120520 48160 120680 48320
rect 120520 48320 120680 48480
rect 120520 48480 120680 48640
rect 120520 48640 120680 48800
rect 120520 48800 120680 48960
rect 120520 48960 120680 49120
rect 120520 49120 120680 49280
rect 120520 49280 120680 49440
rect 120520 49440 120680 49600
rect 120520 49600 120680 49760
rect 120520 49760 120680 49920
rect 120520 49920 120680 50080
rect 120520 50080 120680 50240
rect 120520 50240 120680 50400
rect 120520 50400 120680 50560
rect 120520 50560 120680 50720
rect 120520 50720 120680 50880
rect 120520 50880 120680 51040
rect 120520 51040 120680 51200
rect 120520 51200 120680 51360
rect 120520 51360 120680 51520
rect 120520 51520 120680 51680
rect 120520 51680 120680 51840
rect 120520 51840 120680 52000
rect 120520 52000 120680 52160
rect 120520 52160 120680 52320
rect 120520 52320 120680 52480
rect 120520 52480 120680 52640
rect 120520 52640 120680 52800
rect 120520 52800 120680 52960
rect 120520 52960 120680 53120
rect 120520 53120 120680 53280
rect 120520 53280 120680 53440
rect 120520 53440 120680 53600
rect 120520 53600 120680 53760
rect 120520 53760 120680 53920
rect 120520 53920 120680 54080
rect 120520 54080 120680 54240
rect 120520 54240 120680 54400
rect 120680 48160 120840 48320
rect 120680 48320 120840 48480
rect 120680 48480 120840 48640
rect 120680 48640 120840 48800
rect 120680 48800 120840 48960
rect 120680 48960 120840 49120
rect 120680 49120 120840 49280
rect 120680 49280 120840 49440
rect 120680 49440 120840 49600
rect 120680 49600 120840 49760
rect 120680 49760 120840 49920
rect 120680 49920 120840 50080
rect 120680 50080 120840 50240
rect 120680 50240 120840 50400
rect 120680 50400 120840 50560
rect 120680 50560 120840 50720
rect 120680 50720 120840 50880
rect 120680 50880 120840 51040
rect 120680 51040 120840 51200
rect 120680 51200 120840 51360
rect 120680 51360 120840 51520
rect 120680 51520 120840 51680
rect 120680 51680 120840 51840
rect 120680 51840 120840 52000
rect 120680 52000 120840 52160
rect 120680 52160 120840 52320
rect 120680 52320 120840 52480
rect 120680 52480 120840 52640
rect 120680 52640 120840 52800
rect 120680 52800 120840 52960
rect 120680 52960 120840 53120
rect 120680 53120 120840 53280
rect 120680 53280 120840 53440
rect 120680 53440 120840 53600
rect 120680 53600 120840 53760
rect 120680 53760 120840 53920
rect 120680 53920 120840 54080
rect 120680 54080 120840 54240
rect 120680 54240 120840 54400
rect 120840 48320 121000 48480
rect 120840 48480 121000 48640
rect 120840 48640 121000 48800
rect 120840 48800 121000 48960
rect 120840 48960 121000 49120
rect 120840 49120 121000 49280
rect 120840 49280 121000 49440
rect 120840 49440 121000 49600
rect 120840 49600 121000 49760
rect 120840 49760 121000 49920
rect 120840 49920 121000 50080
rect 120840 50080 121000 50240
rect 120840 50240 121000 50400
rect 120840 50400 121000 50560
rect 120840 50560 121000 50720
rect 120840 50720 121000 50880
rect 120840 50880 121000 51040
rect 120840 51040 121000 51200
rect 120840 51200 121000 51360
rect 120840 51360 121000 51520
rect 120840 51520 121000 51680
rect 120840 51680 121000 51840
rect 120840 51840 121000 52000
rect 120840 52000 121000 52160
rect 120840 52160 121000 52320
rect 120840 52320 121000 52480
rect 120840 52480 121000 52640
rect 120840 52640 121000 52800
rect 120840 52800 121000 52960
rect 120840 52960 121000 53120
rect 120840 53120 121000 53280
rect 120840 53280 121000 53440
rect 120840 53440 121000 53600
rect 120840 53600 121000 53760
rect 120840 53760 121000 53920
rect 120840 53920 121000 54080
rect 120840 54080 121000 54240
rect 121000 48320 121160 48480
rect 121000 48480 121160 48640
rect 121000 48640 121160 48800
rect 121000 48800 121160 48960
rect 121000 48960 121160 49120
rect 121000 49120 121160 49280
rect 121000 49280 121160 49440
rect 121000 49440 121160 49600
rect 121000 49600 121160 49760
rect 121000 49760 121160 49920
rect 121000 49920 121160 50080
rect 121000 50080 121160 50240
rect 121000 50240 121160 50400
rect 121000 50400 121160 50560
rect 121000 50560 121160 50720
rect 121000 50720 121160 50880
rect 121000 50880 121160 51040
rect 121000 51040 121160 51200
rect 121000 51200 121160 51360
rect 121000 51360 121160 51520
rect 121000 51520 121160 51680
rect 121000 51680 121160 51840
rect 121000 51840 121160 52000
rect 121000 52000 121160 52160
rect 121000 52160 121160 52320
rect 121000 52320 121160 52480
rect 121000 52480 121160 52640
rect 121000 52640 121160 52800
rect 121000 52800 121160 52960
rect 121000 52960 121160 53120
rect 121000 53120 121160 53280
rect 121000 53280 121160 53440
rect 121000 53440 121160 53600
rect 121000 53600 121160 53760
rect 121000 53760 121160 53920
rect 121000 53920 121160 54080
rect 121160 48480 121320 48640
rect 121160 48640 121320 48800
rect 121160 48800 121320 48960
rect 121160 48960 121320 49120
rect 121160 49120 121320 49280
rect 121160 49280 121320 49440
rect 121160 49440 121320 49600
rect 121160 49600 121320 49760
rect 121160 49760 121320 49920
rect 121160 49920 121320 50080
rect 121160 50080 121320 50240
rect 121160 50240 121320 50400
rect 121160 50400 121320 50560
rect 121160 50560 121320 50720
rect 121160 50720 121320 50880
rect 121160 50880 121320 51040
rect 121160 51040 121320 51200
rect 121160 51200 121320 51360
rect 121160 51360 121320 51520
rect 121160 51520 121320 51680
rect 121160 51680 121320 51840
rect 121160 51840 121320 52000
rect 121160 52000 121320 52160
rect 121160 52160 121320 52320
rect 121160 52320 121320 52480
rect 121160 52480 121320 52640
rect 121160 52640 121320 52800
rect 121160 52800 121320 52960
rect 121160 52960 121320 53120
rect 121160 53120 121320 53280
rect 121160 53280 121320 53440
rect 121160 53440 121320 53600
rect 121160 53600 121320 53760
rect 121160 53760 121320 53920
rect 121320 48640 121480 48800
rect 121320 48800 121480 48960
rect 121320 48960 121480 49120
rect 121320 49120 121480 49280
rect 121320 49280 121480 49440
rect 121320 49440 121480 49600
rect 121320 49600 121480 49760
rect 121320 49760 121480 49920
rect 121320 49920 121480 50080
rect 121320 50080 121480 50240
rect 121320 50240 121480 50400
rect 121320 50400 121480 50560
rect 121320 50560 121480 50720
rect 121320 50720 121480 50880
rect 121320 50880 121480 51040
rect 121320 51040 121480 51200
rect 121320 51200 121480 51360
rect 121320 51360 121480 51520
rect 121320 51520 121480 51680
rect 121320 51680 121480 51840
rect 121320 51840 121480 52000
rect 121320 52000 121480 52160
rect 121320 52160 121480 52320
rect 121320 52320 121480 52480
rect 121320 52480 121480 52640
rect 121320 52640 121480 52800
rect 121320 52800 121480 52960
rect 121320 52960 121480 53120
rect 121320 53120 121480 53280
rect 121320 53280 121480 53440
rect 121320 53440 121480 53600
rect 121320 53600 121480 53760
rect 121480 48800 121640 48960
rect 121480 48960 121640 49120
rect 121480 49120 121640 49280
rect 121480 49280 121640 49440
rect 121480 49440 121640 49600
rect 121480 49600 121640 49760
rect 121480 49760 121640 49920
rect 121480 49920 121640 50080
rect 121480 50080 121640 50240
rect 121480 50240 121640 50400
rect 121480 50400 121640 50560
rect 121480 50560 121640 50720
rect 121480 50720 121640 50880
rect 121480 50880 121640 51040
rect 121480 51040 121640 51200
rect 121480 51200 121640 51360
rect 121480 51360 121640 51520
rect 121480 51520 121640 51680
rect 121480 51680 121640 51840
rect 121480 51840 121640 52000
rect 121480 52000 121640 52160
rect 121480 52160 121640 52320
rect 121480 52320 121640 52480
rect 121480 52480 121640 52640
rect 121480 52640 121640 52800
rect 121480 52800 121640 52960
rect 121480 52960 121640 53120
rect 121480 53120 121640 53280
rect 121480 53280 121640 53440
rect 121640 48960 121800 49120
rect 121640 49120 121800 49280
rect 121640 49280 121800 49440
rect 121640 49440 121800 49600
rect 121640 49600 121800 49760
rect 121640 49760 121800 49920
rect 121640 49920 121800 50080
rect 121640 50080 121800 50240
rect 121640 50240 121800 50400
rect 121640 50400 121800 50560
rect 121640 50560 121800 50720
rect 121640 50720 121800 50880
rect 121640 50880 121800 51040
rect 121640 51040 121800 51200
rect 121640 51200 121800 51360
rect 121640 51360 121800 51520
rect 121640 51520 121800 51680
rect 121640 51680 121800 51840
rect 121640 51840 121800 52000
rect 121640 52000 121800 52160
rect 121640 52160 121800 52320
rect 121640 52320 121800 52480
rect 121640 52480 121800 52640
rect 121640 52640 121800 52800
rect 121640 52800 121800 52960
rect 121640 52960 121800 53120
rect 121640 53120 121800 53280
rect 121800 49120 121960 49280
rect 121800 49280 121960 49440
rect 121800 49440 121960 49600
rect 121800 49600 121960 49760
rect 121800 49760 121960 49920
rect 121800 49920 121960 50080
rect 121800 50080 121960 50240
rect 121800 50240 121960 50400
rect 121800 50400 121960 50560
rect 121800 50560 121960 50720
rect 121800 50720 121960 50880
rect 121800 50880 121960 51040
rect 121800 51040 121960 51200
rect 121800 51200 121960 51360
rect 121800 51360 121960 51520
rect 121800 51520 121960 51680
rect 121800 51680 121960 51840
rect 121800 51840 121960 52000
rect 121800 52000 121960 52160
rect 121800 52160 121960 52320
rect 121800 52320 121960 52480
rect 121800 52480 121960 52640
rect 121800 52640 121960 52800
rect 121960 49280 122120 49440
rect 121960 49440 122120 49600
rect 121960 49600 122120 49760
rect 121960 49760 122120 49920
rect 121960 49920 122120 50080
rect 121960 50080 122120 50240
rect 121960 50240 122120 50400
rect 121960 50400 122120 50560
rect 121960 50560 122120 50720
rect 121960 50720 122120 50880
rect 121960 50880 122120 51040
rect 121960 51040 122120 51200
rect 121960 51200 122120 51360
rect 121960 51360 122120 51520
rect 121960 51520 122120 51680
rect 121960 51680 122120 51840
rect 121960 51840 122120 52000
rect 121960 52000 122120 52160
rect 121960 52160 122120 52320
rect 121960 52320 122120 52480
rect 122120 49440 122280 49600
rect 122120 49600 122280 49760
rect 122120 49760 122280 49920
rect 122120 49920 122280 50080
rect 122120 50080 122280 50240
rect 122120 50240 122280 50400
rect 122120 50400 122280 50560
rect 122120 50560 122280 50720
rect 122120 50720 122280 50880
rect 122120 50880 122280 51040
rect 122120 51040 122280 51200
rect 122120 51200 122280 51360
rect 122120 51360 122280 51520
rect 122120 51520 122280 51680
rect 122120 51680 122280 51840
rect 122120 51840 122280 52000
rect 122280 49600 122440 49760
rect 122280 49760 122440 49920
rect 122280 49920 122440 50080
rect 122280 50080 122440 50240
rect 122280 50240 122440 50400
rect 122280 50400 122440 50560
rect 122280 50560 122440 50720
rect 122280 50720 122440 50880
rect 122280 50880 122440 51040
rect 122280 51040 122440 51200
rect 122280 51200 122440 51360
rect 122280 51360 122440 51520
rect 122440 36320 122600 36480
rect 122440 36480 122600 36640
rect 122440 36640 122600 36800
rect 122440 36800 122600 36960
rect 122440 36960 122600 37120
rect 122440 37120 122600 37280
rect 122440 37280 122600 37440
rect 122440 37440 122600 37600
rect 122440 37600 122600 37760
rect 122440 37760 122600 37920
rect 122440 37920 122600 38080
rect 122440 38080 122600 38240
rect 122440 38240 122600 38400
rect 122440 38400 122600 38560
rect 122440 38560 122600 38720
rect 122440 38720 122600 38880
rect 122440 38880 122600 39040
rect 122440 39040 122600 39200
rect 122440 39200 122600 39360
rect 122440 39360 122600 39520
rect 122440 39520 122600 39680
rect 122440 39680 122600 39840
rect 122440 40000 122600 40160
rect 122440 50080 122600 50240
rect 122440 50240 122600 50400
rect 122440 50400 122600 50560
rect 122440 50560 122600 50720
rect 122440 50720 122600 50880
rect 122600 35040 122760 35200
rect 122600 35200 122760 35360
rect 122600 35360 122760 35520
rect 122600 35520 122760 35680
rect 122600 35680 122760 35840
rect 122600 35840 122760 36000
rect 122600 36000 122760 36160
rect 122600 36160 122760 36320
rect 122600 36320 122760 36480
rect 122600 36480 122760 36640
rect 122600 36640 122760 36800
rect 122600 36800 122760 36960
rect 122600 36960 122760 37120
rect 122600 37120 122760 37280
rect 122600 37280 122760 37440
rect 122600 37440 122760 37600
rect 122600 37600 122760 37760
rect 122600 37760 122760 37920
rect 122600 37920 122760 38080
rect 122600 38080 122760 38240
rect 122600 38240 122760 38400
rect 122600 38400 122760 38560
rect 122600 38560 122760 38720
rect 122600 38720 122760 38880
rect 122600 38880 122760 39040
rect 122600 39040 122760 39200
rect 122600 39200 122760 39360
rect 122600 39360 122760 39520
rect 122600 39520 122760 39680
rect 122600 39680 122760 39840
rect 122600 39840 122760 40000
rect 122600 40000 122760 40160
rect 122600 40160 122760 40320
rect 122600 40320 122760 40480
rect 122600 40480 122760 40640
rect 122600 40640 122760 40800
rect 122600 40800 122760 40960
rect 122600 40960 122760 41120
rect 122600 41120 122760 41280
rect 122760 34400 122920 34560
rect 122760 34560 122920 34720
rect 122760 34720 122920 34880
rect 122760 34880 122920 35040
rect 122760 35040 122920 35200
rect 122760 35200 122920 35360
rect 122760 35360 122920 35520
rect 122760 35520 122920 35680
rect 122760 35680 122920 35840
rect 122760 35840 122920 36000
rect 122760 36000 122920 36160
rect 122760 36160 122920 36320
rect 122760 36320 122920 36480
rect 122760 36480 122920 36640
rect 122760 36640 122920 36800
rect 122760 36800 122920 36960
rect 122760 36960 122920 37120
rect 122760 37120 122920 37280
rect 122760 37280 122920 37440
rect 122760 37440 122920 37600
rect 122760 37600 122920 37760
rect 122760 37760 122920 37920
rect 122760 37920 122920 38080
rect 122760 38080 122920 38240
rect 122760 38240 122920 38400
rect 122760 38400 122920 38560
rect 122760 38560 122920 38720
rect 122760 38720 122920 38880
rect 122760 38880 122920 39040
rect 122760 39040 122920 39200
rect 122760 39200 122920 39360
rect 122760 39360 122920 39520
rect 122760 39520 122920 39680
rect 122760 39680 122920 39840
rect 122760 39840 122920 40000
rect 122760 40000 122920 40160
rect 122760 40160 122920 40320
rect 122760 40320 122920 40480
rect 122760 40480 122920 40640
rect 122760 40640 122920 40800
rect 122760 40800 122920 40960
rect 122760 40960 122920 41120
rect 122760 41120 122920 41280
rect 122760 41280 122920 41440
rect 122760 41440 122920 41600
rect 122760 41600 122920 41760
rect 122760 41760 122920 41920
rect 122760 41920 122920 42080
rect 122920 33760 123080 33920
rect 122920 33920 123080 34080
rect 122920 34080 123080 34240
rect 122920 34240 123080 34400
rect 122920 34400 123080 34560
rect 122920 34560 123080 34720
rect 122920 34720 123080 34880
rect 122920 34880 123080 35040
rect 122920 35040 123080 35200
rect 122920 35200 123080 35360
rect 122920 35360 123080 35520
rect 122920 35520 123080 35680
rect 122920 35680 123080 35840
rect 122920 35840 123080 36000
rect 122920 36000 123080 36160
rect 122920 36160 123080 36320
rect 122920 36320 123080 36480
rect 122920 36480 123080 36640
rect 122920 36640 123080 36800
rect 122920 36800 123080 36960
rect 122920 36960 123080 37120
rect 122920 37120 123080 37280
rect 122920 37280 123080 37440
rect 122920 37440 123080 37600
rect 122920 37600 123080 37760
rect 122920 37760 123080 37920
rect 122920 37920 123080 38080
rect 122920 38080 123080 38240
rect 122920 38240 123080 38400
rect 122920 38400 123080 38560
rect 122920 38560 123080 38720
rect 122920 38720 123080 38880
rect 122920 38880 123080 39040
rect 122920 39040 123080 39200
rect 122920 39200 123080 39360
rect 122920 39360 123080 39520
rect 122920 39520 123080 39680
rect 122920 39680 123080 39840
rect 122920 39840 123080 40000
rect 122920 40000 123080 40160
rect 122920 40160 123080 40320
rect 122920 40320 123080 40480
rect 122920 40480 123080 40640
rect 122920 40640 123080 40800
rect 122920 40800 123080 40960
rect 122920 40960 123080 41120
rect 122920 41120 123080 41280
rect 122920 41280 123080 41440
rect 122920 41440 123080 41600
rect 122920 41600 123080 41760
rect 122920 41760 123080 41920
rect 122920 41920 123080 42080
rect 122920 42080 123080 42240
rect 122920 42240 123080 42400
rect 122920 42400 123080 42560
rect 122920 42560 123080 42720
rect 123080 33280 123240 33440
rect 123080 33440 123240 33600
rect 123080 33600 123240 33760
rect 123080 33760 123240 33920
rect 123080 33920 123240 34080
rect 123080 34080 123240 34240
rect 123080 34240 123240 34400
rect 123080 34400 123240 34560
rect 123080 34560 123240 34720
rect 123080 34720 123240 34880
rect 123080 34880 123240 35040
rect 123080 35040 123240 35200
rect 123080 35200 123240 35360
rect 123080 35360 123240 35520
rect 123080 35520 123240 35680
rect 123080 35680 123240 35840
rect 123080 35840 123240 36000
rect 123080 36000 123240 36160
rect 123080 36160 123240 36320
rect 123080 36320 123240 36480
rect 123080 36480 123240 36640
rect 123080 36640 123240 36800
rect 123080 36800 123240 36960
rect 123080 36960 123240 37120
rect 123080 37120 123240 37280
rect 123080 37280 123240 37440
rect 123080 37440 123240 37600
rect 123080 37600 123240 37760
rect 123080 37760 123240 37920
rect 123080 37920 123240 38080
rect 123080 38080 123240 38240
rect 123080 38240 123240 38400
rect 123080 38400 123240 38560
rect 123080 38560 123240 38720
rect 123080 38720 123240 38880
rect 123080 38880 123240 39040
rect 123080 39040 123240 39200
rect 123080 39200 123240 39360
rect 123080 39360 123240 39520
rect 123080 39520 123240 39680
rect 123080 39680 123240 39840
rect 123080 39840 123240 40000
rect 123080 40000 123240 40160
rect 123080 40160 123240 40320
rect 123080 40320 123240 40480
rect 123080 40480 123240 40640
rect 123080 40640 123240 40800
rect 123080 40800 123240 40960
rect 123080 40960 123240 41120
rect 123080 41120 123240 41280
rect 123080 41280 123240 41440
rect 123080 41440 123240 41600
rect 123080 41600 123240 41760
rect 123080 41760 123240 41920
rect 123080 41920 123240 42080
rect 123080 42080 123240 42240
rect 123080 42240 123240 42400
rect 123080 42400 123240 42560
rect 123080 42560 123240 42720
rect 123080 42720 123240 42880
rect 123080 42880 123240 43040
rect 123080 43040 123240 43200
rect 123080 43200 123240 43360
rect 123240 32800 123400 32960
rect 123240 32960 123400 33120
rect 123240 33120 123400 33280
rect 123240 33280 123400 33440
rect 123240 33440 123400 33600
rect 123240 33600 123400 33760
rect 123240 33760 123400 33920
rect 123240 33920 123400 34080
rect 123240 34080 123400 34240
rect 123240 34240 123400 34400
rect 123240 34400 123400 34560
rect 123240 34560 123400 34720
rect 123240 34720 123400 34880
rect 123240 34880 123400 35040
rect 123240 35040 123400 35200
rect 123240 35200 123400 35360
rect 123240 35360 123400 35520
rect 123240 35520 123400 35680
rect 123240 35680 123400 35840
rect 123240 35840 123400 36000
rect 123240 36000 123400 36160
rect 123240 36160 123400 36320
rect 123240 36320 123400 36480
rect 123240 36480 123400 36640
rect 123240 36640 123400 36800
rect 123240 36800 123400 36960
rect 123240 36960 123400 37120
rect 123240 37120 123400 37280
rect 123240 37280 123400 37440
rect 123240 37440 123400 37600
rect 123240 37600 123400 37760
rect 123240 37760 123400 37920
rect 123240 37920 123400 38080
rect 123240 38080 123400 38240
rect 123240 38240 123400 38400
rect 123240 38400 123400 38560
rect 123240 38560 123400 38720
rect 123240 38720 123400 38880
rect 123240 38880 123400 39040
rect 123240 39040 123400 39200
rect 123240 39200 123400 39360
rect 123240 39360 123400 39520
rect 123240 39520 123400 39680
rect 123240 39680 123400 39840
rect 123240 39840 123400 40000
rect 123240 40000 123400 40160
rect 123240 40160 123400 40320
rect 123240 40320 123400 40480
rect 123240 40480 123400 40640
rect 123240 40640 123400 40800
rect 123240 40800 123400 40960
rect 123240 40960 123400 41120
rect 123240 41120 123400 41280
rect 123240 41280 123400 41440
rect 123240 41440 123400 41600
rect 123240 41600 123400 41760
rect 123240 41760 123400 41920
rect 123240 41920 123400 42080
rect 123240 42080 123400 42240
rect 123240 42240 123400 42400
rect 123240 42400 123400 42560
rect 123240 42560 123400 42720
rect 123240 42720 123400 42880
rect 123240 42880 123400 43040
rect 123240 43040 123400 43200
rect 123240 43200 123400 43360
rect 123240 43360 123400 43520
rect 123240 43520 123400 43680
rect 123240 43680 123400 43840
rect 123400 32480 123560 32640
rect 123400 32640 123560 32800
rect 123400 32800 123560 32960
rect 123400 32960 123560 33120
rect 123400 33120 123560 33280
rect 123400 33280 123560 33440
rect 123400 33440 123560 33600
rect 123400 33600 123560 33760
rect 123400 33760 123560 33920
rect 123400 33920 123560 34080
rect 123400 34080 123560 34240
rect 123400 34240 123560 34400
rect 123400 34400 123560 34560
rect 123400 34560 123560 34720
rect 123400 34720 123560 34880
rect 123400 34880 123560 35040
rect 123400 35040 123560 35200
rect 123400 35200 123560 35360
rect 123400 35360 123560 35520
rect 123400 35520 123560 35680
rect 123400 35680 123560 35840
rect 123400 35840 123560 36000
rect 123400 36000 123560 36160
rect 123400 36160 123560 36320
rect 123400 36320 123560 36480
rect 123400 36480 123560 36640
rect 123400 36640 123560 36800
rect 123400 36800 123560 36960
rect 123400 36960 123560 37120
rect 123400 37120 123560 37280
rect 123400 37280 123560 37440
rect 123400 37440 123560 37600
rect 123400 37600 123560 37760
rect 123400 37760 123560 37920
rect 123400 37920 123560 38080
rect 123400 38080 123560 38240
rect 123400 38240 123560 38400
rect 123400 38400 123560 38560
rect 123400 38560 123560 38720
rect 123400 38720 123560 38880
rect 123400 38880 123560 39040
rect 123400 39040 123560 39200
rect 123400 39200 123560 39360
rect 123400 39360 123560 39520
rect 123400 39520 123560 39680
rect 123400 39680 123560 39840
rect 123400 39840 123560 40000
rect 123400 40000 123560 40160
rect 123400 40160 123560 40320
rect 123400 40320 123560 40480
rect 123400 40480 123560 40640
rect 123400 40640 123560 40800
rect 123400 40800 123560 40960
rect 123400 40960 123560 41120
rect 123400 41120 123560 41280
rect 123400 41280 123560 41440
rect 123400 41440 123560 41600
rect 123400 41600 123560 41760
rect 123400 41760 123560 41920
rect 123400 41920 123560 42080
rect 123400 42080 123560 42240
rect 123400 42240 123560 42400
rect 123400 42400 123560 42560
rect 123400 42560 123560 42720
rect 123400 42720 123560 42880
rect 123400 42880 123560 43040
rect 123400 43040 123560 43200
rect 123400 43200 123560 43360
rect 123400 43360 123560 43520
rect 123400 43520 123560 43680
rect 123400 43680 123560 43840
rect 123400 43840 123560 44000
rect 123400 44000 123560 44160
rect 123400 44160 123560 44320
rect 123560 32000 123720 32160
rect 123560 32160 123720 32320
rect 123560 32320 123720 32480
rect 123560 32480 123720 32640
rect 123560 32640 123720 32800
rect 123560 32800 123720 32960
rect 123560 32960 123720 33120
rect 123560 33120 123720 33280
rect 123560 33280 123720 33440
rect 123560 33440 123720 33600
rect 123560 33600 123720 33760
rect 123560 33760 123720 33920
rect 123560 33920 123720 34080
rect 123560 34080 123720 34240
rect 123560 34240 123720 34400
rect 123560 34400 123720 34560
rect 123560 34560 123720 34720
rect 123560 34720 123720 34880
rect 123560 34880 123720 35040
rect 123560 35040 123720 35200
rect 123560 35200 123720 35360
rect 123560 35360 123720 35520
rect 123560 35520 123720 35680
rect 123560 35680 123720 35840
rect 123560 35840 123720 36000
rect 123560 36000 123720 36160
rect 123560 36160 123720 36320
rect 123560 36320 123720 36480
rect 123560 36480 123720 36640
rect 123560 36640 123720 36800
rect 123560 36800 123720 36960
rect 123560 36960 123720 37120
rect 123560 37120 123720 37280
rect 123560 37280 123720 37440
rect 123560 37440 123720 37600
rect 123560 37600 123720 37760
rect 123560 37760 123720 37920
rect 123560 37920 123720 38080
rect 123560 38080 123720 38240
rect 123560 38240 123720 38400
rect 123560 38400 123720 38560
rect 123560 38560 123720 38720
rect 123560 38720 123720 38880
rect 123560 38880 123720 39040
rect 123560 39040 123720 39200
rect 123560 39200 123720 39360
rect 123560 39360 123720 39520
rect 123560 39520 123720 39680
rect 123560 39680 123720 39840
rect 123560 39840 123720 40000
rect 123560 40000 123720 40160
rect 123560 40160 123720 40320
rect 123560 40320 123720 40480
rect 123560 40480 123720 40640
rect 123560 40640 123720 40800
rect 123560 40800 123720 40960
rect 123560 40960 123720 41120
rect 123560 41120 123720 41280
rect 123560 41280 123720 41440
rect 123560 41440 123720 41600
rect 123560 41600 123720 41760
rect 123560 41760 123720 41920
rect 123560 41920 123720 42080
rect 123560 42080 123720 42240
rect 123560 42240 123720 42400
rect 123560 42400 123720 42560
rect 123560 42560 123720 42720
rect 123560 42720 123720 42880
rect 123560 42880 123720 43040
rect 123560 43040 123720 43200
rect 123560 43200 123720 43360
rect 123560 43360 123720 43520
rect 123560 43520 123720 43680
rect 123560 43680 123720 43840
rect 123560 43840 123720 44000
rect 123560 44000 123720 44160
rect 123560 44160 123720 44320
rect 123560 44320 123720 44480
rect 123560 44480 123720 44640
rect 123560 44640 123720 44800
rect 123720 31680 123880 31840
rect 123720 31840 123880 32000
rect 123720 32000 123880 32160
rect 123720 32160 123880 32320
rect 123720 32320 123880 32480
rect 123720 32480 123880 32640
rect 123720 32640 123880 32800
rect 123720 32800 123880 32960
rect 123720 32960 123880 33120
rect 123720 33120 123880 33280
rect 123720 33280 123880 33440
rect 123720 33440 123880 33600
rect 123720 33600 123880 33760
rect 123720 33760 123880 33920
rect 123720 33920 123880 34080
rect 123720 34080 123880 34240
rect 123720 34240 123880 34400
rect 123720 34400 123880 34560
rect 123720 34560 123880 34720
rect 123720 34720 123880 34880
rect 123720 34880 123880 35040
rect 123720 35040 123880 35200
rect 123720 35200 123880 35360
rect 123720 35360 123880 35520
rect 123720 35520 123880 35680
rect 123720 35680 123880 35840
rect 123720 35840 123880 36000
rect 123720 36000 123880 36160
rect 123720 36160 123880 36320
rect 123720 36320 123880 36480
rect 123720 36480 123880 36640
rect 123720 36640 123880 36800
rect 123720 36800 123880 36960
rect 123720 36960 123880 37120
rect 123720 37120 123880 37280
rect 123720 37280 123880 37440
rect 123720 37440 123880 37600
rect 123720 37600 123880 37760
rect 123720 37760 123880 37920
rect 123720 37920 123880 38080
rect 123720 38080 123880 38240
rect 123720 38240 123880 38400
rect 123720 38400 123880 38560
rect 123720 38560 123880 38720
rect 123720 38720 123880 38880
rect 123720 38880 123880 39040
rect 123720 39040 123880 39200
rect 123720 39200 123880 39360
rect 123720 39360 123880 39520
rect 123720 39520 123880 39680
rect 123720 39680 123880 39840
rect 123720 39840 123880 40000
rect 123720 40000 123880 40160
rect 123720 40160 123880 40320
rect 123720 40320 123880 40480
rect 123720 40480 123880 40640
rect 123720 40640 123880 40800
rect 123720 40800 123880 40960
rect 123720 40960 123880 41120
rect 123720 41120 123880 41280
rect 123720 41280 123880 41440
rect 123720 41440 123880 41600
rect 123720 41600 123880 41760
rect 123720 41760 123880 41920
rect 123720 41920 123880 42080
rect 123720 42080 123880 42240
rect 123720 42240 123880 42400
rect 123720 42400 123880 42560
rect 123720 42560 123880 42720
rect 123720 42720 123880 42880
rect 123720 42880 123880 43040
rect 123720 43040 123880 43200
rect 123720 43200 123880 43360
rect 123720 43360 123880 43520
rect 123720 43520 123880 43680
rect 123720 43680 123880 43840
rect 123720 43840 123880 44000
rect 123720 44000 123880 44160
rect 123720 44160 123880 44320
rect 123720 44320 123880 44480
rect 123720 44480 123880 44640
rect 123720 44640 123880 44800
rect 123720 44800 123880 44960
rect 123720 44960 123880 45120
rect 123720 45120 123880 45280
rect 123880 31520 124040 31680
rect 123880 31680 124040 31840
rect 123880 31840 124040 32000
rect 123880 32000 124040 32160
rect 123880 32160 124040 32320
rect 123880 32320 124040 32480
rect 123880 32480 124040 32640
rect 123880 32640 124040 32800
rect 123880 32800 124040 32960
rect 123880 32960 124040 33120
rect 123880 33120 124040 33280
rect 123880 33280 124040 33440
rect 123880 33440 124040 33600
rect 123880 33600 124040 33760
rect 123880 33760 124040 33920
rect 123880 33920 124040 34080
rect 123880 34080 124040 34240
rect 123880 34240 124040 34400
rect 123880 34400 124040 34560
rect 123880 34560 124040 34720
rect 123880 34720 124040 34880
rect 123880 34880 124040 35040
rect 123880 35040 124040 35200
rect 123880 35200 124040 35360
rect 123880 35360 124040 35520
rect 123880 35520 124040 35680
rect 123880 35680 124040 35840
rect 123880 35840 124040 36000
rect 123880 36000 124040 36160
rect 123880 36160 124040 36320
rect 123880 36320 124040 36480
rect 123880 36480 124040 36640
rect 123880 36640 124040 36800
rect 123880 36800 124040 36960
rect 123880 36960 124040 37120
rect 123880 37120 124040 37280
rect 123880 37280 124040 37440
rect 123880 37440 124040 37600
rect 123880 37600 124040 37760
rect 123880 37760 124040 37920
rect 123880 37920 124040 38080
rect 123880 38080 124040 38240
rect 123880 38240 124040 38400
rect 123880 38400 124040 38560
rect 123880 38560 124040 38720
rect 123880 38720 124040 38880
rect 123880 38880 124040 39040
rect 123880 39040 124040 39200
rect 123880 39200 124040 39360
rect 123880 39360 124040 39520
rect 123880 39520 124040 39680
rect 123880 39680 124040 39840
rect 123880 39840 124040 40000
rect 123880 40000 124040 40160
rect 123880 40160 124040 40320
rect 123880 40320 124040 40480
rect 123880 40480 124040 40640
rect 123880 40640 124040 40800
rect 123880 40800 124040 40960
rect 123880 40960 124040 41120
rect 123880 41120 124040 41280
rect 123880 41280 124040 41440
rect 123880 41440 124040 41600
rect 123880 41600 124040 41760
rect 123880 41760 124040 41920
rect 123880 41920 124040 42080
rect 123880 42080 124040 42240
rect 123880 42240 124040 42400
rect 123880 42400 124040 42560
rect 123880 42560 124040 42720
rect 123880 42720 124040 42880
rect 123880 42880 124040 43040
rect 123880 43040 124040 43200
rect 123880 43200 124040 43360
rect 123880 43360 124040 43520
rect 123880 43520 124040 43680
rect 123880 43680 124040 43840
rect 123880 43840 124040 44000
rect 123880 44000 124040 44160
rect 123880 44160 124040 44320
rect 123880 44320 124040 44480
rect 123880 44480 124040 44640
rect 123880 44640 124040 44800
rect 123880 44800 124040 44960
rect 123880 44960 124040 45120
rect 123880 45120 124040 45280
rect 123880 45280 124040 45440
rect 123880 45440 124040 45600
rect 124040 31200 124200 31360
rect 124040 31360 124200 31520
rect 124040 31520 124200 31680
rect 124040 31680 124200 31840
rect 124040 31840 124200 32000
rect 124040 32000 124200 32160
rect 124040 32160 124200 32320
rect 124040 32320 124200 32480
rect 124040 32480 124200 32640
rect 124040 32640 124200 32800
rect 124040 32800 124200 32960
rect 124040 32960 124200 33120
rect 124040 33120 124200 33280
rect 124040 33280 124200 33440
rect 124040 33440 124200 33600
rect 124040 33600 124200 33760
rect 124040 33760 124200 33920
rect 124040 33920 124200 34080
rect 124040 34080 124200 34240
rect 124040 34240 124200 34400
rect 124040 34400 124200 34560
rect 124040 34560 124200 34720
rect 124040 34720 124200 34880
rect 124040 34880 124200 35040
rect 124040 35040 124200 35200
rect 124040 35200 124200 35360
rect 124040 35360 124200 35520
rect 124040 35520 124200 35680
rect 124040 35680 124200 35840
rect 124040 35840 124200 36000
rect 124040 36000 124200 36160
rect 124040 36160 124200 36320
rect 124040 36320 124200 36480
rect 124040 36480 124200 36640
rect 124040 36640 124200 36800
rect 124040 36800 124200 36960
rect 124040 36960 124200 37120
rect 124040 37120 124200 37280
rect 124040 37280 124200 37440
rect 124040 37440 124200 37600
rect 124040 37600 124200 37760
rect 124040 37760 124200 37920
rect 124040 37920 124200 38080
rect 124040 38080 124200 38240
rect 124040 38240 124200 38400
rect 124040 38400 124200 38560
rect 124040 38560 124200 38720
rect 124040 38720 124200 38880
rect 124040 38880 124200 39040
rect 124040 39040 124200 39200
rect 124040 39200 124200 39360
rect 124040 39360 124200 39520
rect 124040 39520 124200 39680
rect 124040 39680 124200 39840
rect 124040 39840 124200 40000
rect 124040 40000 124200 40160
rect 124040 40160 124200 40320
rect 124040 40320 124200 40480
rect 124040 40480 124200 40640
rect 124040 40640 124200 40800
rect 124040 40800 124200 40960
rect 124040 40960 124200 41120
rect 124040 41120 124200 41280
rect 124040 41280 124200 41440
rect 124040 41440 124200 41600
rect 124040 41600 124200 41760
rect 124040 41760 124200 41920
rect 124040 41920 124200 42080
rect 124040 42080 124200 42240
rect 124040 42240 124200 42400
rect 124040 42400 124200 42560
rect 124040 42560 124200 42720
rect 124040 42720 124200 42880
rect 124040 42880 124200 43040
rect 124040 43040 124200 43200
rect 124040 43200 124200 43360
rect 124040 43360 124200 43520
rect 124040 43520 124200 43680
rect 124040 43680 124200 43840
rect 124040 43840 124200 44000
rect 124040 44000 124200 44160
rect 124040 44160 124200 44320
rect 124040 44320 124200 44480
rect 124040 44480 124200 44640
rect 124040 44640 124200 44800
rect 124040 44800 124200 44960
rect 124040 44960 124200 45120
rect 124040 45120 124200 45280
rect 124040 45280 124200 45440
rect 124040 45440 124200 45600
rect 124040 45600 124200 45760
rect 124040 45760 124200 45920
rect 124200 30880 124360 31040
rect 124200 31040 124360 31200
rect 124200 31200 124360 31360
rect 124200 31360 124360 31520
rect 124200 31520 124360 31680
rect 124200 31680 124360 31840
rect 124200 31840 124360 32000
rect 124200 32000 124360 32160
rect 124200 32160 124360 32320
rect 124200 32320 124360 32480
rect 124200 32480 124360 32640
rect 124200 32640 124360 32800
rect 124200 32800 124360 32960
rect 124200 32960 124360 33120
rect 124200 33120 124360 33280
rect 124200 33280 124360 33440
rect 124200 33440 124360 33600
rect 124200 33600 124360 33760
rect 124200 33760 124360 33920
rect 124200 33920 124360 34080
rect 124200 34080 124360 34240
rect 124200 34240 124360 34400
rect 124200 34400 124360 34560
rect 124200 34560 124360 34720
rect 124200 34720 124360 34880
rect 124200 34880 124360 35040
rect 124200 35040 124360 35200
rect 124200 35200 124360 35360
rect 124200 35360 124360 35520
rect 124200 35520 124360 35680
rect 124200 35680 124360 35840
rect 124200 35840 124360 36000
rect 124200 36000 124360 36160
rect 124200 36160 124360 36320
rect 124200 36320 124360 36480
rect 124200 36480 124360 36640
rect 124200 36640 124360 36800
rect 124200 36800 124360 36960
rect 124200 36960 124360 37120
rect 124200 37120 124360 37280
rect 124200 37280 124360 37440
rect 124200 37440 124360 37600
rect 124200 37600 124360 37760
rect 124200 37760 124360 37920
rect 124200 37920 124360 38080
rect 124200 38080 124360 38240
rect 124200 38240 124360 38400
rect 124200 38400 124360 38560
rect 124200 38560 124360 38720
rect 124200 38720 124360 38880
rect 124200 38880 124360 39040
rect 124200 39040 124360 39200
rect 124200 39200 124360 39360
rect 124200 39360 124360 39520
rect 124200 39520 124360 39680
rect 124200 39680 124360 39840
rect 124200 39840 124360 40000
rect 124200 40000 124360 40160
rect 124200 40160 124360 40320
rect 124200 40320 124360 40480
rect 124200 40480 124360 40640
rect 124200 40640 124360 40800
rect 124200 40800 124360 40960
rect 124200 40960 124360 41120
rect 124200 41120 124360 41280
rect 124200 41280 124360 41440
rect 124200 41440 124360 41600
rect 124200 41600 124360 41760
rect 124200 41760 124360 41920
rect 124200 41920 124360 42080
rect 124200 42080 124360 42240
rect 124200 42240 124360 42400
rect 124200 42400 124360 42560
rect 124200 42560 124360 42720
rect 124200 42720 124360 42880
rect 124200 42880 124360 43040
rect 124200 43040 124360 43200
rect 124200 43200 124360 43360
rect 124200 43360 124360 43520
rect 124200 43520 124360 43680
rect 124200 43680 124360 43840
rect 124200 43840 124360 44000
rect 124200 44000 124360 44160
rect 124200 44160 124360 44320
rect 124200 44320 124360 44480
rect 124200 44480 124360 44640
rect 124200 44640 124360 44800
rect 124200 44800 124360 44960
rect 124200 44960 124360 45120
rect 124200 45120 124360 45280
rect 124200 45280 124360 45440
rect 124200 45440 124360 45600
rect 124200 45600 124360 45760
rect 124200 45760 124360 45920
rect 124200 45920 124360 46080
rect 124200 46080 124360 46240
rect 124360 30720 124520 30880
rect 124360 30880 124520 31040
rect 124360 31040 124520 31200
rect 124360 31200 124520 31360
rect 124360 31360 124520 31520
rect 124360 31520 124520 31680
rect 124360 31680 124520 31840
rect 124360 31840 124520 32000
rect 124360 32000 124520 32160
rect 124360 32160 124520 32320
rect 124360 32320 124520 32480
rect 124360 32480 124520 32640
rect 124360 32640 124520 32800
rect 124360 32800 124520 32960
rect 124360 32960 124520 33120
rect 124360 33120 124520 33280
rect 124360 33280 124520 33440
rect 124360 33440 124520 33600
rect 124360 33600 124520 33760
rect 124360 33760 124520 33920
rect 124360 33920 124520 34080
rect 124360 34080 124520 34240
rect 124360 34240 124520 34400
rect 124360 34400 124520 34560
rect 124360 34560 124520 34720
rect 124360 34720 124520 34880
rect 124360 34880 124520 35040
rect 124360 35040 124520 35200
rect 124360 35200 124520 35360
rect 124360 35360 124520 35520
rect 124360 35520 124520 35680
rect 124360 35680 124520 35840
rect 124360 35840 124520 36000
rect 124360 36000 124520 36160
rect 124360 36160 124520 36320
rect 124360 36320 124520 36480
rect 124360 36480 124520 36640
rect 124360 36640 124520 36800
rect 124360 36800 124520 36960
rect 124360 36960 124520 37120
rect 124360 37120 124520 37280
rect 124360 37280 124520 37440
rect 124360 37440 124520 37600
rect 124360 37600 124520 37760
rect 124360 37760 124520 37920
rect 124360 37920 124520 38080
rect 124360 38080 124520 38240
rect 124360 38240 124520 38400
rect 124360 38400 124520 38560
rect 124360 38560 124520 38720
rect 124360 38720 124520 38880
rect 124360 38880 124520 39040
rect 124360 39040 124520 39200
rect 124360 39200 124520 39360
rect 124360 39360 124520 39520
rect 124360 39520 124520 39680
rect 124360 39680 124520 39840
rect 124360 39840 124520 40000
rect 124360 40000 124520 40160
rect 124360 40160 124520 40320
rect 124360 40320 124520 40480
rect 124360 40480 124520 40640
rect 124360 40640 124520 40800
rect 124360 40800 124520 40960
rect 124360 40960 124520 41120
rect 124360 41120 124520 41280
rect 124360 41280 124520 41440
rect 124360 41440 124520 41600
rect 124360 41600 124520 41760
rect 124360 41760 124520 41920
rect 124360 41920 124520 42080
rect 124360 42080 124520 42240
rect 124360 42240 124520 42400
rect 124360 42400 124520 42560
rect 124360 42560 124520 42720
rect 124360 42720 124520 42880
rect 124360 42880 124520 43040
rect 124360 43040 124520 43200
rect 124360 43200 124520 43360
rect 124360 43360 124520 43520
rect 124360 43520 124520 43680
rect 124360 43680 124520 43840
rect 124360 43840 124520 44000
rect 124360 44000 124520 44160
rect 124360 44160 124520 44320
rect 124360 44320 124520 44480
rect 124360 44480 124520 44640
rect 124360 44640 124520 44800
rect 124360 44800 124520 44960
rect 124360 44960 124520 45120
rect 124360 45120 124520 45280
rect 124360 45280 124520 45440
rect 124360 45440 124520 45600
rect 124360 45600 124520 45760
rect 124360 45760 124520 45920
rect 124360 45920 124520 46080
rect 124360 46080 124520 46240
rect 124360 46240 124520 46400
rect 124360 46400 124520 46560
rect 124520 30560 124680 30720
rect 124520 30720 124680 30880
rect 124520 30880 124680 31040
rect 124520 31040 124680 31200
rect 124520 31200 124680 31360
rect 124520 31360 124680 31520
rect 124520 31520 124680 31680
rect 124520 31680 124680 31840
rect 124520 31840 124680 32000
rect 124520 32000 124680 32160
rect 124520 32160 124680 32320
rect 124520 32320 124680 32480
rect 124520 32480 124680 32640
rect 124520 32640 124680 32800
rect 124520 32800 124680 32960
rect 124520 32960 124680 33120
rect 124520 33120 124680 33280
rect 124520 33280 124680 33440
rect 124520 33440 124680 33600
rect 124520 33600 124680 33760
rect 124520 33760 124680 33920
rect 124520 33920 124680 34080
rect 124520 34080 124680 34240
rect 124520 34240 124680 34400
rect 124520 34400 124680 34560
rect 124520 34560 124680 34720
rect 124520 34720 124680 34880
rect 124520 34880 124680 35040
rect 124520 35040 124680 35200
rect 124520 35200 124680 35360
rect 124520 35360 124680 35520
rect 124520 35520 124680 35680
rect 124520 35680 124680 35840
rect 124520 35840 124680 36000
rect 124520 36000 124680 36160
rect 124520 36160 124680 36320
rect 124520 36320 124680 36480
rect 124520 36480 124680 36640
rect 124520 36640 124680 36800
rect 124520 36800 124680 36960
rect 124520 36960 124680 37120
rect 124520 37120 124680 37280
rect 124520 37280 124680 37440
rect 124520 37440 124680 37600
rect 124520 37600 124680 37760
rect 124520 37760 124680 37920
rect 124520 37920 124680 38080
rect 124520 38080 124680 38240
rect 124520 38240 124680 38400
rect 124520 38400 124680 38560
rect 124520 38560 124680 38720
rect 124520 38720 124680 38880
rect 124520 38880 124680 39040
rect 124520 39040 124680 39200
rect 124520 39200 124680 39360
rect 124520 39360 124680 39520
rect 124520 39520 124680 39680
rect 124520 39680 124680 39840
rect 124520 39840 124680 40000
rect 124520 40000 124680 40160
rect 124520 40160 124680 40320
rect 124520 40320 124680 40480
rect 124520 40480 124680 40640
rect 124520 40640 124680 40800
rect 124520 40800 124680 40960
rect 124520 40960 124680 41120
rect 124520 41120 124680 41280
rect 124520 41280 124680 41440
rect 124520 41440 124680 41600
rect 124520 41600 124680 41760
rect 124520 41760 124680 41920
rect 124520 41920 124680 42080
rect 124520 42080 124680 42240
rect 124520 42240 124680 42400
rect 124520 42400 124680 42560
rect 124520 42560 124680 42720
rect 124520 42720 124680 42880
rect 124520 42880 124680 43040
rect 124520 43040 124680 43200
rect 124520 43200 124680 43360
rect 124520 43360 124680 43520
rect 124520 43520 124680 43680
rect 124520 43680 124680 43840
rect 124520 43840 124680 44000
rect 124520 44000 124680 44160
rect 124520 44160 124680 44320
rect 124520 44320 124680 44480
rect 124520 44480 124680 44640
rect 124520 44640 124680 44800
rect 124520 44800 124680 44960
rect 124520 44960 124680 45120
rect 124520 45120 124680 45280
rect 124520 45280 124680 45440
rect 124520 45440 124680 45600
rect 124520 45600 124680 45760
rect 124520 45760 124680 45920
rect 124520 45920 124680 46080
rect 124520 46080 124680 46240
rect 124520 46240 124680 46400
rect 124520 46400 124680 46560
rect 124520 46560 124680 46720
rect 124520 46720 124680 46880
rect 124680 30240 124840 30400
rect 124680 30400 124840 30560
rect 124680 30560 124840 30720
rect 124680 30720 124840 30880
rect 124680 30880 124840 31040
rect 124680 31040 124840 31200
rect 124680 31200 124840 31360
rect 124680 31360 124840 31520
rect 124680 31520 124840 31680
rect 124680 31680 124840 31840
rect 124680 31840 124840 32000
rect 124680 32000 124840 32160
rect 124680 32160 124840 32320
rect 124680 32320 124840 32480
rect 124680 32480 124840 32640
rect 124680 32640 124840 32800
rect 124680 32800 124840 32960
rect 124680 32960 124840 33120
rect 124680 33120 124840 33280
rect 124680 33280 124840 33440
rect 124680 33440 124840 33600
rect 124680 33600 124840 33760
rect 124680 33760 124840 33920
rect 124680 33920 124840 34080
rect 124680 34080 124840 34240
rect 124680 34240 124840 34400
rect 124680 34400 124840 34560
rect 124680 34560 124840 34720
rect 124680 34720 124840 34880
rect 124680 34880 124840 35040
rect 124680 35040 124840 35200
rect 124680 35200 124840 35360
rect 124680 35360 124840 35520
rect 124680 35520 124840 35680
rect 124680 35680 124840 35840
rect 124680 35840 124840 36000
rect 124680 36000 124840 36160
rect 124680 36160 124840 36320
rect 124680 36320 124840 36480
rect 124680 36480 124840 36640
rect 124680 36640 124840 36800
rect 124680 36800 124840 36960
rect 124680 36960 124840 37120
rect 124680 37120 124840 37280
rect 124680 37280 124840 37440
rect 124680 37440 124840 37600
rect 124680 37600 124840 37760
rect 124680 37760 124840 37920
rect 124680 37920 124840 38080
rect 124680 38080 124840 38240
rect 124680 38240 124840 38400
rect 124680 38400 124840 38560
rect 124680 38560 124840 38720
rect 124680 38720 124840 38880
rect 124680 38880 124840 39040
rect 124680 39040 124840 39200
rect 124680 39200 124840 39360
rect 124680 39360 124840 39520
rect 124680 39520 124840 39680
rect 124680 39680 124840 39840
rect 124680 39840 124840 40000
rect 124680 40000 124840 40160
rect 124680 40160 124840 40320
rect 124680 40320 124840 40480
rect 124680 40480 124840 40640
rect 124680 40640 124840 40800
rect 124680 40800 124840 40960
rect 124680 40960 124840 41120
rect 124680 41120 124840 41280
rect 124680 41280 124840 41440
rect 124680 41440 124840 41600
rect 124680 41600 124840 41760
rect 124680 41760 124840 41920
rect 124680 41920 124840 42080
rect 124680 42080 124840 42240
rect 124680 42240 124840 42400
rect 124680 42400 124840 42560
rect 124680 42560 124840 42720
rect 124680 42720 124840 42880
rect 124680 42880 124840 43040
rect 124680 43040 124840 43200
rect 124680 43200 124840 43360
rect 124680 43360 124840 43520
rect 124680 43520 124840 43680
rect 124680 43680 124840 43840
rect 124680 43840 124840 44000
rect 124680 44000 124840 44160
rect 124680 44160 124840 44320
rect 124680 44320 124840 44480
rect 124680 44480 124840 44640
rect 124680 44640 124840 44800
rect 124680 44800 124840 44960
rect 124680 44960 124840 45120
rect 124680 45120 124840 45280
rect 124680 45280 124840 45440
rect 124680 45440 124840 45600
rect 124680 45600 124840 45760
rect 124680 45760 124840 45920
rect 124680 45920 124840 46080
rect 124680 46080 124840 46240
rect 124680 46240 124840 46400
rect 124680 46400 124840 46560
rect 124680 46560 124840 46720
rect 124680 46720 124840 46880
rect 124680 46880 124840 47040
rect 124680 47040 124840 47200
rect 124840 30080 125000 30240
rect 124840 30240 125000 30400
rect 124840 30400 125000 30560
rect 124840 30560 125000 30720
rect 124840 30720 125000 30880
rect 124840 30880 125000 31040
rect 124840 31040 125000 31200
rect 124840 31200 125000 31360
rect 124840 31360 125000 31520
rect 124840 31520 125000 31680
rect 124840 31680 125000 31840
rect 124840 31840 125000 32000
rect 124840 32000 125000 32160
rect 124840 32160 125000 32320
rect 124840 32320 125000 32480
rect 124840 32480 125000 32640
rect 124840 32640 125000 32800
rect 124840 32800 125000 32960
rect 124840 32960 125000 33120
rect 124840 33120 125000 33280
rect 124840 33280 125000 33440
rect 124840 33440 125000 33600
rect 124840 33600 125000 33760
rect 124840 33760 125000 33920
rect 124840 33920 125000 34080
rect 124840 34080 125000 34240
rect 124840 34240 125000 34400
rect 124840 34400 125000 34560
rect 124840 34560 125000 34720
rect 124840 34720 125000 34880
rect 124840 34880 125000 35040
rect 124840 35040 125000 35200
rect 124840 35200 125000 35360
rect 124840 35360 125000 35520
rect 124840 35520 125000 35680
rect 124840 35680 125000 35840
rect 124840 35840 125000 36000
rect 124840 36000 125000 36160
rect 124840 36160 125000 36320
rect 124840 36320 125000 36480
rect 124840 36480 125000 36640
rect 124840 36640 125000 36800
rect 124840 36800 125000 36960
rect 124840 36960 125000 37120
rect 124840 37120 125000 37280
rect 124840 37280 125000 37440
rect 124840 37440 125000 37600
rect 124840 37600 125000 37760
rect 124840 37760 125000 37920
rect 124840 37920 125000 38080
rect 124840 38080 125000 38240
rect 124840 38240 125000 38400
rect 124840 38400 125000 38560
rect 124840 38560 125000 38720
rect 124840 38720 125000 38880
rect 124840 38880 125000 39040
rect 124840 39040 125000 39200
rect 124840 39200 125000 39360
rect 124840 39360 125000 39520
rect 124840 39520 125000 39680
rect 124840 39680 125000 39840
rect 124840 39840 125000 40000
rect 124840 40000 125000 40160
rect 124840 40160 125000 40320
rect 124840 40320 125000 40480
rect 124840 40480 125000 40640
rect 124840 40640 125000 40800
rect 124840 40800 125000 40960
rect 124840 40960 125000 41120
rect 124840 41120 125000 41280
rect 124840 41280 125000 41440
rect 124840 41440 125000 41600
rect 124840 41600 125000 41760
rect 124840 41760 125000 41920
rect 124840 41920 125000 42080
rect 124840 42080 125000 42240
rect 124840 42240 125000 42400
rect 124840 42400 125000 42560
rect 124840 42560 125000 42720
rect 124840 42720 125000 42880
rect 124840 42880 125000 43040
rect 124840 43040 125000 43200
rect 124840 43200 125000 43360
rect 124840 43360 125000 43520
rect 124840 43520 125000 43680
rect 124840 43680 125000 43840
rect 124840 43840 125000 44000
rect 124840 44000 125000 44160
rect 124840 44160 125000 44320
rect 124840 44320 125000 44480
rect 124840 44480 125000 44640
rect 124840 44640 125000 44800
rect 124840 44800 125000 44960
rect 124840 44960 125000 45120
rect 124840 45120 125000 45280
rect 124840 45280 125000 45440
rect 124840 45440 125000 45600
rect 124840 45600 125000 45760
rect 124840 45760 125000 45920
rect 124840 45920 125000 46080
rect 124840 46080 125000 46240
rect 124840 46240 125000 46400
rect 124840 46400 125000 46560
rect 124840 46560 125000 46720
rect 124840 46720 125000 46880
rect 124840 46880 125000 47040
rect 124840 47040 125000 47200
rect 124840 47200 125000 47360
rect 124840 47360 125000 47520
rect 125000 29920 125160 30080
rect 125000 30080 125160 30240
rect 125000 30240 125160 30400
rect 125000 30400 125160 30560
rect 125000 30560 125160 30720
rect 125000 30720 125160 30880
rect 125000 30880 125160 31040
rect 125000 31040 125160 31200
rect 125000 31200 125160 31360
rect 125000 31360 125160 31520
rect 125000 31520 125160 31680
rect 125000 31680 125160 31840
rect 125000 31840 125160 32000
rect 125000 32000 125160 32160
rect 125000 32160 125160 32320
rect 125000 32320 125160 32480
rect 125000 32480 125160 32640
rect 125000 32640 125160 32800
rect 125000 32800 125160 32960
rect 125000 32960 125160 33120
rect 125000 33120 125160 33280
rect 125000 33280 125160 33440
rect 125000 33440 125160 33600
rect 125000 33600 125160 33760
rect 125000 33760 125160 33920
rect 125000 33920 125160 34080
rect 125000 34080 125160 34240
rect 125000 34240 125160 34400
rect 125000 34400 125160 34560
rect 125000 34560 125160 34720
rect 125000 34720 125160 34880
rect 125000 34880 125160 35040
rect 125000 35040 125160 35200
rect 125000 35200 125160 35360
rect 125000 35360 125160 35520
rect 125000 35520 125160 35680
rect 125000 35680 125160 35840
rect 125000 35840 125160 36000
rect 125000 36000 125160 36160
rect 125000 36160 125160 36320
rect 125000 36320 125160 36480
rect 125000 36480 125160 36640
rect 125000 36640 125160 36800
rect 125000 36800 125160 36960
rect 125000 36960 125160 37120
rect 125000 37120 125160 37280
rect 125000 37280 125160 37440
rect 125000 37440 125160 37600
rect 125000 37600 125160 37760
rect 125000 37760 125160 37920
rect 125000 37920 125160 38080
rect 125000 38080 125160 38240
rect 125000 38240 125160 38400
rect 125000 38400 125160 38560
rect 125000 38560 125160 38720
rect 125000 38720 125160 38880
rect 125000 38880 125160 39040
rect 125000 39040 125160 39200
rect 125000 39200 125160 39360
rect 125000 39360 125160 39520
rect 125000 39520 125160 39680
rect 125000 39680 125160 39840
rect 125000 39840 125160 40000
rect 125000 40000 125160 40160
rect 125000 40160 125160 40320
rect 125000 40320 125160 40480
rect 125000 40480 125160 40640
rect 125000 40640 125160 40800
rect 125000 40800 125160 40960
rect 125000 40960 125160 41120
rect 125000 41120 125160 41280
rect 125000 41280 125160 41440
rect 125000 41440 125160 41600
rect 125000 41600 125160 41760
rect 125000 41760 125160 41920
rect 125000 41920 125160 42080
rect 125000 42080 125160 42240
rect 125000 42240 125160 42400
rect 125000 42400 125160 42560
rect 125000 42560 125160 42720
rect 125000 42720 125160 42880
rect 125000 42880 125160 43040
rect 125000 43040 125160 43200
rect 125000 43200 125160 43360
rect 125000 43360 125160 43520
rect 125000 43520 125160 43680
rect 125000 43680 125160 43840
rect 125000 43840 125160 44000
rect 125000 44000 125160 44160
rect 125000 44160 125160 44320
rect 125000 44320 125160 44480
rect 125000 44480 125160 44640
rect 125000 44640 125160 44800
rect 125000 44800 125160 44960
rect 125000 44960 125160 45120
rect 125000 45120 125160 45280
rect 125000 45280 125160 45440
rect 125000 45440 125160 45600
rect 125000 45600 125160 45760
rect 125000 45760 125160 45920
rect 125000 45920 125160 46080
rect 125000 46080 125160 46240
rect 125000 46240 125160 46400
rect 125000 46400 125160 46560
rect 125000 46560 125160 46720
rect 125000 46720 125160 46880
rect 125000 46880 125160 47040
rect 125000 47040 125160 47200
rect 125000 47200 125160 47360
rect 125000 47360 125160 47520
rect 125000 47520 125160 47680
rect 125000 47680 125160 47840
rect 125160 29760 125320 29920
rect 125160 29920 125320 30080
rect 125160 30080 125320 30240
rect 125160 30240 125320 30400
rect 125160 30400 125320 30560
rect 125160 30560 125320 30720
rect 125160 30720 125320 30880
rect 125160 30880 125320 31040
rect 125160 31040 125320 31200
rect 125160 31200 125320 31360
rect 125160 31360 125320 31520
rect 125160 31520 125320 31680
rect 125160 31680 125320 31840
rect 125160 31840 125320 32000
rect 125160 32000 125320 32160
rect 125160 32160 125320 32320
rect 125160 32320 125320 32480
rect 125160 32480 125320 32640
rect 125160 32640 125320 32800
rect 125160 32800 125320 32960
rect 125160 32960 125320 33120
rect 125160 33120 125320 33280
rect 125160 33280 125320 33440
rect 125160 33440 125320 33600
rect 125160 33600 125320 33760
rect 125160 33760 125320 33920
rect 125160 33920 125320 34080
rect 125160 34080 125320 34240
rect 125160 34240 125320 34400
rect 125160 34400 125320 34560
rect 125160 34560 125320 34720
rect 125160 34720 125320 34880
rect 125160 34880 125320 35040
rect 125160 35040 125320 35200
rect 125160 35200 125320 35360
rect 125160 35360 125320 35520
rect 125160 35520 125320 35680
rect 125160 35680 125320 35840
rect 125160 35840 125320 36000
rect 125160 36000 125320 36160
rect 125160 36160 125320 36320
rect 125160 36320 125320 36480
rect 125160 36480 125320 36640
rect 125160 36640 125320 36800
rect 125160 36800 125320 36960
rect 125160 36960 125320 37120
rect 125160 37120 125320 37280
rect 125160 37280 125320 37440
rect 125160 37440 125320 37600
rect 125160 37600 125320 37760
rect 125160 37760 125320 37920
rect 125160 37920 125320 38080
rect 125160 38080 125320 38240
rect 125160 38240 125320 38400
rect 125160 38400 125320 38560
rect 125160 38560 125320 38720
rect 125160 38720 125320 38880
rect 125160 38880 125320 39040
rect 125160 39040 125320 39200
rect 125160 39200 125320 39360
rect 125160 39360 125320 39520
rect 125160 39520 125320 39680
rect 125160 39680 125320 39840
rect 125160 39840 125320 40000
rect 125160 40000 125320 40160
rect 125160 40160 125320 40320
rect 125160 40320 125320 40480
rect 125160 40480 125320 40640
rect 125160 40640 125320 40800
rect 125160 40800 125320 40960
rect 125160 40960 125320 41120
rect 125160 41120 125320 41280
rect 125160 41280 125320 41440
rect 125160 41440 125320 41600
rect 125160 41600 125320 41760
rect 125160 41760 125320 41920
rect 125160 41920 125320 42080
rect 125160 42080 125320 42240
rect 125160 42240 125320 42400
rect 125160 42400 125320 42560
rect 125160 42560 125320 42720
rect 125160 42720 125320 42880
rect 125160 42880 125320 43040
rect 125160 43040 125320 43200
rect 125160 43200 125320 43360
rect 125160 43360 125320 43520
rect 125160 43520 125320 43680
rect 125160 43680 125320 43840
rect 125160 43840 125320 44000
rect 125160 44000 125320 44160
rect 125160 44160 125320 44320
rect 125160 44320 125320 44480
rect 125160 44480 125320 44640
rect 125160 44640 125320 44800
rect 125160 44800 125320 44960
rect 125160 44960 125320 45120
rect 125160 45120 125320 45280
rect 125160 45280 125320 45440
rect 125160 45440 125320 45600
rect 125160 45600 125320 45760
rect 125160 45760 125320 45920
rect 125160 45920 125320 46080
rect 125160 46080 125320 46240
rect 125160 46240 125320 46400
rect 125160 46400 125320 46560
rect 125160 46560 125320 46720
rect 125160 46720 125320 46880
rect 125160 46880 125320 47040
rect 125160 47040 125320 47200
rect 125160 47200 125320 47360
rect 125160 47360 125320 47520
rect 125160 47520 125320 47680
rect 125160 47680 125320 47840
rect 125160 47840 125320 48000
rect 125320 29600 125480 29760
rect 125320 29760 125480 29920
rect 125320 29920 125480 30080
rect 125320 30080 125480 30240
rect 125320 30240 125480 30400
rect 125320 30400 125480 30560
rect 125320 30560 125480 30720
rect 125320 30720 125480 30880
rect 125320 30880 125480 31040
rect 125320 31040 125480 31200
rect 125320 31200 125480 31360
rect 125320 31360 125480 31520
rect 125320 31520 125480 31680
rect 125320 31680 125480 31840
rect 125320 31840 125480 32000
rect 125320 32000 125480 32160
rect 125320 32160 125480 32320
rect 125320 32320 125480 32480
rect 125320 32480 125480 32640
rect 125320 32640 125480 32800
rect 125320 32800 125480 32960
rect 125320 32960 125480 33120
rect 125320 33120 125480 33280
rect 125320 33280 125480 33440
rect 125320 33440 125480 33600
rect 125320 33600 125480 33760
rect 125320 33760 125480 33920
rect 125320 33920 125480 34080
rect 125320 34080 125480 34240
rect 125320 34240 125480 34400
rect 125320 34400 125480 34560
rect 125320 34560 125480 34720
rect 125320 34720 125480 34880
rect 125320 34880 125480 35040
rect 125320 35040 125480 35200
rect 125320 35200 125480 35360
rect 125320 35360 125480 35520
rect 125320 35520 125480 35680
rect 125320 35680 125480 35840
rect 125320 35840 125480 36000
rect 125320 36000 125480 36160
rect 125320 36160 125480 36320
rect 125320 36320 125480 36480
rect 125320 36480 125480 36640
rect 125320 36640 125480 36800
rect 125320 36800 125480 36960
rect 125320 36960 125480 37120
rect 125320 37120 125480 37280
rect 125320 37280 125480 37440
rect 125320 37440 125480 37600
rect 125320 37600 125480 37760
rect 125320 37760 125480 37920
rect 125320 37920 125480 38080
rect 125320 38080 125480 38240
rect 125320 38240 125480 38400
rect 125320 38400 125480 38560
rect 125320 38560 125480 38720
rect 125320 38720 125480 38880
rect 125320 38880 125480 39040
rect 125320 39040 125480 39200
rect 125320 39200 125480 39360
rect 125320 39360 125480 39520
rect 125320 39520 125480 39680
rect 125320 39680 125480 39840
rect 125320 39840 125480 40000
rect 125320 40000 125480 40160
rect 125320 40160 125480 40320
rect 125320 40320 125480 40480
rect 125320 40480 125480 40640
rect 125320 40640 125480 40800
rect 125320 40800 125480 40960
rect 125320 40960 125480 41120
rect 125320 41120 125480 41280
rect 125320 41280 125480 41440
rect 125320 41440 125480 41600
rect 125320 41600 125480 41760
rect 125320 41760 125480 41920
rect 125320 41920 125480 42080
rect 125320 42080 125480 42240
rect 125320 42240 125480 42400
rect 125320 42400 125480 42560
rect 125320 42560 125480 42720
rect 125320 42720 125480 42880
rect 125320 42880 125480 43040
rect 125320 43040 125480 43200
rect 125320 43200 125480 43360
rect 125320 43360 125480 43520
rect 125320 43520 125480 43680
rect 125320 43680 125480 43840
rect 125320 43840 125480 44000
rect 125320 44000 125480 44160
rect 125320 44160 125480 44320
rect 125320 44320 125480 44480
rect 125320 44480 125480 44640
rect 125320 44640 125480 44800
rect 125320 44800 125480 44960
rect 125320 44960 125480 45120
rect 125320 45120 125480 45280
rect 125320 45280 125480 45440
rect 125320 45440 125480 45600
rect 125320 45600 125480 45760
rect 125320 45760 125480 45920
rect 125320 45920 125480 46080
rect 125320 46080 125480 46240
rect 125320 46240 125480 46400
rect 125320 46400 125480 46560
rect 125320 46560 125480 46720
rect 125320 46720 125480 46880
rect 125320 46880 125480 47040
rect 125320 47040 125480 47200
rect 125320 47200 125480 47360
rect 125320 47360 125480 47520
rect 125320 47520 125480 47680
rect 125320 47680 125480 47840
rect 125320 47840 125480 48000
rect 125320 48000 125480 48160
rect 125320 48160 125480 48320
rect 125480 29440 125640 29600
rect 125480 29600 125640 29760
rect 125480 29760 125640 29920
rect 125480 29920 125640 30080
rect 125480 30080 125640 30240
rect 125480 30240 125640 30400
rect 125480 30400 125640 30560
rect 125480 30560 125640 30720
rect 125480 30720 125640 30880
rect 125480 30880 125640 31040
rect 125480 31040 125640 31200
rect 125480 31200 125640 31360
rect 125480 31360 125640 31520
rect 125480 31520 125640 31680
rect 125480 31680 125640 31840
rect 125480 31840 125640 32000
rect 125480 32000 125640 32160
rect 125480 32160 125640 32320
rect 125480 32320 125640 32480
rect 125480 32480 125640 32640
rect 125480 32640 125640 32800
rect 125480 32800 125640 32960
rect 125480 32960 125640 33120
rect 125480 33120 125640 33280
rect 125480 33280 125640 33440
rect 125480 33440 125640 33600
rect 125480 33600 125640 33760
rect 125480 33760 125640 33920
rect 125480 33920 125640 34080
rect 125480 34080 125640 34240
rect 125480 34240 125640 34400
rect 125480 34400 125640 34560
rect 125480 34560 125640 34720
rect 125480 34720 125640 34880
rect 125480 34880 125640 35040
rect 125480 35040 125640 35200
rect 125480 35200 125640 35360
rect 125480 35360 125640 35520
rect 125480 35520 125640 35680
rect 125480 35680 125640 35840
rect 125480 35840 125640 36000
rect 125480 36000 125640 36160
rect 125480 36160 125640 36320
rect 125480 36320 125640 36480
rect 125480 36480 125640 36640
rect 125480 36640 125640 36800
rect 125480 36800 125640 36960
rect 125480 36960 125640 37120
rect 125480 37120 125640 37280
rect 125480 37280 125640 37440
rect 125480 37440 125640 37600
rect 125480 37600 125640 37760
rect 125480 37760 125640 37920
rect 125480 37920 125640 38080
rect 125480 38080 125640 38240
rect 125480 38240 125640 38400
rect 125480 38400 125640 38560
rect 125480 38560 125640 38720
rect 125480 38720 125640 38880
rect 125480 38880 125640 39040
rect 125480 39040 125640 39200
rect 125480 39200 125640 39360
rect 125480 39360 125640 39520
rect 125480 39520 125640 39680
rect 125480 39680 125640 39840
rect 125480 39840 125640 40000
rect 125480 40000 125640 40160
rect 125480 40160 125640 40320
rect 125480 40320 125640 40480
rect 125480 40480 125640 40640
rect 125480 40640 125640 40800
rect 125480 40800 125640 40960
rect 125480 40960 125640 41120
rect 125480 41120 125640 41280
rect 125480 41280 125640 41440
rect 125480 41440 125640 41600
rect 125480 41600 125640 41760
rect 125480 41760 125640 41920
rect 125480 41920 125640 42080
rect 125480 42080 125640 42240
rect 125480 42240 125640 42400
rect 125480 42400 125640 42560
rect 125480 42560 125640 42720
rect 125480 42720 125640 42880
rect 125480 42880 125640 43040
rect 125480 43040 125640 43200
rect 125480 43200 125640 43360
rect 125480 43360 125640 43520
rect 125480 43520 125640 43680
rect 125480 43680 125640 43840
rect 125480 43840 125640 44000
rect 125480 44000 125640 44160
rect 125480 44160 125640 44320
rect 125480 44320 125640 44480
rect 125480 44480 125640 44640
rect 125480 44640 125640 44800
rect 125480 44800 125640 44960
rect 125480 44960 125640 45120
rect 125480 45120 125640 45280
rect 125480 45280 125640 45440
rect 125480 45440 125640 45600
rect 125480 45600 125640 45760
rect 125480 45760 125640 45920
rect 125480 45920 125640 46080
rect 125480 46080 125640 46240
rect 125480 46240 125640 46400
rect 125480 46400 125640 46560
rect 125480 46560 125640 46720
rect 125480 46720 125640 46880
rect 125480 46880 125640 47040
rect 125480 47040 125640 47200
rect 125480 47200 125640 47360
rect 125480 47360 125640 47520
rect 125480 47520 125640 47680
rect 125480 47680 125640 47840
rect 125480 47840 125640 48000
rect 125480 48000 125640 48160
rect 125480 48160 125640 48320
rect 125480 48320 125640 48480
rect 125640 29280 125800 29440
rect 125640 29440 125800 29600
rect 125640 29600 125800 29760
rect 125640 29760 125800 29920
rect 125640 29920 125800 30080
rect 125640 30080 125800 30240
rect 125640 30240 125800 30400
rect 125640 30400 125800 30560
rect 125640 30560 125800 30720
rect 125640 30720 125800 30880
rect 125640 30880 125800 31040
rect 125640 31040 125800 31200
rect 125640 31200 125800 31360
rect 125640 31360 125800 31520
rect 125640 31520 125800 31680
rect 125640 31680 125800 31840
rect 125640 31840 125800 32000
rect 125640 32000 125800 32160
rect 125640 32160 125800 32320
rect 125640 32320 125800 32480
rect 125640 32480 125800 32640
rect 125640 32640 125800 32800
rect 125640 32800 125800 32960
rect 125640 32960 125800 33120
rect 125640 33120 125800 33280
rect 125640 33280 125800 33440
rect 125640 33440 125800 33600
rect 125640 33600 125800 33760
rect 125640 33760 125800 33920
rect 125640 33920 125800 34080
rect 125640 34080 125800 34240
rect 125640 34240 125800 34400
rect 125640 34400 125800 34560
rect 125640 34560 125800 34720
rect 125640 34720 125800 34880
rect 125640 34880 125800 35040
rect 125640 35040 125800 35200
rect 125640 35200 125800 35360
rect 125640 35360 125800 35520
rect 125640 35520 125800 35680
rect 125640 35680 125800 35840
rect 125640 35840 125800 36000
rect 125640 36000 125800 36160
rect 125640 36160 125800 36320
rect 125640 36320 125800 36480
rect 125640 36480 125800 36640
rect 125640 36640 125800 36800
rect 125640 36960 125800 37120
rect 125640 39360 125800 39520
rect 125640 39520 125800 39680
rect 125640 39680 125800 39840
rect 125640 39840 125800 40000
rect 125640 40000 125800 40160
rect 125640 40160 125800 40320
rect 125640 40320 125800 40480
rect 125640 40480 125800 40640
rect 125640 40640 125800 40800
rect 125640 40800 125800 40960
rect 125640 40960 125800 41120
rect 125640 41120 125800 41280
rect 125640 41280 125800 41440
rect 125640 41440 125800 41600
rect 125640 41600 125800 41760
rect 125640 41760 125800 41920
rect 125640 41920 125800 42080
rect 125640 42080 125800 42240
rect 125640 42240 125800 42400
rect 125640 42400 125800 42560
rect 125640 42560 125800 42720
rect 125640 42720 125800 42880
rect 125640 42880 125800 43040
rect 125640 43040 125800 43200
rect 125640 43200 125800 43360
rect 125640 43360 125800 43520
rect 125640 43520 125800 43680
rect 125640 43680 125800 43840
rect 125640 43840 125800 44000
rect 125640 44000 125800 44160
rect 125640 44160 125800 44320
rect 125640 44320 125800 44480
rect 125640 44480 125800 44640
rect 125640 44640 125800 44800
rect 125640 44800 125800 44960
rect 125640 44960 125800 45120
rect 125640 45120 125800 45280
rect 125640 45280 125800 45440
rect 125640 45440 125800 45600
rect 125640 45600 125800 45760
rect 125640 45760 125800 45920
rect 125640 45920 125800 46080
rect 125640 46080 125800 46240
rect 125640 46240 125800 46400
rect 125640 46400 125800 46560
rect 125640 46560 125800 46720
rect 125640 46720 125800 46880
rect 125640 46880 125800 47040
rect 125640 47040 125800 47200
rect 125640 47200 125800 47360
rect 125640 47360 125800 47520
rect 125640 47520 125800 47680
rect 125640 47680 125800 47840
rect 125640 47840 125800 48000
rect 125640 48000 125800 48160
rect 125640 48160 125800 48320
rect 125640 48320 125800 48480
rect 125640 48480 125800 48640
rect 125640 48640 125800 48800
rect 125800 29120 125960 29280
rect 125800 29280 125960 29440
rect 125800 29440 125960 29600
rect 125800 29600 125960 29760
rect 125800 29760 125960 29920
rect 125800 29920 125960 30080
rect 125800 30080 125960 30240
rect 125800 30240 125960 30400
rect 125800 30400 125960 30560
rect 125800 30560 125960 30720
rect 125800 30720 125960 30880
rect 125800 30880 125960 31040
rect 125800 31040 125960 31200
rect 125800 31200 125960 31360
rect 125800 31360 125960 31520
rect 125800 31520 125960 31680
rect 125800 31680 125960 31840
rect 125800 31840 125960 32000
rect 125800 32000 125960 32160
rect 125800 32160 125960 32320
rect 125800 32320 125960 32480
rect 125800 32480 125960 32640
rect 125800 32640 125960 32800
rect 125800 32800 125960 32960
rect 125800 32960 125960 33120
rect 125800 33120 125960 33280
rect 125800 33280 125960 33440
rect 125800 33440 125960 33600
rect 125800 33600 125960 33760
rect 125800 33760 125960 33920
rect 125800 33920 125960 34080
rect 125800 34080 125960 34240
rect 125800 34240 125960 34400
rect 125800 34400 125960 34560
rect 125800 34560 125960 34720
rect 125800 34720 125960 34880
rect 125800 34880 125960 35040
rect 125800 35040 125960 35200
rect 125800 35200 125960 35360
rect 125800 35360 125960 35520
rect 125800 35520 125960 35680
rect 125800 40640 125960 40800
rect 125800 40800 125960 40960
rect 125800 40960 125960 41120
rect 125800 41120 125960 41280
rect 125800 41280 125960 41440
rect 125800 41440 125960 41600
rect 125800 41600 125960 41760
rect 125800 41760 125960 41920
rect 125800 41920 125960 42080
rect 125800 42080 125960 42240
rect 125800 42240 125960 42400
rect 125800 42400 125960 42560
rect 125800 42560 125960 42720
rect 125800 42720 125960 42880
rect 125800 42880 125960 43040
rect 125800 43040 125960 43200
rect 125800 43200 125960 43360
rect 125800 43360 125960 43520
rect 125800 43520 125960 43680
rect 125800 43680 125960 43840
rect 125800 43840 125960 44000
rect 125800 44000 125960 44160
rect 125800 44160 125960 44320
rect 125800 44320 125960 44480
rect 125800 44480 125960 44640
rect 125800 44640 125960 44800
rect 125800 44800 125960 44960
rect 125800 44960 125960 45120
rect 125800 45120 125960 45280
rect 125800 45280 125960 45440
rect 125800 45440 125960 45600
rect 125800 45600 125960 45760
rect 125800 45760 125960 45920
rect 125800 45920 125960 46080
rect 125800 46080 125960 46240
rect 125800 46240 125960 46400
rect 125800 46400 125960 46560
rect 125800 46560 125960 46720
rect 125800 46720 125960 46880
rect 125800 46880 125960 47040
rect 125800 47040 125960 47200
rect 125800 47200 125960 47360
rect 125800 47360 125960 47520
rect 125800 47520 125960 47680
rect 125800 47680 125960 47840
rect 125800 47840 125960 48000
rect 125800 48000 125960 48160
rect 125800 48160 125960 48320
rect 125800 48320 125960 48480
rect 125800 48480 125960 48640
rect 125800 48640 125960 48800
rect 125800 48800 125960 48960
rect 125960 28960 126120 29120
rect 125960 29120 126120 29280
rect 125960 29280 126120 29440
rect 125960 29440 126120 29600
rect 125960 29600 126120 29760
rect 125960 29760 126120 29920
rect 125960 29920 126120 30080
rect 125960 30080 126120 30240
rect 125960 30240 126120 30400
rect 125960 30400 126120 30560
rect 125960 30560 126120 30720
rect 125960 30720 126120 30880
rect 125960 30880 126120 31040
rect 125960 31040 126120 31200
rect 125960 31200 126120 31360
rect 125960 31360 126120 31520
rect 125960 31520 126120 31680
rect 125960 31680 126120 31840
rect 125960 31840 126120 32000
rect 125960 32000 126120 32160
rect 125960 32160 126120 32320
rect 125960 32320 126120 32480
rect 125960 32480 126120 32640
rect 125960 32640 126120 32800
rect 125960 32800 126120 32960
rect 125960 32960 126120 33120
rect 125960 33120 126120 33280
rect 125960 33280 126120 33440
rect 125960 33440 126120 33600
rect 125960 33600 126120 33760
rect 125960 33760 126120 33920
rect 125960 33920 126120 34080
rect 125960 34080 126120 34240
rect 125960 34240 126120 34400
rect 125960 34400 126120 34560
rect 125960 34560 126120 34720
rect 125960 34720 126120 34880
rect 125960 41440 126120 41600
rect 125960 41600 126120 41760
rect 125960 41760 126120 41920
rect 125960 41920 126120 42080
rect 125960 42080 126120 42240
rect 125960 42240 126120 42400
rect 125960 42400 126120 42560
rect 125960 42560 126120 42720
rect 125960 42720 126120 42880
rect 125960 42880 126120 43040
rect 125960 43040 126120 43200
rect 125960 43200 126120 43360
rect 125960 43360 126120 43520
rect 125960 43520 126120 43680
rect 125960 43680 126120 43840
rect 125960 43840 126120 44000
rect 125960 44000 126120 44160
rect 125960 44160 126120 44320
rect 125960 44320 126120 44480
rect 125960 44480 126120 44640
rect 125960 44640 126120 44800
rect 125960 44800 126120 44960
rect 125960 44960 126120 45120
rect 125960 45120 126120 45280
rect 125960 45280 126120 45440
rect 125960 45440 126120 45600
rect 125960 45600 126120 45760
rect 125960 45760 126120 45920
rect 125960 45920 126120 46080
rect 125960 46080 126120 46240
rect 125960 46240 126120 46400
rect 125960 46400 126120 46560
rect 125960 46560 126120 46720
rect 125960 46720 126120 46880
rect 125960 46880 126120 47040
rect 125960 47040 126120 47200
rect 125960 47200 126120 47360
rect 125960 47360 126120 47520
rect 125960 47520 126120 47680
rect 125960 47680 126120 47840
rect 125960 47840 126120 48000
rect 125960 48000 126120 48160
rect 125960 48160 126120 48320
rect 125960 48320 126120 48480
rect 125960 48480 126120 48640
rect 125960 48640 126120 48800
rect 125960 48800 126120 48960
rect 125960 48960 126120 49120
rect 125960 49120 126120 49280
rect 126120 28800 126280 28960
rect 126120 28960 126280 29120
rect 126120 29120 126280 29280
rect 126120 29280 126280 29440
rect 126120 29440 126280 29600
rect 126120 29600 126280 29760
rect 126120 29760 126280 29920
rect 126120 29920 126280 30080
rect 126120 30080 126280 30240
rect 126120 30240 126280 30400
rect 126120 30400 126280 30560
rect 126120 30560 126280 30720
rect 126120 30720 126280 30880
rect 126120 30880 126280 31040
rect 126120 31040 126280 31200
rect 126120 31200 126280 31360
rect 126120 31360 126280 31520
rect 126120 31520 126280 31680
rect 126120 31680 126280 31840
rect 126120 31840 126280 32000
rect 126120 32000 126280 32160
rect 126120 32160 126280 32320
rect 126120 32320 126280 32480
rect 126120 32480 126280 32640
rect 126120 32640 126280 32800
rect 126120 32800 126280 32960
rect 126120 32960 126280 33120
rect 126120 33120 126280 33280
rect 126120 33280 126280 33440
rect 126120 33440 126280 33600
rect 126120 33600 126280 33760
rect 126120 33760 126280 33920
rect 126120 33920 126280 34080
rect 126120 34080 126280 34240
rect 126120 34240 126280 34400
rect 126120 42080 126280 42240
rect 126120 42240 126280 42400
rect 126120 42400 126280 42560
rect 126120 42560 126280 42720
rect 126120 42720 126280 42880
rect 126120 42880 126280 43040
rect 126120 43040 126280 43200
rect 126120 43200 126280 43360
rect 126120 43360 126280 43520
rect 126120 43520 126280 43680
rect 126120 43680 126280 43840
rect 126120 43840 126280 44000
rect 126120 44000 126280 44160
rect 126120 44160 126280 44320
rect 126120 44320 126280 44480
rect 126120 44480 126280 44640
rect 126120 44640 126280 44800
rect 126120 44800 126280 44960
rect 126120 44960 126280 45120
rect 126120 45120 126280 45280
rect 126120 45280 126280 45440
rect 126120 45440 126280 45600
rect 126120 45600 126280 45760
rect 126120 45760 126280 45920
rect 126120 45920 126280 46080
rect 126120 46080 126280 46240
rect 126120 46240 126280 46400
rect 126120 46400 126280 46560
rect 126120 46560 126280 46720
rect 126120 46720 126280 46880
rect 126120 46880 126280 47040
rect 126120 47040 126280 47200
rect 126120 47200 126280 47360
rect 126120 47360 126280 47520
rect 126120 47520 126280 47680
rect 126120 47680 126280 47840
rect 126120 47840 126280 48000
rect 126120 48000 126280 48160
rect 126120 48160 126280 48320
rect 126120 48320 126280 48480
rect 126120 48480 126280 48640
rect 126120 48640 126280 48800
rect 126120 48800 126280 48960
rect 126120 48960 126280 49120
rect 126120 49120 126280 49280
rect 126120 49280 126280 49440
rect 126280 28800 126440 28960
rect 126280 28960 126440 29120
rect 126280 29120 126440 29280
rect 126280 29280 126440 29440
rect 126280 29440 126440 29600
rect 126280 29600 126440 29760
rect 126280 29760 126440 29920
rect 126280 29920 126440 30080
rect 126280 30080 126440 30240
rect 126280 30240 126440 30400
rect 126280 30400 126440 30560
rect 126280 30560 126440 30720
rect 126280 30720 126440 30880
rect 126280 30880 126440 31040
rect 126280 31040 126440 31200
rect 126280 31200 126440 31360
rect 126280 31360 126440 31520
rect 126280 31520 126440 31680
rect 126280 31680 126440 31840
rect 126280 31840 126440 32000
rect 126280 32000 126440 32160
rect 126280 32160 126440 32320
rect 126280 32320 126440 32480
rect 126280 32480 126440 32640
rect 126280 32640 126440 32800
rect 126280 32800 126440 32960
rect 126280 32960 126440 33120
rect 126280 33120 126440 33280
rect 126280 33280 126440 33440
rect 126280 33440 126440 33600
rect 126280 33600 126440 33760
rect 126280 33760 126440 33920
rect 126280 33920 126440 34080
rect 126280 42720 126440 42880
rect 126280 42880 126440 43040
rect 126280 43040 126440 43200
rect 126280 43200 126440 43360
rect 126280 43360 126440 43520
rect 126280 43520 126440 43680
rect 126280 43680 126440 43840
rect 126280 43840 126440 44000
rect 126280 44000 126440 44160
rect 126280 44160 126440 44320
rect 126280 44320 126440 44480
rect 126280 44480 126440 44640
rect 126280 44640 126440 44800
rect 126280 44800 126440 44960
rect 126280 44960 126440 45120
rect 126280 45120 126440 45280
rect 126280 45280 126440 45440
rect 126280 45440 126440 45600
rect 126280 45600 126440 45760
rect 126280 45760 126440 45920
rect 126280 45920 126440 46080
rect 126280 46080 126440 46240
rect 126280 46240 126440 46400
rect 126280 46400 126440 46560
rect 126280 46560 126440 46720
rect 126280 46720 126440 46880
rect 126280 46880 126440 47040
rect 126280 47040 126440 47200
rect 126280 47200 126440 47360
rect 126280 47360 126440 47520
rect 126280 47520 126440 47680
rect 126280 47680 126440 47840
rect 126280 47840 126440 48000
rect 126280 48000 126440 48160
rect 126280 48160 126440 48320
rect 126280 48320 126440 48480
rect 126280 48480 126440 48640
rect 126280 48640 126440 48800
rect 126280 48800 126440 48960
rect 126280 48960 126440 49120
rect 126280 49120 126440 49280
rect 126280 49280 126440 49440
rect 126280 49440 126440 49600
rect 126440 28640 126600 28800
rect 126440 28800 126600 28960
rect 126440 28960 126600 29120
rect 126440 29120 126600 29280
rect 126440 29280 126600 29440
rect 126440 29440 126600 29600
rect 126440 29600 126600 29760
rect 126440 29760 126600 29920
rect 126440 29920 126600 30080
rect 126440 30080 126600 30240
rect 126440 30240 126600 30400
rect 126440 30400 126600 30560
rect 126440 30560 126600 30720
rect 126440 30720 126600 30880
rect 126440 30880 126600 31040
rect 126440 31040 126600 31200
rect 126440 31200 126600 31360
rect 126440 31360 126600 31520
rect 126440 31520 126600 31680
rect 126440 31680 126600 31840
rect 126440 31840 126600 32000
rect 126440 32000 126600 32160
rect 126440 32160 126600 32320
rect 126440 32320 126600 32480
rect 126440 32480 126600 32640
rect 126440 32640 126600 32800
rect 126440 32800 126600 32960
rect 126440 32960 126600 33120
rect 126440 33120 126600 33280
rect 126440 33280 126600 33440
rect 126440 33440 126600 33600
rect 126440 43040 126600 43200
rect 126440 43200 126600 43360
rect 126440 43360 126600 43520
rect 126440 43520 126600 43680
rect 126440 43680 126600 43840
rect 126440 43840 126600 44000
rect 126440 44000 126600 44160
rect 126440 44160 126600 44320
rect 126440 44320 126600 44480
rect 126440 44480 126600 44640
rect 126440 44640 126600 44800
rect 126440 44800 126600 44960
rect 126440 44960 126600 45120
rect 126440 45120 126600 45280
rect 126440 45280 126600 45440
rect 126440 45440 126600 45600
rect 126440 45600 126600 45760
rect 126440 45760 126600 45920
rect 126440 45920 126600 46080
rect 126440 46080 126600 46240
rect 126440 46240 126600 46400
rect 126440 46400 126600 46560
rect 126440 46560 126600 46720
rect 126440 46720 126600 46880
rect 126440 46880 126600 47040
rect 126440 47040 126600 47200
rect 126440 47200 126600 47360
rect 126440 47360 126600 47520
rect 126440 47520 126600 47680
rect 126440 47680 126600 47840
rect 126440 47840 126600 48000
rect 126440 48000 126600 48160
rect 126440 48160 126600 48320
rect 126440 48320 126600 48480
rect 126440 48480 126600 48640
rect 126440 48640 126600 48800
rect 126440 48800 126600 48960
rect 126440 48960 126600 49120
rect 126440 49120 126600 49280
rect 126440 49280 126600 49440
rect 126440 49440 126600 49600
rect 126440 49600 126600 49760
rect 126600 28480 126760 28640
rect 126600 28640 126760 28800
rect 126600 28800 126760 28960
rect 126600 28960 126760 29120
rect 126600 29120 126760 29280
rect 126600 29280 126760 29440
rect 126600 29440 126760 29600
rect 126600 29600 126760 29760
rect 126600 29760 126760 29920
rect 126600 29920 126760 30080
rect 126600 30080 126760 30240
rect 126600 30240 126760 30400
rect 126600 30400 126760 30560
rect 126600 30560 126760 30720
rect 126600 30720 126760 30880
rect 126600 30880 126760 31040
rect 126600 31040 126760 31200
rect 126600 31200 126760 31360
rect 126600 31360 126760 31520
rect 126600 31520 126760 31680
rect 126600 31680 126760 31840
rect 126600 31840 126760 32000
rect 126600 32000 126760 32160
rect 126600 32160 126760 32320
rect 126600 32320 126760 32480
rect 126600 32480 126760 32640
rect 126600 32640 126760 32800
rect 126600 32800 126760 32960
rect 126600 32960 126760 33120
rect 126600 33120 126760 33280
rect 126600 33280 126760 33440
rect 126600 43520 126760 43680
rect 126600 43680 126760 43840
rect 126600 43840 126760 44000
rect 126600 44000 126760 44160
rect 126600 44160 126760 44320
rect 126600 44320 126760 44480
rect 126600 44480 126760 44640
rect 126600 44640 126760 44800
rect 126600 44800 126760 44960
rect 126600 44960 126760 45120
rect 126600 45120 126760 45280
rect 126600 45280 126760 45440
rect 126600 45440 126760 45600
rect 126600 45600 126760 45760
rect 126600 45760 126760 45920
rect 126600 45920 126760 46080
rect 126600 46080 126760 46240
rect 126600 46240 126760 46400
rect 126600 46400 126760 46560
rect 126600 46560 126760 46720
rect 126600 46720 126760 46880
rect 126600 46880 126760 47040
rect 126600 47040 126760 47200
rect 126600 47200 126760 47360
rect 126600 47360 126760 47520
rect 126600 47520 126760 47680
rect 126600 47680 126760 47840
rect 126600 47840 126760 48000
rect 126600 48000 126760 48160
rect 126600 48160 126760 48320
rect 126600 48320 126760 48480
rect 126600 48480 126760 48640
rect 126600 48640 126760 48800
rect 126600 48800 126760 48960
rect 126600 48960 126760 49120
rect 126600 49120 126760 49280
rect 126600 49280 126760 49440
rect 126600 49440 126760 49600
rect 126600 49600 126760 49760
rect 126600 49760 126760 49920
rect 126760 28320 126920 28480
rect 126760 28480 126920 28640
rect 126760 28640 126920 28800
rect 126760 28800 126920 28960
rect 126760 28960 126920 29120
rect 126760 29120 126920 29280
rect 126760 29280 126920 29440
rect 126760 29440 126920 29600
rect 126760 29600 126920 29760
rect 126760 29760 126920 29920
rect 126760 29920 126920 30080
rect 126760 30080 126920 30240
rect 126760 30240 126920 30400
rect 126760 30400 126920 30560
rect 126760 30560 126920 30720
rect 126760 30720 126920 30880
rect 126760 30880 126920 31040
rect 126760 31040 126920 31200
rect 126760 31200 126920 31360
rect 126760 31360 126920 31520
rect 126760 31520 126920 31680
rect 126760 31680 126920 31840
rect 126760 31840 126920 32000
rect 126760 32000 126920 32160
rect 126760 32160 126920 32320
rect 126760 32320 126920 32480
rect 126760 32480 126920 32640
rect 126760 32640 126920 32800
rect 126760 32800 126920 32960
rect 126760 32960 126920 33120
rect 126760 44000 126920 44160
rect 126760 44160 126920 44320
rect 126760 44320 126920 44480
rect 126760 44480 126920 44640
rect 126760 44640 126920 44800
rect 126760 44800 126920 44960
rect 126760 44960 126920 45120
rect 126760 45120 126920 45280
rect 126760 45280 126920 45440
rect 126760 45440 126920 45600
rect 126760 45600 126920 45760
rect 126760 45760 126920 45920
rect 126760 45920 126920 46080
rect 126760 46080 126920 46240
rect 126760 46240 126920 46400
rect 126760 46400 126920 46560
rect 126760 46560 126920 46720
rect 126760 46720 126920 46880
rect 126760 46880 126920 47040
rect 126760 47040 126920 47200
rect 126760 47200 126920 47360
rect 126760 47360 126920 47520
rect 126760 47520 126920 47680
rect 126760 47680 126920 47840
rect 126760 47840 126920 48000
rect 126760 48000 126920 48160
rect 126760 48160 126920 48320
rect 126760 48320 126920 48480
rect 126760 48480 126920 48640
rect 126760 48640 126920 48800
rect 126760 48800 126920 48960
rect 126760 48960 126920 49120
rect 126760 49120 126920 49280
rect 126760 49280 126920 49440
rect 126760 49440 126920 49600
rect 126760 49600 126920 49760
rect 126760 49760 126920 49920
rect 126760 49920 126920 50080
rect 126920 28320 127080 28480
rect 126920 28480 127080 28640
rect 126920 28640 127080 28800
rect 126920 28800 127080 28960
rect 126920 28960 127080 29120
rect 126920 29120 127080 29280
rect 126920 29280 127080 29440
rect 126920 29440 127080 29600
rect 126920 29600 127080 29760
rect 126920 29760 127080 29920
rect 126920 29920 127080 30080
rect 126920 30080 127080 30240
rect 126920 30240 127080 30400
rect 126920 30400 127080 30560
rect 126920 30560 127080 30720
rect 126920 30720 127080 30880
rect 126920 30880 127080 31040
rect 126920 31040 127080 31200
rect 126920 31200 127080 31360
rect 126920 31360 127080 31520
rect 126920 31520 127080 31680
rect 126920 31680 127080 31840
rect 126920 31840 127080 32000
rect 126920 32000 127080 32160
rect 126920 32160 127080 32320
rect 126920 32320 127080 32480
rect 126920 32480 127080 32640
rect 126920 32640 127080 32800
rect 126920 44320 127080 44480
rect 126920 44480 127080 44640
rect 126920 44640 127080 44800
rect 126920 44800 127080 44960
rect 126920 44960 127080 45120
rect 126920 45120 127080 45280
rect 126920 45280 127080 45440
rect 126920 45440 127080 45600
rect 126920 45600 127080 45760
rect 126920 45760 127080 45920
rect 126920 45920 127080 46080
rect 126920 46080 127080 46240
rect 126920 46240 127080 46400
rect 126920 46400 127080 46560
rect 126920 46560 127080 46720
rect 126920 46720 127080 46880
rect 126920 46880 127080 47040
rect 126920 47040 127080 47200
rect 126920 47200 127080 47360
rect 126920 47360 127080 47520
rect 126920 47520 127080 47680
rect 126920 47680 127080 47840
rect 126920 47840 127080 48000
rect 126920 48000 127080 48160
rect 126920 48160 127080 48320
rect 126920 48320 127080 48480
rect 126920 48480 127080 48640
rect 126920 48640 127080 48800
rect 126920 48800 127080 48960
rect 126920 48960 127080 49120
rect 126920 49120 127080 49280
rect 126920 49280 127080 49440
rect 126920 49440 127080 49600
rect 126920 49600 127080 49760
rect 126920 49760 127080 49920
rect 126920 49920 127080 50080
rect 126920 50080 127080 50240
rect 127080 28160 127240 28320
rect 127080 28320 127240 28480
rect 127080 28480 127240 28640
rect 127080 28640 127240 28800
rect 127080 28800 127240 28960
rect 127080 28960 127240 29120
rect 127080 29120 127240 29280
rect 127080 29280 127240 29440
rect 127080 29440 127240 29600
rect 127080 29600 127240 29760
rect 127080 29760 127240 29920
rect 127080 29920 127240 30080
rect 127080 30080 127240 30240
rect 127080 30240 127240 30400
rect 127080 30400 127240 30560
rect 127080 30560 127240 30720
rect 127080 30720 127240 30880
rect 127080 30880 127240 31040
rect 127080 31040 127240 31200
rect 127080 31200 127240 31360
rect 127080 31360 127240 31520
rect 127080 31520 127240 31680
rect 127080 31680 127240 31840
rect 127080 31840 127240 32000
rect 127080 32000 127240 32160
rect 127080 32160 127240 32320
rect 127080 32320 127240 32480
rect 127080 32480 127240 32640
rect 127080 44640 127240 44800
rect 127080 44800 127240 44960
rect 127080 44960 127240 45120
rect 127080 45120 127240 45280
rect 127080 45280 127240 45440
rect 127080 45440 127240 45600
rect 127080 45600 127240 45760
rect 127080 45760 127240 45920
rect 127080 45920 127240 46080
rect 127080 46080 127240 46240
rect 127080 46240 127240 46400
rect 127080 46400 127240 46560
rect 127080 46560 127240 46720
rect 127080 46720 127240 46880
rect 127080 46880 127240 47040
rect 127080 47040 127240 47200
rect 127080 47200 127240 47360
rect 127080 47360 127240 47520
rect 127080 47520 127240 47680
rect 127080 47680 127240 47840
rect 127080 47840 127240 48000
rect 127080 48000 127240 48160
rect 127080 48160 127240 48320
rect 127080 48320 127240 48480
rect 127080 48480 127240 48640
rect 127080 48640 127240 48800
rect 127080 48800 127240 48960
rect 127080 48960 127240 49120
rect 127080 49120 127240 49280
rect 127080 49280 127240 49440
rect 127080 49440 127240 49600
rect 127080 49600 127240 49760
rect 127080 49760 127240 49920
rect 127080 49920 127240 50080
rect 127080 50080 127240 50240
rect 127080 50240 127240 50400
rect 127240 28000 127400 28160
rect 127240 28160 127400 28320
rect 127240 28320 127400 28480
rect 127240 28480 127400 28640
rect 127240 28640 127400 28800
rect 127240 28800 127400 28960
rect 127240 28960 127400 29120
rect 127240 29120 127400 29280
rect 127240 29280 127400 29440
rect 127240 29440 127400 29600
rect 127240 29600 127400 29760
rect 127240 29760 127400 29920
rect 127240 29920 127400 30080
rect 127240 30080 127400 30240
rect 127240 30240 127400 30400
rect 127240 30400 127400 30560
rect 127240 30560 127400 30720
rect 127240 30720 127400 30880
rect 127240 30880 127400 31040
rect 127240 31040 127400 31200
rect 127240 31200 127400 31360
rect 127240 31360 127400 31520
rect 127240 31520 127400 31680
rect 127240 31680 127400 31840
rect 127240 31840 127400 32000
rect 127240 32000 127400 32160
rect 127240 32160 127400 32320
rect 127240 32320 127400 32480
rect 127240 44960 127400 45120
rect 127240 45120 127400 45280
rect 127240 45280 127400 45440
rect 127240 45440 127400 45600
rect 127240 45600 127400 45760
rect 127240 45760 127400 45920
rect 127240 45920 127400 46080
rect 127240 46080 127400 46240
rect 127240 46240 127400 46400
rect 127240 46400 127400 46560
rect 127240 46560 127400 46720
rect 127240 46720 127400 46880
rect 127240 46880 127400 47040
rect 127240 47040 127400 47200
rect 127240 47200 127400 47360
rect 127240 47360 127400 47520
rect 127240 47520 127400 47680
rect 127240 47680 127400 47840
rect 127240 47840 127400 48000
rect 127240 48000 127400 48160
rect 127240 48160 127400 48320
rect 127240 48320 127400 48480
rect 127240 48480 127400 48640
rect 127240 48640 127400 48800
rect 127240 48800 127400 48960
rect 127240 48960 127400 49120
rect 127240 49120 127400 49280
rect 127240 49280 127400 49440
rect 127240 49440 127400 49600
rect 127240 49600 127400 49760
rect 127240 49760 127400 49920
rect 127240 49920 127400 50080
rect 127240 50080 127400 50240
rect 127240 50240 127400 50400
rect 127240 50400 127400 50560
rect 127400 28000 127560 28160
rect 127400 28160 127560 28320
rect 127400 28320 127560 28480
rect 127400 28480 127560 28640
rect 127400 28640 127560 28800
rect 127400 28800 127560 28960
rect 127400 28960 127560 29120
rect 127400 29120 127560 29280
rect 127400 29280 127560 29440
rect 127400 29440 127560 29600
rect 127400 29600 127560 29760
rect 127400 29760 127560 29920
rect 127400 29920 127560 30080
rect 127400 30080 127560 30240
rect 127400 30240 127560 30400
rect 127400 30400 127560 30560
rect 127400 30560 127560 30720
rect 127400 30720 127560 30880
rect 127400 30880 127560 31040
rect 127400 31040 127560 31200
rect 127400 31200 127560 31360
rect 127400 31360 127560 31520
rect 127400 31520 127560 31680
rect 127400 31680 127560 31840
rect 127400 31840 127560 32000
rect 127400 32000 127560 32160
rect 127400 32160 127560 32320
rect 127400 45280 127560 45440
rect 127400 45440 127560 45600
rect 127400 45600 127560 45760
rect 127400 45760 127560 45920
rect 127400 45920 127560 46080
rect 127400 46080 127560 46240
rect 127400 46240 127560 46400
rect 127400 46400 127560 46560
rect 127400 46560 127560 46720
rect 127400 46720 127560 46880
rect 127400 46880 127560 47040
rect 127400 47040 127560 47200
rect 127400 47200 127560 47360
rect 127400 47360 127560 47520
rect 127400 47520 127560 47680
rect 127400 47680 127560 47840
rect 127400 47840 127560 48000
rect 127400 48000 127560 48160
rect 127400 48160 127560 48320
rect 127400 48320 127560 48480
rect 127400 48480 127560 48640
rect 127400 48640 127560 48800
rect 127400 48800 127560 48960
rect 127400 48960 127560 49120
rect 127400 49120 127560 49280
rect 127400 49280 127560 49440
rect 127400 49440 127560 49600
rect 127400 49600 127560 49760
rect 127400 49760 127560 49920
rect 127400 49920 127560 50080
rect 127400 50080 127560 50240
rect 127400 50240 127560 50400
rect 127400 50400 127560 50560
rect 127400 50560 127560 50720
rect 127560 27840 127720 28000
rect 127560 28000 127720 28160
rect 127560 28160 127720 28320
rect 127560 28320 127720 28480
rect 127560 28480 127720 28640
rect 127560 28640 127720 28800
rect 127560 28800 127720 28960
rect 127560 28960 127720 29120
rect 127560 29120 127720 29280
rect 127560 29280 127720 29440
rect 127560 29440 127720 29600
rect 127560 29600 127720 29760
rect 127560 29760 127720 29920
rect 127560 29920 127720 30080
rect 127560 30080 127720 30240
rect 127560 30240 127720 30400
rect 127560 30400 127720 30560
rect 127560 30560 127720 30720
rect 127560 30720 127720 30880
rect 127560 30880 127720 31040
rect 127560 31040 127720 31200
rect 127560 31200 127720 31360
rect 127560 31360 127720 31520
rect 127560 31520 127720 31680
rect 127560 31680 127720 31840
rect 127560 31840 127720 32000
rect 127560 32000 127720 32160
rect 127560 45600 127720 45760
rect 127560 45760 127720 45920
rect 127560 45920 127720 46080
rect 127560 46080 127720 46240
rect 127560 46240 127720 46400
rect 127560 46400 127720 46560
rect 127560 46560 127720 46720
rect 127560 46720 127720 46880
rect 127560 46880 127720 47040
rect 127560 47040 127720 47200
rect 127560 47200 127720 47360
rect 127560 47360 127720 47520
rect 127560 47520 127720 47680
rect 127560 47680 127720 47840
rect 127560 47840 127720 48000
rect 127560 48000 127720 48160
rect 127560 48160 127720 48320
rect 127560 48320 127720 48480
rect 127560 48480 127720 48640
rect 127560 48640 127720 48800
rect 127560 48800 127720 48960
rect 127560 48960 127720 49120
rect 127560 49120 127720 49280
rect 127560 49280 127720 49440
rect 127560 49440 127720 49600
rect 127560 49600 127720 49760
rect 127560 49760 127720 49920
rect 127560 49920 127720 50080
rect 127560 50080 127720 50240
rect 127560 50240 127720 50400
rect 127560 50400 127720 50560
rect 127560 50560 127720 50720
rect 127560 50720 127720 50880
rect 127720 27840 127880 28000
rect 127720 28000 127880 28160
rect 127720 28160 127880 28320
rect 127720 28320 127880 28480
rect 127720 28480 127880 28640
rect 127720 28640 127880 28800
rect 127720 28800 127880 28960
rect 127720 28960 127880 29120
rect 127720 29120 127880 29280
rect 127720 29280 127880 29440
rect 127720 29440 127880 29600
rect 127720 29600 127880 29760
rect 127720 29760 127880 29920
rect 127720 29920 127880 30080
rect 127720 30080 127880 30240
rect 127720 30240 127880 30400
rect 127720 30400 127880 30560
rect 127720 30560 127880 30720
rect 127720 30720 127880 30880
rect 127720 30880 127880 31040
rect 127720 31040 127880 31200
rect 127720 31200 127880 31360
rect 127720 31360 127880 31520
rect 127720 31520 127880 31680
rect 127720 31680 127880 31840
rect 127720 31840 127880 32000
rect 127720 45920 127880 46080
rect 127720 46080 127880 46240
rect 127720 46240 127880 46400
rect 127720 46400 127880 46560
rect 127720 46560 127880 46720
rect 127720 46720 127880 46880
rect 127720 46880 127880 47040
rect 127720 47040 127880 47200
rect 127720 47200 127880 47360
rect 127720 47360 127880 47520
rect 127720 47520 127880 47680
rect 127720 47680 127880 47840
rect 127720 47840 127880 48000
rect 127720 48000 127880 48160
rect 127720 48160 127880 48320
rect 127720 48320 127880 48480
rect 127720 48480 127880 48640
rect 127720 48640 127880 48800
rect 127720 48800 127880 48960
rect 127720 48960 127880 49120
rect 127720 49120 127880 49280
rect 127720 49280 127880 49440
rect 127720 49440 127880 49600
rect 127720 49600 127880 49760
rect 127720 49760 127880 49920
rect 127720 49920 127880 50080
rect 127720 50080 127880 50240
rect 127720 50240 127880 50400
rect 127720 50400 127880 50560
rect 127720 50560 127880 50720
rect 127720 50720 127880 50880
rect 127720 50880 127880 51040
rect 127880 27680 128040 27840
rect 127880 27840 128040 28000
rect 127880 28000 128040 28160
rect 127880 28160 128040 28320
rect 127880 28320 128040 28480
rect 127880 28480 128040 28640
rect 127880 28640 128040 28800
rect 127880 28800 128040 28960
rect 127880 28960 128040 29120
rect 127880 29120 128040 29280
rect 127880 29280 128040 29440
rect 127880 29440 128040 29600
rect 127880 29600 128040 29760
rect 127880 29760 128040 29920
rect 127880 29920 128040 30080
rect 127880 30080 128040 30240
rect 127880 30240 128040 30400
rect 127880 30400 128040 30560
rect 127880 30560 128040 30720
rect 127880 30720 128040 30880
rect 127880 30880 128040 31040
rect 127880 31040 128040 31200
rect 127880 31200 128040 31360
rect 127880 31360 128040 31520
rect 127880 31520 128040 31680
rect 127880 31680 128040 31840
rect 127880 46080 128040 46240
rect 127880 46240 128040 46400
rect 127880 46400 128040 46560
rect 127880 46560 128040 46720
rect 127880 46720 128040 46880
rect 127880 46880 128040 47040
rect 127880 47040 128040 47200
rect 127880 47200 128040 47360
rect 127880 47360 128040 47520
rect 127880 47520 128040 47680
rect 127880 47680 128040 47840
rect 127880 47840 128040 48000
rect 127880 48000 128040 48160
rect 127880 48160 128040 48320
rect 127880 48320 128040 48480
rect 127880 48480 128040 48640
rect 127880 48640 128040 48800
rect 127880 48800 128040 48960
rect 127880 48960 128040 49120
rect 127880 49120 128040 49280
rect 127880 49280 128040 49440
rect 127880 49440 128040 49600
rect 127880 49600 128040 49760
rect 127880 49760 128040 49920
rect 127880 49920 128040 50080
rect 127880 50080 128040 50240
rect 127880 50240 128040 50400
rect 127880 50400 128040 50560
rect 127880 50560 128040 50720
rect 127880 50720 128040 50880
rect 127880 50880 128040 51040
rect 127880 51040 128040 51200
rect 128040 27680 128200 27840
rect 128040 27840 128200 28000
rect 128040 28000 128200 28160
rect 128040 28160 128200 28320
rect 128040 28320 128200 28480
rect 128040 28480 128200 28640
rect 128040 28640 128200 28800
rect 128040 28800 128200 28960
rect 128040 28960 128200 29120
rect 128040 29120 128200 29280
rect 128040 29280 128200 29440
rect 128040 29440 128200 29600
rect 128040 29600 128200 29760
rect 128040 29760 128200 29920
rect 128040 29920 128200 30080
rect 128040 30080 128200 30240
rect 128040 30240 128200 30400
rect 128040 30400 128200 30560
rect 128040 30560 128200 30720
rect 128040 30720 128200 30880
rect 128040 30880 128200 31040
rect 128040 31040 128200 31200
rect 128040 31200 128200 31360
rect 128040 31360 128200 31520
rect 128040 31520 128200 31680
rect 128040 46400 128200 46560
rect 128040 46560 128200 46720
rect 128040 46720 128200 46880
rect 128040 46880 128200 47040
rect 128040 47040 128200 47200
rect 128040 47200 128200 47360
rect 128040 47360 128200 47520
rect 128040 47520 128200 47680
rect 128040 47680 128200 47840
rect 128040 47840 128200 48000
rect 128040 48000 128200 48160
rect 128040 48160 128200 48320
rect 128040 48320 128200 48480
rect 128040 48480 128200 48640
rect 128040 48640 128200 48800
rect 128040 48800 128200 48960
rect 128040 48960 128200 49120
rect 128040 49120 128200 49280
rect 128040 49280 128200 49440
rect 128040 49440 128200 49600
rect 128040 49600 128200 49760
rect 128040 49760 128200 49920
rect 128040 49920 128200 50080
rect 128040 50080 128200 50240
rect 128040 50240 128200 50400
rect 128040 50400 128200 50560
rect 128040 50560 128200 50720
rect 128040 50720 128200 50880
rect 128040 50880 128200 51040
rect 128040 51040 128200 51200
rect 128200 27520 128360 27680
rect 128200 27680 128360 27840
rect 128200 27840 128360 28000
rect 128200 28000 128360 28160
rect 128200 28160 128360 28320
rect 128200 28320 128360 28480
rect 128200 28480 128360 28640
rect 128200 28640 128360 28800
rect 128200 28800 128360 28960
rect 128200 28960 128360 29120
rect 128200 29120 128360 29280
rect 128200 29280 128360 29440
rect 128200 29440 128360 29600
rect 128200 29600 128360 29760
rect 128200 29760 128360 29920
rect 128200 29920 128360 30080
rect 128200 30080 128360 30240
rect 128200 30240 128360 30400
rect 128200 30400 128360 30560
rect 128200 30560 128360 30720
rect 128200 30720 128360 30880
rect 128200 30880 128360 31040
rect 128200 31040 128360 31200
rect 128200 31200 128360 31360
rect 128200 31360 128360 31520
rect 128200 46560 128360 46720
rect 128200 46720 128360 46880
rect 128200 46880 128360 47040
rect 128200 47040 128360 47200
rect 128200 47200 128360 47360
rect 128200 47360 128360 47520
rect 128200 47520 128360 47680
rect 128200 47680 128360 47840
rect 128200 47840 128360 48000
rect 128200 48000 128360 48160
rect 128200 48160 128360 48320
rect 128200 48320 128360 48480
rect 128200 48480 128360 48640
rect 128200 48640 128360 48800
rect 128200 48800 128360 48960
rect 128200 48960 128360 49120
rect 128200 49120 128360 49280
rect 128200 49280 128360 49440
rect 128200 49440 128360 49600
rect 128200 49600 128360 49760
rect 128200 49760 128360 49920
rect 128200 49920 128360 50080
rect 128200 50080 128360 50240
rect 128200 50240 128360 50400
rect 128200 50400 128360 50560
rect 128200 50560 128360 50720
rect 128200 50720 128360 50880
rect 128200 50880 128360 51040
rect 128200 51040 128360 51200
rect 128200 51200 128360 51360
rect 128360 27520 128520 27680
rect 128360 27680 128520 27840
rect 128360 27840 128520 28000
rect 128360 28000 128520 28160
rect 128360 28160 128520 28320
rect 128360 28320 128520 28480
rect 128360 28480 128520 28640
rect 128360 28640 128520 28800
rect 128360 28800 128520 28960
rect 128360 28960 128520 29120
rect 128360 29120 128520 29280
rect 128360 29280 128520 29440
rect 128360 29440 128520 29600
rect 128360 29600 128520 29760
rect 128360 29760 128520 29920
rect 128360 29920 128520 30080
rect 128360 30080 128520 30240
rect 128360 30240 128520 30400
rect 128360 30400 128520 30560
rect 128360 30560 128520 30720
rect 128360 30720 128520 30880
rect 128360 30880 128520 31040
rect 128360 31040 128520 31200
rect 128360 31200 128520 31360
rect 128360 46880 128520 47040
rect 128360 47040 128520 47200
rect 128360 47200 128520 47360
rect 128360 47360 128520 47520
rect 128360 47520 128520 47680
rect 128360 47680 128520 47840
rect 128360 47840 128520 48000
rect 128360 48000 128520 48160
rect 128360 48160 128520 48320
rect 128360 48320 128520 48480
rect 128360 48480 128520 48640
rect 128360 48640 128520 48800
rect 128360 48800 128520 48960
rect 128360 48960 128520 49120
rect 128360 49120 128520 49280
rect 128360 49280 128520 49440
rect 128360 49440 128520 49600
rect 128360 49600 128520 49760
rect 128360 49760 128520 49920
rect 128360 49920 128520 50080
rect 128360 50080 128520 50240
rect 128360 50240 128520 50400
rect 128360 50400 128520 50560
rect 128360 50560 128520 50720
rect 128360 50720 128520 50880
rect 128360 50880 128520 51040
rect 128360 51040 128520 51200
rect 128360 51200 128520 51360
rect 128360 51360 128520 51520
rect 128520 27360 128680 27520
rect 128520 27520 128680 27680
rect 128520 27680 128680 27840
rect 128520 27840 128680 28000
rect 128520 28000 128680 28160
rect 128520 28160 128680 28320
rect 128520 28320 128680 28480
rect 128520 28480 128680 28640
rect 128520 28640 128680 28800
rect 128520 28800 128680 28960
rect 128520 28960 128680 29120
rect 128520 29120 128680 29280
rect 128520 29280 128680 29440
rect 128520 29440 128680 29600
rect 128520 29600 128680 29760
rect 128520 29760 128680 29920
rect 128520 29920 128680 30080
rect 128520 30080 128680 30240
rect 128520 30240 128680 30400
rect 128520 30400 128680 30560
rect 128520 30560 128680 30720
rect 128520 30720 128680 30880
rect 128520 30880 128680 31040
rect 128520 31040 128680 31200
rect 128520 31200 128680 31360
rect 128520 47040 128680 47200
rect 128520 47200 128680 47360
rect 128520 47360 128680 47520
rect 128520 47520 128680 47680
rect 128520 47680 128680 47840
rect 128520 47840 128680 48000
rect 128520 48000 128680 48160
rect 128520 48160 128680 48320
rect 128520 48320 128680 48480
rect 128520 48480 128680 48640
rect 128520 48640 128680 48800
rect 128520 48800 128680 48960
rect 128520 48960 128680 49120
rect 128520 49120 128680 49280
rect 128520 49280 128680 49440
rect 128520 49440 128680 49600
rect 128520 49600 128680 49760
rect 128520 49760 128680 49920
rect 128520 49920 128680 50080
rect 128520 50080 128680 50240
rect 128520 50240 128680 50400
rect 128520 50400 128680 50560
rect 128520 50560 128680 50720
rect 128520 50720 128680 50880
rect 128520 50880 128680 51040
rect 128520 51040 128680 51200
rect 128520 51200 128680 51360
rect 128520 51360 128680 51520
rect 128520 51520 128680 51680
rect 128680 27360 128840 27520
rect 128680 27520 128840 27680
rect 128680 27680 128840 27840
rect 128680 27840 128840 28000
rect 128680 28000 128840 28160
rect 128680 28160 128840 28320
rect 128680 28320 128840 28480
rect 128680 28480 128840 28640
rect 128680 28640 128840 28800
rect 128680 28800 128840 28960
rect 128680 28960 128840 29120
rect 128680 29120 128840 29280
rect 128680 29280 128840 29440
rect 128680 29440 128840 29600
rect 128680 29600 128840 29760
rect 128680 29760 128840 29920
rect 128680 29920 128840 30080
rect 128680 30080 128840 30240
rect 128680 30240 128840 30400
rect 128680 30400 128840 30560
rect 128680 30560 128840 30720
rect 128680 30720 128840 30880
rect 128680 30880 128840 31040
rect 128680 31040 128840 31200
rect 128680 47200 128840 47360
rect 128680 47360 128840 47520
rect 128680 47520 128840 47680
rect 128680 47680 128840 47840
rect 128680 47840 128840 48000
rect 128680 48000 128840 48160
rect 128680 48160 128840 48320
rect 128680 48320 128840 48480
rect 128680 48480 128840 48640
rect 128680 48640 128840 48800
rect 128680 48800 128840 48960
rect 128680 48960 128840 49120
rect 128680 49120 128840 49280
rect 128680 49280 128840 49440
rect 128680 49440 128840 49600
rect 128680 49600 128840 49760
rect 128680 49760 128840 49920
rect 128680 49920 128840 50080
rect 128680 50080 128840 50240
rect 128680 50240 128840 50400
rect 128680 50400 128840 50560
rect 128680 50560 128840 50720
rect 128680 50720 128840 50880
rect 128680 50880 128840 51040
rect 128680 51040 128840 51200
rect 128680 51200 128840 51360
rect 128680 51360 128840 51520
rect 128680 51520 128840 51680
rect 128840 27200 129000 27360
rect 128840 27360 129000 27520
rect 128840 27520 129000 27680
rect 128840 27680 129000 27840
rect 128840 27840 129000 28000
rect 128840 28000 129000 28160
rect 128840 28160 129000 28320
rect 128840 28320 129000 28480
rect 128840 28480 129000 28640
rect 128840 28640 129000 28800
rect 128840 28800 129000 28960
rect 128840 28960 129000 29120
rect 128840 29120 129000 29280
rect 128840 29280 129000 29440
rect 128840 29440 129000 29600
rect 128840 29600 129000 29760
rect 128840 29760 129000 29920
rect 128840 29920 129000 30080
rect 128840 30080 129000 30240
rect 128840 30240 129000 30400
rect 128840 30400 129000 30560
rect 128840 30560 129000 30720
rect 128840 30720 129000 30880
rect 128840 30880 129000 31040
rect 128840 47360 129000 47520
rect 128840 47520 129000 47680
rect 128840 47680 129000 47840
rect 128840 47840 129000 48000
rect 128840 48000 129000 48160
rect 128840 48160 129000 48320
rect 128840 48320 129000 48480
rect 128840 48480 129000 48640
rect 128840 48640 129000 48800
rect 128840 48800 129000 48960
rect 128840 48960 129000 49120
rect 128840 49120 129000 49280
rect 128840 49280 129000 49440
rect 128840 49440 129000 49600
rect 128840 49600 129000 49760
rect 128840 49760 129000 49920
rect 128840 49920 129000 50080
rect 128840 50080 129000 50240
rect 128840 50240 129000 50400
rect 128840 50400 129000 50560
rect 128840 50560 129000 50720
rect 128840 50720 129000 50880
rect 128840 50880 129000 51040
rect 128840 51040 129000 51200
rect 128840 51200 129000 51360
rect 128840 51360 129000 51520
rect 128840 51520 129000 51680
rect 128840 51680 129000 51840
rect 129000 27200 129160 27360
rect 129000 27360 129160 27520
rect 129000 27520 129160 27680
rect 129000 27680 129160 27840
rect 129000 27840 129160 28000
rect 129000 28000 129160 28160
rect 129000 28160 129160 28320
rect 129000 28320 129160 28480
rect 129000 28480 129160 28640
rect 129000 28640 129160 28800
rect 129000 28800 129160 28960
rect 129000 28960 129160 29120
rect 129000 29120 129160 29280
rect 129000 29280 129160 29440
rect 129000 29440 129160 29600
rect 129000 29600 129160 29760
rect 129000 29760 129160 29920
rect 129000 29920 129160 30080
rect 129000 30080 129160 30240
rect 129000 30240 129160 30400
rect 129000 30400 129160 30560
rect 129000 30560 129160 30720
rect 129000 30720 129160 30880
rect 129000 30880 129160 31040
rect 129000 47680 129160 47840
rect 129000 47840 129160 48000
rect 129000 48000 129160 48160
rect 129000 48160 129160 48320
rect 129000 48320 129160 48480
rect 129000 48480 129160 48640
rect 129000 48640 129160 48800
rect 129000 48800 129160 48960
rect 129000 48960 129160 49120
rect 129000 49120 129160 49280
rect 129000 49280 129160 49440
rect 129000 49440 129160 49600
rect 129000 49600 129160 49760
rect 129000 49760 129160 49920
rect 129000 49920 129160 50080
rect 129000 50080 129160 50240
rect 129000 50240 129160 50400
rect 129000 50400 129160 50560
rect 129000 50560 129160 50720
rect 129000 50720 129160 50880
rect 129000 50880 129160 51040
rect 129000 51040 129160 51200
rect 129000 51200 129160 51360
rect 129000 51360 129160 51520
rect 129000 51520 129160 51680
rect 129000 51680 129160 51840
rect 129160 27200 129320 27360
rect 129160 27360 129320 27520
rect 129160 27520 129320 27680
rect 129160 27680 129320 27840
rect 129160 27840 129320 28000
rect 129160 28000 129320 28160
rect 129160 28160 129320 28320
rect 129160 28320 129320 28480
rect 129160 28480 129320 28640
rect 129160 28640 129320 28800
rect 129160 28800 129320 28960
rect 129160 28960 129320 29120
rect 129160 29120 129320 29280
rect 129160 29280 129320 29440
rect 129160 29440 129320 29600
rect 129160 29600 129320 29760
rect 129160 29760 129320 29920
rect 129160 29920 129320 30080
rect 129160 30080 129320 30240
rect 129160 30240 129320 30400
rect 129160 30400 129320 30560
rect 129160 30560 129320 30720
rect 129160 30720 129320 30880
rect 129160 47680 129320 47840
rect 129160 47840 129320 48000
rect 129160 48000 129320 48160
rect 129160 48160 129320 48320
rect 129160 48320 129320 48480
rect 129160 48480 129320 48640
rect 129160 48640 129320 48800
rect 129160 48800 129320 48960
rect 129160 48960 129320 49120
rect 129160 49120 129320 49280
rect 129160 49280 129320 49440
rect 129160 49440 129320 49600
rect 129160 49600 129320 49760
rect 129160 49760 129320 49920
rect 129160 49920 129320 50080
rect 129160 50080 129320 50240
rect 129160 50240 129320 50400
rect 129160 50400 129320 50560
rect 129160 50560 129320 50720
rect 129160 50720 129320 50880
rect 129160 50880 129320 51040
rect 129160 51040 129320 51200
rect 129160 51200 129320 51360
rect 129160 51360 129320 51520
rect 129160 51520 129320 51680
rect 129160 51680 129320 51840
rect 129160 51840 129320 52000
rect 129320 27040 129480 27200
rect 129320 27200 129480 27360
rect 129320 27360 129480 27520
rect 129320 27520 129480 27680
rect 129320 27680 129480 27840
rect 129320 27840 129480 28000
rect 129320 28000 129480 28160
rect 129320 28160 129480 28320
rect 129320 28320 129480 28480
rect 129320 28480 129480 28640
rect 129320 28640 129480 28800
rect 129320 28800 129480 28960
rect 129320 28960 129480 29120
rect 129320 29120 129480 29280
rect 129320 29280 129480 29440
rect 129320 29440 129480 29600
rect 129320 29600 129480 29760
rect 129320 29760 129480 29920
rect 129320 29920 129480 30080
rect 129320 30080 129480 30240
rect 129320 30240 129480 30400
rect 129320 30400 129480 30560
rect 129320 30560 129480 30720
rect 129320 30720 129480 30880
rect 129320 48000 129480 48160
rect 129320 48160 129480 48320
rect 129320 48320 129480 48480
rect 129320 48480 129480 48640
rect 129320 48640 129480 48800
rect 129320 48800 129480 48960
rect 129320 48960 129480 49120
rect 129320 49120 129480 49280
rect 129320 49280 129480 49440
rect 129320 49440 129480 49600
rect 129320 49600 129480 49760
rect 129320 49760 129480 49920
rect 129320 49920 129480 50080
rect 129320 50080 129480 50240
rect 129320 50240 129480 50400
rect 129320 50400 129480 50560
rect 129320 50560 129480 50720
rect 129320 50720 129480 50880
rect 129320 50880 129480 51040
rect 129320 51040 129480 51200
rect 129320 51200 129480 51360
rect 129320 51360 129480 51520
rect 129320 51520 129480 51680
rect 129320 51680 129480 51840
rect 129320 51840 129480 52000
rect 129320 52000 129480 52160
rect 129480 27040 129640 27200
rect 129480 27200 129640 27360
rect 129480 27360 129640 27520
rect 129480 27520 129640 27680
rect 129480 27680 129640 27840
rect 129480 27840 129640 28000
rect 129480 28000 129640 28160
rect 129480 28160 129640 28320
rect 129480 28320 129640 28480
rect 129480 28480 129640 28640
rect 129480 28640 129640 28800
rect 129480 28800 129640 28960
rect 129480 28960 129640 29120
rect 129480 29120 129640 29280
rect 129480 29280 129640 29440
rect 129480 29440 129640 29600
rect 129480 29600 129640 29760
rect 129480 29760 129640 29920
rect 129480 29920 129640 30080
rect 129480 30080 129640 30240
rect 129480 30240 129640 30400
rect 129480 30400 129640 30560
rect 129480 30560 129640 30720
rect 129480 48000 129640 48160
rect 129480 48160 129640 48320
rect 129480 48320 129640 48480
rect 129480 48480 129640 48640
rect 129480 48640 129640 48800
rect 129480 48800 129640 48960
rect 129480 48960 129640 49120
rect 129480 49120 129640 49280
rect 129480 49280 129640 49440
rect 129480 49440 129640 49600
rect 129480 49600 129640 49760
rect 129480 49760 129640 49920
rect 129480 49920 129640 50080
rect 129480 50080 129640 50240
rect 129480 50240 129640 50400
rect 129480 50400 129640 50560
rect 129480 50560 129640 50720
rect 129480 50720 129640 50880
rect 129480 50880 129640 51040
rect 129480 51040 129640 51200
rect 129480 51200 129640 51360
rect 129480 51360 129640 51520
rect 129480 51520 129640 51680
rect 129480 51680 129640 51840
rect 129480 51840 129640 52000
rect 129480 52000 129640 52160
rect 129640 27040 129800 27200
rect 129640 27200 129800 27360
rect 129640 27360 129800 27520
rect 129640 27520 129800 27680
rect 129640 27680 129800 27840
rect 129640 27840 129800 28000
rect 129640 28000 129800 28160
rect 129640 28160 129800 28320
rect 129640 28320 129800 28480
rect 129640 28480 129800 28640
rect 129640 28640 129800 28800
rect 129640 28800 129800 28960
rect 129640 28960 129800 29120
rect 129640 29120 129800 29280
rect 129640 29280 129800 29440
rect 129640 29440 129800 29600
rect 129640 29600 129800 29760
rect 129640 29760 129800 29920
rect 129640 29920 129800 30080
rect 129640 30080 129800 30240
rect 129640 30240 129800 30400
rect 129640 30400 129800 30560
rect 129640 30560 129800 30720
rect 129640 48160 129800 48320
rect 129640 48320 129800 48480
rect 129640 48480 129800 48640
rect 129640 48640 129800 48800
rect 129640 48800 129800 48960
rect 129640 48960 129800 49120
rect 129640 49120 129800 49280
rect 129640 49280 129800 49440
rect 129640 49440 129800 49600
rect 129640 49600 129800 49760
rect 129640 49760 129800 49920
rect 129640 49920 129800 50080
rect 129640 50080 129800 50240
rect 129640 50240 129800 50400
rect 129640 50400 129800 50560
rect 129640 50560 129800 50720
rect 129640 50720 129800 50880
rect 129640 50880 129800 51040
rect 129640 51040 129800 51200
rect 129640 51200 129800 51360
rect 129640 51360 129800 51520
rect 129640 51520 129800 51680
rect 129640 51680 129800 51840
rect 129640 51840 129800 52000
rect 129640 52000 129800 52160
rect 129640 52160 129800 52320
rect 129800 26880 129960 27040
rect 129800 27040 129960 27200
rect 129800 27200 129960 27360
rect 129800 27360 129960 27520
rect 129800 27520 129960 27680
rect 129800 27680 129960 27840
rect 129800 27840 129960 28000
rect 129800 28000 129960 28160
rect 129800 28160 129960 28320
rect 129800 28320 129960 28480
rect 129800 28480 129960 28640
rect 129800 28640 129960 28800
rect 129800 28800 129960 28960
rect 129800 28960 129960 29120
rect 129800 29120 129960 29280
rect 129800 29280 129960 29440
rect 129800 29440 129960 29600
rect 129800 29600 129960 29760
rect 129800 29760 129960 29920
rect 129800 29920 129960 30080
rect 129800 30080 129960 30240
rect 129800 30240 129960 30400
rect 129800 30400 129960 30560
rect 129800 48320 129960 48480
rect 129800 48480 129960 48640
rect 129800 48640 129960 48800
rect 129800 48800 129960 48960
rect 129800 48960 129960 49120
rect 129800 49120 129960 49280
rect 129800 49280 129960 49440
rect 129800 49440 129960 49600
rect 129800 49600 129960 49760
rect 129800 49760 129960 49920
rect 129800 49920 129960 50080
rect 129800 50080 129960 50240
rect 129800 50240 129960 50400
rect 129800 50400 129960 50560
rect 129800 50560 129960 50720
rect 129800 50720 129960 50880
rect 129800 50880 129960 51040
rect 129800 51040 129960 51200
rect 129800 51200 129960 51360
rect 129800 51360 129960 51520
rect 129800 51520 129960 51680
rect 129800 51680 129960 51840
rect 129800 51840 129960 52000
rect 129800 52000 129960 52160
rect 129800 52160 129960 52320
rect 129960 26880 130120 27040
rect 129960 27040 130120 27200
rect 129960 27200 130120 27360
rect 129960 27360 130120 27520
rect 129960 27520 130120 27680
rect 129960 27680 130120 27840
rect 129960 27840 130120 28000
rect 129960 28000 130120 28160
rect 129960 28160 130120 28320
rect 129960 28320 130120 28480
rect 129960 28480 130120 28640
rect 129960 28640 130120 28800
rect 129960 28800 130120 28960
rect 129960 28960 130120 29120
rect 129960 29120 130120 29280
rect 129960 29280 130120 29440
rect 129960 29440 130120 29600
rect 129960 29600 130120 29760
rect 129960 29760 130120 29920
rect 129960 29920 130120 30080
rect 129960 30080 130120 30240
rect 129960 30240 130120 30400
rect 129960 30400 130120 30560
rect 129960 48480 130120 48640
rect 129960 48640 130120 48800
rect 129960 48800 130120 48960
rect 129960 48960 130120 49120
rect 129960 49120 130120 49280
rect 129960 49280 130120 49440
rect 129960 49440 130120 49600
rect 129960 49600 130120 49760
rect 129960 49760 130120 49920
rect 129960 49920 130120 50080
rect 129960 50080 130120 50240
rect 129960 50240 130120 50400
rect 129960 50400 130120 50560
rect 129960 50560 130120 50720
rect 129960 50720 130120 50880
rect 129960 50880 130120 51040
rect 129960 51040 130120 51200
rect 129960 51200 130120 51360
rect 129960 51360 130120 51520
rect 129960 51520 130120 51680
rect 129960 51680 130120 51840
rect 129960 51840 130120 52000
rect 129960 52000 130120 52160
rect 129960 52160 130120 52320
rect 129960 52320 130120 52480
rect 130120 26880 130280 27040
rect 130120 27040 130280 27200
rect 130120 27200 130280 27360
rect 130120 27360 130280 27520
rect 130120 27520 130280 27680
rect 130120 27680 130280 27840
rect 130120 27840 130280 28000
rect 130120 28000 130280 28160
rect 130120 28160 130280 28320
rect 130120 28320 130280 28480
rect 130120 28480 130280 28640
rect 130120 28640 130280 28800
rect 130120 28800 130280 28960
rect 130120 28960 130280 29120
rect 130120 29120 130280 29280
rect 130120 29280 130280 29440
rect 130120 29440 130280 29600
rect 130120 29600 130280 29760
rect 130120 29760 130280 29920
rect 130120 29920 130280 30080
rect 130120 30080 130280 30240
rect 130120 30240 130280 30400
rect 130120 48640 130280 48800
rect 130120 48800 130280 48960
rect 130120 48960 130280 49120
rect 130120 49120 130280 49280
rect 130120 49280 130280 49440
rect 130120 49440 130280 49600
rect 130120 49600 130280 49760
rect 130120 49760 130280 49920
rect 130120 49920 130280 50080
rect 130120 50080 130280 50240
rect 130120 50240 130280 50400
rect 130120 50400 130280 50560
rect 130120 50560 130280 50720
rect 130120 50720 130280 50880
rect 130120 50880 130280 51040
rect 130120 51040 130280 51200
rect 130120 51200 130280 51360
rect 130120 51360 130280 51520
rect 130120 51520 130280 51680
rect 130120 51680 130280 51840
rect 130120 51840 130280 52000
rect 130120 52000 130280 52160
rect 130120 52160 130280 52320
rect 130120 52320 130280 52480
rect 130280 26720 130440 26880
rect 130280 26880 130440 27040
rect 130280 27040 130440 27200
rect 130280 27200 130440 27360
rect 130280 27360 130440 27520
rect 130280 27520 130440 27680
rect 130280 27680 130440 27840
rect 130280 27840 130440 28000
rect 130280 28000 130440 28160
rect 130280 28160 130440 28320
rect 130280 28320 130440 28480
rect 130280 28480 130440 28640
rect 130280 28640 130440 28800
rect 130280 28800 130440 28960
rect 130280 28960 130440 29120
rect 130280 29120 130440 29280
rect 130280 29280 130440 29440
rect 130280 29440 130440 29600
rect 130280 29600 130440 29760
rect 130280 29760 130440 29920
rect 130280 29920 130440 30080
rect 130280 30080 130440 30240
rect 130280 30240 130440 30400
rect 130280 48640 130440 48800
rect 130280 48800 130440 48960
rect 130280 48960 130440 49120
rect 130280 49120 130440 49280
rect 130280 49280 130440 49440
rect 130280 49440 130440 49600
rect 130280 49600 130440 49760
rect 130280 49760 130440 49920
rect 130280 49920 130440 50080
rect 130280 50080 130440 50240
rect 130280 50240 130440 50400
rect 130280 50400 130440 50560
rect 130280 50560 130440 50720
rect 130280 50720 130440 50880
rect 130280 50880 130440 51040
rect 130280 51040 130440 51200
rect 130280 51200 130440 51360
rect 130280 51360 130440 51520
rect 130280 51520 130440 51680
rect 130280 51680 130440 51840
rect 130280 51840 130440 52000
rect 130280 52000 130440 52160
rect 130280 52160 130440 52320
rect 130280 52320 130440 52480
rect 130440 26720 130600 26880
rect 130440 26880 130600 27040
rect 130440 27040 130600 27200
rect 130440 27200 130600 27360
rect 130440 27360 130600 27520
rect 130440 27520 130600 27680
rect 130440 27680 130600 27840
rect 130440 27840 130600 28000
rect 130440 28000 130600 28160
rect 130440 28160 130600 28320
rect 130440 28320 130600 28480
rect 130440 28480 130600 28640
rect 130440 28640 130600 28800
rect 130440 28800 130600 28960
rect 130440 28960 130600 29120
rect 130440 29120 130600 29280
rect 130440 29280 130600 29440
rect 130440 29440 130600 29600
rect 130440 29600 130600 29760
rect 130440 29760 130600 29920
rect 130440 29920 130600 30080
rect 130440 30080 130600 30240
rect 130440 30240 130600 30400
rect 130440 48800 130600 48960
rect 130440 48960 130600 49120
rect 130440 49120 130600 49280
rect 130440 49280 130600 49440
rect 130440 49440 130600 49600
rect 130440 49600 130600 49760
rect 130440 49760 130600 49920
rect 130440 49920 130600 50080
rect 130440 50080 130600 50240
rect 130440 50240 130600 50400
rect 130440 50400 130600 50560
rect 130440 50560 130600 50720
rect 130440 50720 130600 50880
rect 130440 50880 130600 51040
rect 130440 51040 130600 51200
rect 130440 51200 130600 51360
rect 130440 51360 130600 51520
rect 130440 51520 130600 51680
rect 130440 51680 130600 51840
rect 130440 51840 130600 52000
rect 130440 52000 130600 52160
rect 130440 52160 130600 52320
rect 130440 52320 130600 52480
rect 130440 52480 130600 52640
rect 130600 26720 130760 26880
rect 130600 26880 130760 27040
rect 130600 27040 130760 27200
rect 130600 27200 130760 27360
rect 130600 27360 130760 27520
rect 130600 27520 130760 27680
rect 130600 27680 130760 27840
rect 130600 27840 130760 28000
rect 130600 28000 130760 28160
rect 130600 28160 130760 28320
rect 130600 28320 130760 28480
rect 130600 28480 130760 28640
rect 130600 28640 130760 28800
rect 130600 28800 130760 28960
rect 130600 28960 130760 29120
rect 130600 29120 130760 29280
rect 130600 29280 130760 29440
rect 130600 29440 130760 29600
rect 130600 29600 130760 29760
rect 130600 29760 130760 29920
rect 130600 29920 130760 30080
rect 130600 30080 130760 30240
rect 130600 48800 130760 48960
rect 130600 48960 130760 49120
rect 130600 49120 130760 49280
rect 130600 49280 130760 49440
rect 130600 49440 130760 49600
rect 130600 49600 130760 49760
rect 130600 49760 130760 49920
rect 130600 49920 130760 50080
rect 130600 50080 130760 50240
rect 130600 50240 130760 50400
rect 130600 50400 130760 50560
rect 130600 50560 130760 50720
rect 130600 50720 130760 50880
rect 130600 50880 130760 51040
rect 130600 51040 130760 51200
rect 130600 51200 130760 51360
rect 130600 51360 130760 51520
rect 130600 51520 130760 51680
rect 130600 51680 130760 51840
rect 130600 51840 130760 52000
rect 130600 52000 130760 52160
rect 130600 52160 130760 52320
rect 130600 52320 130760 52480
rect 130600 52480 130760 52640
rect 130760 26720 130920 26880
rect 130760 26880 130920 27040
rect 130760 27040 130920 27200
rect 130760 27200 130920 27360
rect 130760 27360 130920 27520
rect 130760 27520 130920 27680
rect 130760 27680 130920 27840
rect 130760 27840 130920 28000
rect 130760 28000 130920 28160
rect 130760 28160 130920 28320
rect 130760 28320 130920 28480
rect 130760 28480 130920 28640
rect 130760 28640 130920 28800
rect 130760 28800 130920 28960
rect 130760 28960 130920 29120
rect 130760 29120 130920 29280
rect 130760 29280 130920 29440
rect 130760 29440 130920 29600
rect 130760 29600 130920 29760
rect 130760 29760 130920 29920
rect 130760 29920 130920 30080
rect 130760 30080 130920 30240
rect 130760 48960 130920 49120
rect 130760 49120 130920 49280
rect 130760 49280 130920 49440
rect 130760 49440 130920 49600
rect 130760 49600 130920 49760
rect 130760 49760 130920 49920
rect 130760 49920 130920 50080
rect 130760 50080 130920 50240
rect 130760 50240 130920 50400
rect 130760 50400 130920 50560
rect 130760 50560 130920 50720
rect 130760 50720 130920 50880
rect 130760 50880 130920 51040
rect 130760 51040 130920 51200
rect 130760 51200 130920 51360
rect 130760 51360 130920 51520
rect 130760 51520 130920 51680
rect 130760 51680 130920 51840
rect 130760 51840 130920 52000
rect 130760 52000 130920 52160
rect 130760 52160 130920 52320
rect 130760 52320 130920 52480
rect 130760 52480 130920 52640
rect 130920 26720 131080 26880
rect 130920 26880 131080 27040
rect 130920 27040 131080 27200
rect 130920 27200 131080 27360
rect 130920 27360 131080 27520
rect 130920 27520 131080 27680
rect 130920 27680 131080 27840
rect 130920 27840 131080 28000
rect 130920 28000 131080 28160
rect 130920 28160 131080 28320
rect 130920 28320 131080 28480
rect 130920 28480 131080 28640
rect 130920 28640 131080 28800
rect 130920 28800 131080 28960
rect 130920 28960 131080 29120
rect 130920 29120 131080 29280
rect 130920 29280 131080 29440
rect 130920 29440 131080 29600
rect 130920 29600 131080 29760
rect 130920 29760 131080 29920
rect 130920 29920 131080 30080
rect 130920 30080 131080 30240
rect 130920 48960 131080 49120
rect 130920 49120 131080 49280
rect 130920 49280 131080 49440
rect 130920 49440 131080 49600
rect 130920 49600 131080 49760
rect 130920 49760 131080 49920
rect 130920 49920 131080 50080
rect 130920 50080 131080 50240
rect 130920 50240 131080 50400
rect 130920 50400 131080 50560
rect 130920 50560 131080 50720
rect 130920 50720 131080 50880
rect 130920 50880 131080 51040
rect 130920 51040 131080 51200
rect 130920 51200 131080 51360
rect 130920 51360 131080 51520
rect 130920 51520 131080 51680
rect 130920 51680 131080 51840
rect 130920 51840 131080 52000
rect 130920 52000 131080 52160
rect 130920 52160 131080 52320
rect 130920 52320 131080 52480
rect 130920 52480 131080 52640
rect 130920 52640 131080 52800
rect 131080 26720 131240 26880
rect 131080 26880 131240 27040
rect 131080 27040 131240 27200
rect 131080 27200 131240 27360
rect 131080 27360 131240 27520
rect 131080 27520 131240 27680
rect 131080 27680 131240 27840
rect 131080 27840 131240 28000
rect 131080 28000 131240 28160
rect 131080 28160 131240 28320
rect 131080 28320 131240 28480
rect 131080 28480 131240 28640
rect 131080 28640 131240 28800
rect 131080 28800 131240 28960
rect 131080 28960 131240 29120
rect 131080 29120 131240 29280
rect 131080 29280 131240 29440
rect 131080 29440 131240 29600
rect 131080 29600 131240 29760
rect 131080 29760 131240 29920
rect 131080 29920 131240 30080
rect 131080 30080 131240 30240
rect 131080 49120 131240 49280
rect 131080 49280 131240 49440
rect 131080 49440 131240 49600
rect 131080 49600 131240 49760
rect 131080 49760 131240 49920
rect 131080 49920 131240 50080
rect 131080 50080 131240 50240
rect 131080 50240 131240 50400
rect 131080 50400 131240 50560
rect 131080 50560 131240 50720
rect 131080 50720 131240 50880
rect 131080 50880 131240 51040
rect 131080 51040 131240 51200
rect 131080 51200 131240 51360
rect 131080 51360 131240 51520
rect 131080 51520 131240 51680
rect 131080 51680 131240 51840
rect 131080 51840 131240 52000
rect 131080 52000 131240 52160
rect 131080 52160 131240 52320
rect 131080 52320 131240 52480
rect 131080 52480 131240 52640
rect 131080 52640 131240 52800
rect 131240 26560 131400 26720
rect 131240 26720 131400 26880
rect 131240 26880 131400 27040
rect 131240 27040 131400 27200
rect 131240 27200 131400 27360
rect 131240 27360 131400 27520
rect 131240 27520 131400 27680
rect 131240 27680 131400 27840
rect 131240 27840 131400 28000
rect 131240 28000 131400 28160
rect 131240 28160 131400 28320
rect 131240 28320 131400 28480
rect 131240 28480 131400 28640
rect 131240 28640 131400 28800
rect 131240 28800 131400 28960
rect 131240 28960 131400 29120
rect 131240 29120 131400 29280
rect 131240 29280 131400 29440
rect 131240 29440 131400 29600
rect 131240 29600 131400 29760
rect 131240 29760 131400 29920
rect 131240 29920 131400 30080
rect 131240 49120 131400 49280
rect 131240 49280 131400 49440
rect 131240 49440 131400 49600
rect 131240 49600 131400 49760
rect 131240 49760 131400 49920
rect 131240 49920 131400 50080
rect 131240 50080 131400 50240
rect 131240 50240 131400 50400
rect 131240 50400 131400 50560
rect 131240 50560 131400 50720
rect 131240 50720 131400 50880
rect 131240 50880 131400 51040
rect 131240 51040 131400 51200
rect 131240 51200 131400 51360
rect 131240 51360 131400 51520
rect 131240 51520 131400 51680
rect 131240 51680 131400 51840
rect 131240 51840 131400 52000
rect 131240 52000 131400 52160
rect 131240 52160 131400 52320
rect 131240 52320 131400 52480
rect 131240 52480 131400 52640
rect 131240 52640 131400 52800
rect 131400 26560 131560 26720
rect 131400 26720 131560 26880
rect 131400 26880 131560 27040
rect 131400 27040 131560 27200
rect 131400 27200 131560 27360
rect 131400 27360 131560 27520
rect 131400 27520 131560 27680
rect 131400 27680 131560 27840
rect 131400 27840 131560 28000
rect 131400 28000 131560 28160
rect 131400 28160 131560 28320
rect 131400 28320 131560 28480
rect 131400 28480 131560 28640
rect 131400 28640 131560 28800
rect 131400 28800 131560 28960
rect 131400 28960 131560 29120
rect 131400 29120 131560 29280
rect 131400 29280 131560 29440
rect 131400 29440 131560 29600
rect 131400 29600 131560 29760
rect 131400 29760 131560 29920
rect 131400 29920 131560 30080
rect 131400 49280 131560 49440
rect 131400 49440 131560 49600
rect 131400 49600 131560 49760
rect 131400 49760 131560 49920
rect 131400 49920 131560 50080
rect 131400 50080 131560 50240
rect 131400 50240 131560 50400
rect 131400 50400 131560 50560
rect 131400 50560 131560 50720
rect 131400 50720 131560 50880
rect 131400 50880 131560 51040
rect 131400 51040 131560 51200
rect 131400 51200 131560 51360
rect 131400 51360 131560 51520
rect 131400 51520 131560 51680
rect 131400 51680 131560 51840
rect 131400 51840 131560 52000
rect 131400 52000 131560 52160
rect 131400 52160 131560 52320
rect 131400 52320 131560 52480
rect 131400 52480 131560 52640
rect 131400 52640 131560 52800
rect 131400 52800 131560 52960
rect 131560 26560 131720 26720
rect 131560 26720 131720 26880
rect 131560 26880 131720 27040
rect 131560 27040 131720 27200
rect 131560 27200 131720 27360
rect 131560 27360 131720 27520
rect 131560 27520 131720 27680
rect 131560 27680 131720 27840
rect 131560 27840 131720 28000
rect 131560 28000 131720 28160
rect 131560 28160 131720 28320
rect 131560 28320 131720 28480
rect 131560 28480 131720 28640
rect 131560 28640 131720 28800
rect 131560 28800 131720 28960
rect 131560 28960 131720 29120
rect 131560 29120 131720 29280
rect 131560 29280 131720 29440
rect 131560 29440 131720 29600
rect 131560 29600 131720 29760
rect 131560 29760 131720 29920
rect 131560 29920 131720 30080
rect 131560 49280 131720 49440
rect 131560 49440 131720 49600
rect 131560 49600 131720 49760
rect 131560 49760 131720 49920
rect 131560 49920 131720 50080
rect 131560 50080 131720 50240
rect 131560 50240 131720 50400
rect 131560 50400 131720 50560
rect 131560 50560 131720 50720
rect 131560 50720 131720 50880
rect 131560 50880 131720 51040
rect 131560 51040 131720 51200
rect 131560 51200 131720 51360
rect 131560 51360 131720 51520
rect 131560 51520 131720 51680
rect 131560 51680 131720 51840
rect 131560 51840 131720 52000
rect 131560 52000 131720 52160
rect 131560 52160 131720 52320
rect 131560 52320 131720 52480
rect 131560 52480 131720 52640
rect 131560 52640 131720 52800
rect 131560 52800 131720 52960
rect 131720 26560 131880 26720
rect 131720 26720 131880 26880
rect 131720 26880 131880 27040
rect 131720 27040 131880 27200
rect 131720 27200 131880 27360
rect 131720 27360 131880 27520
rect 131720 27520 131880 27680
rect 131720 27680 131880 27840
rect 131720 27840 131880 28000
rect 131720 28000 131880 28160
rect 131720 28160 131880 28320
rect 131720 28320 131880 28480
rect 131720 28480 131880 28640
rect 131720 28640 131880 28800
rect 131720 28800 131880 28960
rect 131720 28960 131880 29120
rect 131720 29120 131880 29280
rect 131720 29280 131880 29440
rect 131720 29440 131880 29600
rect 131720 29600 131880 29760
rect 131720 29760 131880 29920
rect 131720 29920 131880 30080
rect 131720 49440 131880 49600
rect 131720 49600 131880 49760
rect 131720 49760 131880 49920
rect 131720 49920 131880 50080
rect 131720 50080 131880 50240
rect 131720 50240 131880 50400
rect 131720 50400 131880 50560
rect 131720 50560 131880 50720
rect 131720 50720 131880 50880
rect 131720 50880 131880 51040
rect 131720 51040 131880 51200
rect 131720 51200 131880 51360
rect 131720 51360 131880 51520
rect 131720 51520 131880 51680
rect 131720 51680 131880 51840
rect 131720 51840 131880 52000
rect 131720 52000 131880 52160
rect 131720 52160 131880 52320
rect 131720 52320 131880 52480
rect 131720 52480 131880 52640
rect 131720 52640 131880 52800
rect 131720 52800 131880 52960
rect 131880 26560 132040 26720
rect 131880 26720 132040 26880
rect 131880 26880 132040 27040
rect 131880 27040 132040 27200
rect 131880 27200 132040 27360
rect 131880 27360 132040 27520
rect 131880 27520 132040 27680
rect 131880 27680 132040 27840
rect 131880 27840 132040 28000
rect 131880 28000 132040 28160
rect 131880 28160 132040 28320
rect 131880 28320 132040 28480
rect 131880 28480 132040 28640
rect 131880 28640 132040 28800
rect 131880 28800 132040 28960
rect 131880 28960 132040 29120
rect 131880 29120 132040 29280
rect 131880 29280 132040 29440
rect 131880 29440 132040 29600
rect 131880 29600 132040 29760
rect 131880 29760 132040 29920
rect 131880 29920 132040 30080
rect 131880 49440 132040 49600
rect 131880 49600 132040 49760
rect 131880 49760 132040 49920
rect 131880 49920 132040 50080
rect 131880 50080 132040 50240
rect 131880 50240 132040 50400
rect 131880 50400 132040 50560
rect 131880 50560 132040 50720
rect 131880 50720 132040 50880
rect 131880 50880 132040 51040
rect 131880 51040 132040 51200
rect 131880 51200 132040 51360
rect 131880 51360 132040 51520
rect 131880 51520 132040 51680
rect 131880 51680 132040 51840
rect 131880 51840 132040 52000
rect 131880 52000 132040 52160
rect 131880 52160 132040 52320
rect 131880 52320 132040 52480
rect 131880 52480 132040 52640
rect 131880 52640 132040 52800
rect 131880 52800 132040 52960
rect 132040 26560 132200 26720
rect 132040 26720 132200 26880
rect 132040 26880 132200 27040
rect 132040 27040 132200 27200
rect 132040 27200 132200 27360
rect 132040 27360 132200 27520
rect 132040 27520 132200 27680
rect 132040 27680 132200 27840
rect 132040 27840 132200 28000
rect 132040 28000 132200 28160
rect 132040 28160 132200 28320
rect 132040 28320 132200 28480
rect 132040 28480 132200 28640
rect 132040 28640 132200 28800
rect 132040 28800 132200 28960
rect 132040 28960 132200 29120
rect 132040 29120 132200 29280
rect 132040 29280 132200 29440
rect 132040 29440 132200 29600
rect 132040 29600 132200 29760
rect 132040 29760 132200 29920
rect 132040 29920 132200 30080
rect 132040 49440 132200 49600
rect 132040 49600 132200 49760
rect 132040 49760 132200 49920
rect 132040 49920 132200 50080
rect 132040 50080 132200 50240
rect 132040 50240 132200 50400
rect 132040 50400 132200 50560
rect 132040 50560 132200 50720
rect 132040 50720 132200 50880
rect 132040 50880 132200 51040
rect 132040 51040 132200 51200
rect 132040 51200 132200 51360
rect 132040 51360 132200 51520
rect 132040 51520 132200 51680
rect 132040 51680 132200 51840
rect 132040 51840 132200 52000
rect 132040 52000 132200 52160
rect 132040 52160 132200 52320
rect 132040 52320 132200 52480
rect 132040 52480 132200 52640
rect 132040 52640 132200 52800
rect 132040 52800 132200 52960
rect 132040 52960 132200 53120
rect 132200 26560 132360 26720
rect 132200 26720 132360 26880
rect 132200 26880 132360 27040
rect 132200 27040 132360 27200
rect 132200 27200 132360 27360
rect 132200 27360 132360 27520
rect 132200 27520 132360 27680
rect 132200 27680 132360 27840
rect 132200 27840 132360 28000
rect 132200 28000 132360 28160
rect 132200 28160 132360 28320
rect 132200 28320 132360 28480
rect 132200 28480 132360 28640
rect 132200 28640 132360 28800
rect 132200 28800 132360 28960
rect 132200 28960 132360 29120
rect 132200 29120 132360 29280
rect 132200 29280 132360 29440
rect 132200 29440 132360 29600
rect 132200 29600 132360 29760
rect 132200 29760 132360 29920
rect 132200 29920 132360 30080
rect 132200 49600 132360 49760
rect 132200 49760 132360 49920
rect 132200 49920 132360 50080
rect 132200 50080 132360 50240
rect 132200 50240 132360 50400
rect 132200 50400 132360 50560
rect 132200 50560 132360 50720
rect 132200 50720 132360 50880
rect 132200 50880 132360 51040
rect 132200 51040 132360 51200
rect 132200 51200 132360 51360
rect 132200 51360 132360 51520
rect 132200 51520 132360 51680
rect 132200 51680 132360 51840
rect 132200 51840 132360 52000
rect 132200 52000 132360 52160
rect 132200 52160 132360 52320
rect 132200 52320 132360 52480
rect 132200 52480 132360 52640
rect 132200 52640 132360 52800
rect 132200 52800 132360 52960
rect 132200 52960 132360 53120
rect 132360 26560 132520 26720
rect 132360 26720 132520 26880
rect 132360 26880 132520 27040
rect 132360 27040 132520 27200
rect 132360 27200 132520 27360
rect 132360 27360 132520 27520
rect 132360 27520 132520 27680
rect 132360 27680 132520 27840
rect 132360 27840 132520 28000
rect 132360 28000 132520 28160
rect 132360 28160 132520 28320
rect 132360 28320 132520 28480
rect 132360 28480 132520 28640
rect 132360 28640 132520 28800
rect 132360 28800 132520 28960
rect 132360 28960 132520 29120
rect 132360 29120 132520 29280
rect 132360 29280 132520 29440
rect 132360 29440 132520 29600
rect 132360 29600 132520 29760
rect 132360 29760 132520 29920
rect 132360 29920 132520 30080
rect 132360 49600 132520 49760
rect 132360 49760 132520 49920
rect 132360 49920 132520 50080
rect 132360 50080 132520 50240
rect 132360 50240 132520 50400
rect 132360 50400 132520 50560
rect 132360 50560 132520 50720
rect 132360 50720 132520 50880
rect 132360 50880 132520 51040
rect 132360 51040 132520 51200
rect 132360 51200 132520 51360
rect 132360 51360 132520 51520
rect 132360 51520 132520 51680
rect 132360 51680 132520 51840
rect 132360 51840 132520 52000
rect 132360 52000 132520 52160
rect 132360 52160 132520 52320
rect 132360 52320 132520 52480
rect 132360 52480 132520 52640
rect 132360 52640 132520 52800
rect 132360 52800 132520 52960
rect 132360 52960 132520 53120
rect 132520 26560 132680 26720
rect 132520 26720 132680 26880
rect 132520 26880 132680 27040
rect 132520 27040 132680 27200
rect 132520 27200 132680 27360
rect 132520 27360 132680 27520
rect 132520 27520 132680 27680
rect 132520 27680 132680 27840
rect 132520 27840 132680 28000
rect 132520 28000 132680 28160
rect 132520 28160 132680 28320
rect 132520 28320 132680 28480
rect 132520 28480 132680 28640
rect 132520 28640 132680 28800
rect 132520 28800 132680 28960
rect 132520 28960 132680 29120
rect 132520 29120 132680 29280
rect 132520 29280 132680 29440
rect 132520 29440 132680 29600
rect 132520 29600 132680 29760
rect 132520 29760 132680 29920
rect 132520 29920 132680 30080
rect 132520 49600 132680 49760
rect 132520 49760 132680 49920
rect 132520 49920 132680 50080
rect 132520 50080 132680 50240
rect 132520 50240 132680 50400
rect 132520 50400 132680 50560
rect 132520 50560 132680 50720
rect 132520 50720 132680 50880
rect 132520 50880 132680 51040
rect 132520 51040 132680 51200
rect 132520 51200 132680 51360
rect 132520 51360 132680 51520
rect 132520 51520 132680 51680
rect 132520 51680 132680 51840
rect 132520 51840 132680 52000
rect 132520 52000 132680 52160
rect 132520 52160 132680 52320
rect 132520 52320 132680 52480
rect 132520 52480 132680 52640
rect 132520 52640 132680 52800
rect 132520 52800 132680 52960
rect 132520 52960 132680 53120
rect 132680 26560 132840 26720
rect 132680 26720 132840 26880
rect 132680 26880 132840 27040
rect 132680 27040 132840 27200
rect 132680 27200 132840 27360
rect 132680 27360 132840 27520
rect 132680 27520 132840 27680
rect 132680 27680 132840 27840
rect 132680 27840 132840 28000
rect 132680 28000 132840 28160
rect 132680 28160 132840 28320
rect 132680 28320 132840 28480
rect 132680 28480 132840 28640
rect 132680 28640 132840 28800
rect 132680 28800 132840 28960
rect 132680 28960 132840 29120
rect 132680 29120 132840 29280
rect 132680 29280 132840 29440
rect 132680 29440 132840 29600
rect 132680 29600 132840 29760
rect 132680 29760 132840 29920
rect 132680 29920 132840 30080
rect 132680 49600 132840 49760
rect 132680 49760 132840 49920
rect 132680 49920 132840 50080
rect 132680 50080 132840 50240
rect 132680 50240 132840 50400
rect 132680 50400 132840 50560
rect 132680 50560 132840 50720
rect 132680 50720 132840 50880
rect 132680 50880 132840 51040
rect 132680 51040 132840 51200
rect 132680 51200 132840 51360
rect 132680 51360 132840 51520
rect 132680 51520 132840 51680
rect 132680 51680 132840 51840
rect 132680 51840 132840 52000
rect 132680 52000 132840 52160
rect 132680 52160 132840 52320
rect 132680 52320 132840 52480
rect 132680 52480 132840 52640
rect 132680 52640 132840 52800
rect 132680 52800 132840 52960
rect 132680 52960 132840 53120
rect 132840 26560 133000 26720
rect 132840 26720 133000 26880
rect 132840 26880 133000 27040
rect 132840 27040 133000 27200
rect 132840 27200 133000 27360
rect 132840 27360 133000 27520
rect 132840 27520 133000 27680
rect 132840 27680 133000 27840
rect 132840 27840 133000 28000
rect 132840 28000 133000 28160
rect 132840 28160 133000 28320
rect 132840 28320 133000 28480
rect 132840 28480 133000 28640
rect 132840 28640 133000 28800
rect 132840 28800 133000 28960
rect 132840 28960 133000 29120
rect 132840 29120 133000 29280
rect 132840 29280 133000 29440
rect 132840 29440 133000 29600
rect 132840 29600 133000 29760
rect 132840 29760 133000 29920
rect 132840 29920 133000 30080
rect 132840 49600 133000 49760
rect 132840 49760 133000 49920
rect 132840 49920 133000 50080
rect 132840 50080 133000 50240
rect 132840 50240 133000 50400
rect 132840 50400 133000 50560
rect 132840 50560 133000 50720
rect 132840 50720 133000 50880
rect 132840 50880 133000 51040
rect 132840 51040 133000 51200
rect 132840 51200 133000 51360
rect 132840 51360 133000 51520
rect 132840 51520 133000 51680
rect 132840 51680 133000 51840
rect 132840 51840 133000 52000
rect 132840 52000 133000 52160
rect 132840 52160 133000 52320
rect 132840 52320 133000 52480
rect 132840 52480 133000 52640
rect 132840 52640 133000 52800
rect 132840 52800 133000 52960
rect 132840 52960 133000 53120
rect 133000 26560 133160 26720
rect 133000 26720 133160 26880
rect 133000 26880 133160 27040
rect 133000 27040 133160 27200
rect 133000 27200 133160 27360
rect 133000 27360 133160 27520
rect 133000 27520 133160 27680
rect 133000 27680 133160 27840
rect 133000 27840 133160 28000
rect 133000 28000 133160 28160
rect 133000 28160 133160 28320
rect 133000 28320 133160 28480
rect 133000 28480 133160 28640
rect 133000 28640 133160 28800
rect 133000 28800 133160 28960
rect 133000 28960 133160 29120
rect 133000 29120 133160 29280
rect 133000 29280 133160 29440
rect 133000 29440 133160 29600
rect 133000 29600 133160 29760
rect 133000 29760 133160 29920
rect 133000 29920 133160 30080
rect 133000 49760 133160 49920
rect 133000 49920 133160 50080
rect 133000 50080 133160 50240
rect 133000 50240 133160 50400
rect 133000 50400 133160 50560
rect 133000 50560 133160 50720
rect 133000 50720 133160 50880
rect 133000 50880 133160 51040
rect 133000 51040 133160 51200
rect 133000 51200 133160 51360
rect 133000 51360 133160 51520
rect 133000 51520 133160 51680
rect 133000 51680 133160 51840
rect 133000 51840 133160 52000
rect 133000 52000 133160 52160
rect 133000 52160 133160 52320
rect 133000 52320 133160 52480
rect 133000 52480 133160 52640
rect 133000 52640 133160 52800
rect 133000 52800 133160 52960
rect 133000 52960 133160 53120
rect 133160 26560 133320 26720
rect 133160 26720 133320 26880
rect 133160 26880 133320 27040
rect 133160 27040 133320 27200
rect 133160 27200 133320 27360
rect 133160 27360 133320 27520
rect 133160 27520 133320 27680
rect 133160 27680 133320 27840
rect 133160 27840 133320 28000
rect 133160 28000 133320 28160
rect 133160 28160 133320 28320
rect 133160 28320 133320 28480
rect 133160 28480 133320 28640
rect 133160 28640 133320 28800
rect 133160 28800 133320 28960
rect 133160 28960 133320 29120
rect 133160 29120 133320 29280
rect 133160 29280 133320 29440
rect 133160 29440 133320 29600
rect 133160 29600 133320 29760
rect 133160 29760 133320 29920
rect 133160 29920 133320 30080
rect 133160 49760 133320 49920
rect 133160 49920 133320 50080
rect 133160 50080 133320 50240
rect 133160 50240 133320 50400
rect 133160 50400 133320 50560
rect 133160 50560 133320 50720
rect 133160 50720 133320 50880
rect 133160 50880 133320 51040
rect 133160 51040 133320 51200
rect 133160 51200 133320 51360
rect 133160 51360 133320 51520
rect 133160 51520 133320 51680
rect 133160 51680 133320 51840
rect 133160 51840 133320 52000
rect 133160 52000 133320 52160
rect 133160 52160 133320 52320
rect 133160 52320 133320 52480
rect 133160 52480 133320 52640
rect 133160 52640 133320 52800
rect 133160 52800 133320 52960
rect 133160 52960 133320 53120
rect 133160 53120 133320 53280
rect 133320 26560 133480 26720
rect 133320 26720 133480 26880
rect 133320 26880 133480 27040
rect 133320 27040 133480 27200
rect 133320 27200 133480 27360
rect 133320 27360 133480 27520
rect 133320 27520 133480 27680
rect 133320 27680 133480 27840
rect 133320 27840 133480 28000
rect 133320 28000 133480 28160
rect 133320 28160 133480 28320
rect 133320 28320 133480 28480
rect 133320 28480 133480 28640
rect 133320 28640 133480 28800
rect 133320 28800 133480 28960
rect 133320 28960 133480 29120
rect 133320 29120 133480 29280
rect 133320 29280 133480 29440
rect 133320 29440 133480 29600
rect 133320 29600 133480 29760
rect 133320 29760 133480 29920
rect 133320 29920 133480 30080
rect 133320 49760 133480 49920
rect 133320 49920 133480 50080
rect 133320 50080 133480 50240
rect 133320 50240 133480 50400
rect 133320 50400 133480 50560
rect 133320 50560 133480 50720
rect 133320 50720 133480 50880
rect 133320 50880 133480 51040
rect 133320 51040 133480 51200
rect 133320 51200 133480 51360
rect 133320 51360 133480 51520
rect 133320 51520 133480 51680
rect 133320 51680 133480 51840
rect 133320 51840 133480 52000
rect 133320 52000 133480 52160
rect 133320 52160 133480 52320
rect 133320 52320 133480 52480
rect 133320 52480 133480 52640
rect 133320 52640 133480 52800
rect 133320 52800 133480 52960
rect 133320 52960 133480 53120
rect 133320 53120 133480 53280
rect 133480 26560 133640 26720
rect 133480 26720 133640 26880
rect 133480 26880 133640 27040
rect 133480 27040 133640 27200
rect 133480 27200 133640 27360
rect 133480 27360 133640 27520
rect 133480 27520 133640 27680
rect 133480 27680 133640 27840
rect 133480 27840 133640 28000
rect 133480 28000 133640 28160
rect 133480 28160 133640 28320
rect 133480 28320 133640 28480
rect 133480 28480 133640 28640
rect 133480 28640 133640 28800
rect 133480 28800 133640 28960
rect 133480 28960 133640 29120
rect 133480 29120 133640 29280
rect 133480 29280 133640 29440
rect 133480 29440 133640 29600
rect 133480 29600 133640 29760
rect 133480 29760 133640 29920
rect 133480 29920 133640 30080
rect 133480 49760 133640 49920
rect 133480 49920 133640 50080
rect 133480 50080 133640 50240
rect 133480 50240 133640 50400
rect 133480 50400 133640 50560
rect 133480 50560 133640 50720
rect 133480 50720 133640 50880
rect 133480 50880 133640 51040
rect 133480 51040 133640 51200
rect 133480 51200 133640 51360
rect 133480 51360 133640 51520
rect 133480 51520 133640 51680
rect 133480 51680 133640 51840
rect 133480 51840 133640 52000
rect 133480 52000 133640 52160
rect 133480 52160 133640 52320
rect 133480 52320 133640 52480
rect 133480 52480 133640 52640
rect 133480 52640 133640 52800
rect 133480 52800 133640 52960
rect 133480 52960 133640 53120
rect 133480 53120 133640 53280
rect 133640 26560 133800 26720
rect 133640 26720 133800 26880
rect 133640 26880 133800 27040
rect 133640 27040 133800 27200
rect 133640 27200 133800 27360
rect 133640 27360 133800 27520
rect 133640 27520 133800 27680
rect 133640 27680 133800 27840
rect 133640 27840 133800 28000
rect 133640 28000 133800 28160
rect 133640 28160 133800 28320
rect 133640 28320 133800 28480
rect 133640 28480 133800 28640
rect 133640 28640 133800 28800
rect 133640 28800 133800 28960
rect 133640 28960 133800 29120
rect 133640 29120 133800 29280
rect 133640 29280 133800 29440
rect 133640 29440 133800 29600
rect 133640 29600 133800 29760
rect 133640 29760 133800 29920
rect 133640 29920 133800 30080
rect 133640 49760 133800 49920
rect 133640 49920 133800 50080
rect 133640 50080 133800 50240
rect 133640 50240 133800 50400
rect 133640 50400 133800 50560
rect 133640 50560 133800 50720
rect 133640 50720 133800 50880
rect 133640 50880 133800 51040
rect 133640 51040 133800 51200
rect 133640 51200 133800 51360
rect 133640 51360 133800 51520
rect 133640 51520 133800 51680
rect 133640 51680 133800 51840
rect 133640 51840 133800 52000
rect 133640 52000 133800 52160
rect 133640 52160 133800 52320
rect 133640 52320 133800 52480
rect 133640 52480 133800 52640
rect 133640 52640 133800 52800
rect 133640 52800 133800 52960
rect 133640 52960 133800 53120
rect 133640 53120 133800 53280
rect 133800 26560 133960 26720
rect 133800 26720 133960 26880
rect 133800 26880 133960 27040
rect 133800 27040 133960 27200
rect 133800 27200 133960 27360
rect 133800 27360 133960 27520
rect 133800 27520 133960 27680
rect 133800 27680 133960 27840
rect 133800 27840 133960 28000
rect 133800 28000 133960 28160
rect 133800 28160 133960 28320
rect 133800 28320 133960 28480
rect 133800 28480 133960 28640
rect 133800 28640 133960 28800
rect 133800 28800 133960 28960
rect 133800 28960 133960 29120
rect 133800 29120 133960 29280
rect 133800 29280 133960 29440
rect 133800 29440 133960 29600
rect 133800 29600 133960 29760
rect 133800 29760 133960 29920
rect 133800 29920 133960 30080
rect 133800 49760 133960 49920
rect 133800 49920 133960 50080
rect 133800 50080 133960 50240
rect 133800 50240 133960 50400
rect 133800 50400 133960 50560
rect 133800 50560 133960 50720
rect 133800 50720 133960 50880
rect 133800 50880 133960 51040
rect 133800 51040 133960 51200
rect 133800 51200 133960 51360
rect 133800 51360 133960 51520
rect 133800 51520 133960 51680
rect 133800 51680 133960 51840
rect 133800 51840 133960 52000
rect 133800 52000 133960 52160
rect 133800 52160 133960 52320
rect 133800 52320 133960 52480
rect 133800 52480 133960 52640
rect 133800 52640 133960 52800
rect 133800 52800 133960 52960
rect 133800 52960 133960 53120
rect 133800 53120 133960 53280
rect 133960 26560 134120 26720
rect 133960 26720 134120 26880
rect 133960 26880 134120 27040
rect 133960 27040 134120 27200
rect 133960 27200 134120 27360
rect 133960 27360 134120 27520
rect 133960 27520 134120 27680
rect 133960 27680 134120 27840
rect 133960 27840 134120 28000
rect 133960 28000 134120 28160
rect 133960 28160 134120 28320
rect 133960 28320 134120 28480
rect 133960 28480 134120 28640
rect 133960 28640 134120 28800
rect 133960 28800 134120 28960
rect 133960 28960 134120 29120
rect 133960 29120 134120 29280
rect 133960 29280 134120 29440
rect 133960 29440 134120 29600
rect 133960 29600 134120 29760
rect 133960 29760 134120 29920
rect 133960 29920 134120 30080
rect 133960 49760 134120 49920
rect 133960 49920 134120 50080
rect 133960 50080 134120 50240
rect 133960 50240 134120 50400
rect 133960 50400 134120 50560
rect 133960 50560 134120 50720
rect 133960 50720 134120 50880
rect 133960 50880 134120 51040
rect 133960 51040 134120 51200
rect 133960 51200 134120 51360
rect 133960 51360 134120 51520
rect 133960 51520 134120 51680
rect 133960 51680 134120 51840
rect 133960 51840 134120 52000
rect 133960 52000 134120 52160
rect 133960 52160 134120 52320
rect 133960 52320 134120 52480
rect 133960 52480 134120 52640
rect 133960 52640 134120 52800
rect 133960 52800 134120 52960
rect 133960 52960 134120 53120
rect 133960 53120 134120 53280
rect 134120 26720 134280 26880
rect 134120 26880 134280 27040
rect 134120 27040 134280 27200
rect 134120 27200 134280 27360
rect 134120 27360 134280 27520
rect 134120 27520 134280 27680
rect 134120 27680 134280 27840
rect 134120 27840 134280 28000
rect 134120 28000 134280 28160
rect 134120 28160 134280 28320
rect 134120 28320 134280 28480
rect 134120 28480 134280 28640
rect 134120 28640 134280 28800
rect 134120 28800 134280 28960
rect 134120 28960 134280 29120
rect 134120 29120 134280 29280
rect 134120 29280 134280 29440
rect 134120 29440 134280 29600
rect 134120 29600 134280 29760
rect 134120 29760 134280 29920
rect 134120 29920 134280 30080
rect 134120 49760 134280 49920
rect 134120 49920 134280 50080
rect 134120 50080 134280 50240
rect 134120 50240 134280 50400
rect 134120 50400 134280 50560
rect 134120 50560 134280 50720
rect 134120 50720 134280 50880
rect 134120 50880 134280 51040
rect 134120 51040 134280 51200
rect 134120 51200 134280 51360
rect 134120 51360 134280 51520
rect 134120 51520 134280 51680
rect 134120 51680 134280 51840
rect 134120 51840 134280 52000
rect 134120 52000 134280 52160
rect 134120 52160 134280 52320
rect 134120 52320 134280 52480
rect 134120 52480 134280 52640
rect 134120 52640 134280 52800
rect 134120 52800 134280 52960
rect 134120 52960 134280 53120
rect 134120 53120 134280 53280
rect 134280 26720 134440 26880
rect 134280 26880 134440 27040
rect 134280 27040 134440 27200
rect 134280 27200 134440 27360
rect 134280 27360 134440 27520
rect 134280 27520 134440 27680
rect 134280 27680 134440 27840
rect 134280 27840 134440 28000
rect 134280 28000 134440 28160
rect 134280 28160 134440 28320
rect 134280 28320 134440 28480
rect 134280 28480 134440 28640
rect 134280 28640 134440 28800
rect 134280 28800 134440 28960
rect 134280 28960 134440 29120
rect 134280 29120 134440 29280
rect 134280 29280 134440 29440
rect 134280 29440 134440 29600
rect 134280 29600 134440 29760
rect 134280 29760 134440 29920
rect 134280 29920 134440 30080
rect 134280 30080 134440 30240
rect 134280 49760 134440 49920
rect 134280 49920 134440 50080
rect 134280 50080 134440 50240
rect 134280 50240 134440 50400
rect 134280 50400 134440 50560
rect 134280 50560 134440 50720
rect 134280 50720 134440 50880
rect 134280 50880 134440 51040
rect 134280 51040 134440 51200
rect 134280 51200 134440 51360
rect 134280 51360 134440 51520
rect 134280 51520 134440 51680
rect 134280 51680 134440 51840
rect 134280 51840 134440 52000
rect 134280 52000 134440 52160
rect 134280 52160 134440 52320
rect 134280 52320 134440 52480
rect 134280 52480 134440 52640
rect 134280 52640 134440 52800
rect 134280 52800 134440 52960
rect 134280 52960 134440 53120
rect 134280 53120 134440 53280
rect 134440 26720 134600 26880
rect 134440 26880 134600 27040
rect 134440 27040 134600 27200
rect 134440 27200 134600 27360
rect 134440 27360 134600 27520
rect 134440 27520 134600 27680
rect 134440 27680 134600 27840
rect 134440 27840 134600 28000
rect 134440 28000 134600 28160
rect 134440 28160 134600 28320
rect 134440 28320 134600 28480
rect 134440 28480 134600 28640
rect 134440 28640 134600 28800
rect 134440 28800 134600 28960
rect 134440 28960 134600 29120
rect 134440 29120 134600 29280
rect 134440 29280 134600 29440
rect 134440 29440 134600 29600
rect 134440 29600 134600 29760
rect 134440 29760 134600 29920
rect 134440 29920 134600 30080
rect 134440 30080 134600 30240
rect 134440 49760 134600 49920
rect 134440 49920 134600 50080
rect 134440 50080 134600 50240
rect 134440 50240 134600 50400
rect 134440 50400 134600 50560
rect 134440 50560 134600 50720
rect 134440 50720 134600 50880
rect 134440 50880 134600 51040
rect 134440 51040 134600 51200
rect 134440 51200 134600 51360
rect 134440 51360 134600 51520
rect 134440 51520 134600 51680
rect 134440 51680 134600 51840
rect 134440 51840 134600 52000
rect 134440 52000 134600 52160
rect 134440 52160 134600 52320
rect 134440 52320 134600 52480
rect 134440 52480 134600 52640
rect 134440 52640 134600 52800
rect 134440 52800 134600 52960
rect 134440 52960 134600 53120
rect 134440 53120 134600 53280
rect 134600 26720 134760 26880
rect 134600 26880 134760 27040
rect 134600 27040 134760 27200
rect 134600 27200 134760 27360
rect 134600 27360 134760 27520
rect 134600 27520 134760 27680
rect 134600 27680 134760 27840
rect 134600 27840 134760 28000
rect 134600 28000 134760 28160
rect 134600 28160 134760 28320
rect 134600 28320 134760 28480
rect 134600 28480 134760 28640
rect 134600 28640 134760 28800
rect 134600 28800 134760 28960
rect 134600 28960 134760 29120
rect 134600 29120 134760 29280
rect 134600 29280 134760 29440
rect 134600 29440 134760 29600
rect 134600 29600 134760 29760
rect 134600 29760 134760 29920
rect 134600 29920 134760 30080
rect 134600 30080 134760 30240
rect 134600 49920 134760 50080
rect 134600 50080 134760 50240
rect 134600 50240 134760 50400
rect 134600 50400 134760 50560
rect 134600 50560 134760 50720
rect 134600 50720 134760 50880
rect 134600 50880 134760 51040
rect 134600 51040 134760 51200
rect 134600 51200 134760 51360
rect 134600 51360 134760 51520
rect 134600 51520 134760 51680
rect 134600 51680 134760 51840
rect 134600 51840 134760 52000
rect 134600 52000 134760 52160
rect 134600 52160 134760 52320
rect 134600 52320 134760 52480
rect 134600 52480 134760 52640
rect 134600 52640 134760 52800
rect 134600 52800 134760 52960
rect 134600 52960 134760 53120
rect 134600 53120 134760 53280
rect 134760 26720 134920 26880
rect 134760 26880 134920 27040
rect 134760 27040 134920 27200
rect 134760 27200 134920 27360
rect 134760 27360 134920 27520
rect 134760 27520 134920 27680
rect 134760 27680 134920 27840
rect 134760 27840 134920 28000
rect 134760 28000 134920 28160
rect 134760 28160 134920 28320
rect 134760 28320 134920 28480
rect 134760 28480 134920 28640
rect 134760 28640 134920 28800
rect 134760 28800 134920 28960
rect 134760 28960 134920 29120
rect 134760 29120 134920 29280
rect 134760 29280 134920 29440
rect 134760 29440 134920 29600
rect 134760 29600 134920 29760
rect 134760 29760 134920 29920
rect 134760 29920 134920 30080
rect 134760 30080 134920 30240
rect 134760 49760 134920 49920
rect 134760 49920 134920 50080
rect 134760 50080 134920 50240
rect 134760 50240 134920 50400
rect 134760 50400 134920 50560
rect 134760 50560 134920 50720
rect 134760 50720 134920 50880
rect 134760 50880 134920 51040
rect 134760 51040 134920 51200
rect 134760 51200 134920 51360
rect 134760 51360 134920 51520
rect 134760 51520 134920 51680
rect 134760 51680 134920 51840
rect 134760 51840 134920 52000
rect 134760 52000 134920 52160
rect 134760 52160 134920 52320
rect 134760 52320 134920 52480
rect 134760 52480 134920 52640
rect 134760 52640 134920 52800
rect 134760 52800 134920 52960
rect 134760 52960 134920 53120
rect 134760 53120 134920 53280
rect 134920 26720 135080 26880
rect 134920 26880 135080 27040
rect 134920 27040 135080 27200
rect 134920 27200 135080 27360
rect 134920 27360 135080 27520
rect 134920 27520 135080 27680
rect 134920 27680 135080 27840
rect 134920 27840 135080 28000
rect 134920 28000 135080 28160
rect 134920 28160 135080 28320
rect 134920 28320 135080 28480
rect 134920 28480 135080 28640
rect 134920 28640 135080 28800
rect 134920 28800 135080 28960
rect 134920 28960 135080 29120
rect 134920 29120 135080 29280
rect 134920 29280 135080 29440
rect 134920 29440 135080 29600
rect 134920 29600 135080 29760
rect 134920 29760 135080 29920
rect 134920 29920 135080 30080
rect 134920 30080 135080 30240
rect 134920 30240 135080 30400
rect 134920 49920 135080 50080
rect 134920 50080 135080 50240
rect 134920 50240 135080 50400
rect 134920 50400 135080 50560
rect 134920 50560 135080 50720
rect 134920 50720 135080 50880
rect 134920 50880 135080 51040
rect 134920 51040 135080 51200
rect 134920 51200 135080 51360
rect 134920 51360 135080 51520
rect 134920 51520 135080 51680
rect 134920 51680 135080 51840
rect 134920 51840 135080 52000
rect 134920 52000 135080 52160
rect 134920 52160 135080 52320
rect 134920 52320 135080 52480
rect 134920 52480 135080 52640
rect 134920 52640 135080 52800
rect 134920 52800 135080 52960
rect 134920 52960 135080 53120
rect 134920 53120 135080 53280
rect 135080 26720 135240 26880
rect 135080 26880 135240 27040
rect 135080 27040 135240 27200
rect 135080 27200 135240 27360
rect 135080 27360 135240 27520
rect 135080 27520 135240 27680
rect 135080 27680 135240 27840
rect 135080 27840 135240 28000
rect 135080 28000 135240 28160
rect 135080 28160 135240 28320
rect 135080 28320 135240 28480
rect 135080 28480 135240 28640
rect 135080 28640 135240 28800
rect 135080 28800 135240 28960
rect 135080 28960 135240 29120
rect 135080 29120 135240 29280
rect 135080 29280 135240 29440
rect 135080 29440 135240 29600
rect 135080 29600 135240 29760
rect 135080 29760 135240 29920
rect 135080 29920 135240 30080
rect 135080 30080 135240 30240
rect 135080 30240 135240 30400
rect 135080 49760 135240 49920
rect 135080 49920 135240 50080
rect 135080 50080 135240 50240
rect 135080 50240 135240 50400
rect 135080 50400 135240 50560
rect 135080 50560 135240 50720
rect 135080 50720 135240 50880
rect 135080 50880 135240 51040
rect 135080 51040 135240 51200
rect 135080 51200 135240 51360
rect 135080 51360 135240 51520
rect 135080 51520 135240 51680
rect 135080 51680 135240 51840
rect 135080 51840 135240 52000
rect 135080 52000 135240 52160
rect 135080 52160 135240 52320
rect 135080 52320 135240 52480
rect 135080 52480 135240 52640
rect 135080 52640 135240 52800
rect 135080 52800 135240 52960
rect 135080 52960 135240 53120
rect 135080 53120 135240 53280
rect 135240 26880 135400 27040
rect 135240 27040 135400 27200
rect 135240 27200 135400 27360
rect 135240 27360 135400 27520
rect 135240 27520 135400 27680
rect 135240 27680 135400 27840
rect 135240 27840 135400 28000
rect 135240 28000 135400 28160
rect 135240 28160 135400 28320
rect 135240 28320 135400 28480
rect 135240 28480 135400 28640
rect 135240 28640 135400 28800
rect 135240 28800 135400 28960
rect 135240 28960 135400 29120
rect 135240 29120 135400 29280
rect 135240 29280 135400 29440
rect 135240 29440 135400 29600
rect 135240 29600 135400 29760
rect 135240 29760 135400 29920
rect 135240 29920 135400 30080
rect 135240 30080 135400 30240
rect 135240 30240 135400 30400
rect 135240 49760 135400 49920
rect 135240 49920 135400 50080
rect 135240 50080 135400 50240
rect 135240 50240 135400 50400
rect 135240 50400 135400 50560
rect 135240 50560 135400 50720
rect 135240 50720 135400 50880
rect 135240 50880 135400 51040
rect 135240 51040 135400 51200
rect 135240 51200 135400 51360
rect 135240 51360 135400 51520
rect 135240 51520 135400 51680
rect 135240 51680 135400 51840
rect 135240 51840 135400 52000
rect 135240 52000 135400 52160
rect 135240 52160 135400 52320
rect 135240 52320 135400 52480
rect 135240 52480 135400 52640
rect 135240 52640 135400 52800
rect 135240 52800 135400 52960
rect 135240 52960 135400 53120
rect 135240 53120 135400 53280
rect 135400 26880 135560 27040
rect 135400 27040 135560 27200
rect 135400 27200 135560 27360
rect 135400 27360 135560 27520
rect 135400 27520 135560 27680
rect 135400 27680 135560 27840
rect 135400 27840 135560 28000
rect 135400 28000 135560 28160
rect 135400 28160 135560 28320
rect 135400 28320 135560 28480
rect 135400 28480 135560 28640
rect 135400 28640 135560 28800
rect 135400 28800 135560 28960
rect 135400 28960 135560 29120
rect 135400 29120 135560 29280
rect 135400 29280 135560 29440
rect 135400 29440 135560 29600
rect 135400 29600 135560 29760
rect 135400 29760 135560 29920
rect 135400 29920 135560 30080
rect 135400 30080 135560 30240
rect 135400 30240 135560 30400
rect 135400 30400 135560 30560
rect 135400 49920 135560 50080
rect 135400 50080 135560 50240
rect 135400 50240 135560 50400
rect 135400 50400 135560 50560
rect 135400 50560 135560 50720
rect 135400 50720 135560 50880
rect 135400 50880 135560 51040
rect 135400 51040 135560 51200
rect 135400 51200 135560 51360
rect 135400 51360 135560 51520
rect 135400 51520 135560 51680
rect 135400 51680 135560 51840
rect 135400 51840 135560 52000
rect 135400 52000 135560 52160
rect 135400 52160 135560 52320
rect 135400 52320 135560 52480
rect 135400 52480 135560 52640
rect 135400 52640 135560 52800
rect 135400 52800 135560 52960
rect 135400 52960 135560 53120
rect 135400 53120 135560 53280
rect 135560 26880 135720 27040
rect 135560 27040 135720 27200
rect 135560 27200 135720 27360
rect 135560 27360 135720 27520
rect 135560 27520 135720 27680
rect 135560 27680 135720 27840
rect 135560 27840 135720 28000
rect 135560 28000 135720 28160
rect 135560 28160 135720 28320
rect 135560 28320 135720 28480
rect 135560 28480 135720 28640
rect 135560 28640 135720 28800
rect 135560 28800 135720 28960
rect 135560 28960 135720 29120
rect 135560 29120 135720 29280
rect 135560 29280 135720 29440
rect 135560 29440 135720 29600
rect 135560 29600 135720 29760
rect 135560 29760 135720 29920
rect 135560 29920 135720 30080
rect 135560 30080 135720 30240
rect 135560 30240 135720 30400
rect 135560 30400 135720 30560
rect 135560 49760 135720 49920
rect 135560 49920 135720 50080
rect 135560 50080 135720 50240
rect 135560 50240 135720 50400
rect 135560 50400 135720 50560
rect 135560 50560 135720 50720
rect 135560 50720 135720 50880
rect 135560 50880 135720 51040
rect 135560 51040 135720 51200
rect 135560 51200 135720 51360
rect 135560 51360 135720 51520
rect 135560 51520 135720 51680
rect 135560 51680 135720 51840
rect 135560 51840 135720 52000
rect 135560 52000 135720 52160
rect 135560 52160 135720 52320
rect 135560 52320 135720 52480
rect 135560 52480 135720 52640
rect 135560 52640 135720 52800
rect 135560 52800 135720 52960
rect 135560 52960 135720 53120
rect 135560 53120 135720 53280
rect 135720 26880 135880 27040
rect 135720 27040 135880 27200
rect 135720 27200 135880 27360
rect 135720 27360 135880 27520
rect 135720 27520 135880 27680
rect 135720 27680 135880 27840
rect 135720 27840 135880 28000
rect 135720 28000 135880 28160
rect 135720 28160 135880 28320
rect 135720 28320 135880 28480
rect 135720 28480 135880 28640
rect 135720 28640 135880 28800
rect 135720 28800 135880 28960
rect 135720 28960 135880 29120
rect 135720 29120 135880 29280
rect 135720 29280 135880 29440
rect 135720 29440 135880 29600
rect 135720 29600 135880 29760
rect 135720 29760 135880 29920
rect 135720 29920 135880 30080
rect 135720 30080 135880 30240
rect 135720 30240 135880 30400
rect 135720 30400 135880 30560
rect 135720 49760 135880 49920
rect 135720 49920 135880 50080
rect 135720 50080 135880 50240
rect 135720 50240 135880 50400
rect 135720 50400 135880 50560
rect 135720 50560 135880 50720
rect 135720 50720 135880 50880
rect 135720 50880 135880 51040
rect 135720 51040 135880 51200
rect 135720 51200 135880 51360
rect 135720 51360 135880 51520
rect 135720 51520 135880 51680
rect 135720 51680 135880 51840
rect 135720 51840 135880 52000
rect 135720 52000 135880 52160
rect 135720 52160 135880 52320
rect 135720 52320 135880 52480
rect 135720 52480 135880 52640
rect 135720 52640 135880 52800
rect 135720 52800 135880 52960
rect 135720 52960 135880 53120
rect 135720 53120 135880 53280
rect 135880 27040 136040 27200
rect 135880 27200 136040 27360
rect 135880 27360 136040 27520
rect 135880 27520 136040 27680
rect 135880 27680 136040 27840
rect 135880 27840 136040 28000
rect 135880 28000 136040 28160
rect 135880 28160 136040 28320
rect 135880 28320 136040 28480
rect 135880 28480 136040 28640
rect 135880 28640 136040 28800
rect 135880 28800 136040 28960
rect 135880 28960 136040 29120
rect 135880 29120 136040 29280
rect 135880 29280 136040 29440
rect 135880 29440 136040 29600
rect 135880 29600 136040 29760
rect 135880 29760 136040 29920
rect 135880 29920 136040 30080
rect 135880 30080 136040 30240
rect 135880 30240 136040 30400
rect 135880 30400 136040 30560
rect 135880 30560 136040 30720
rect 135880 49760 136040 49920
rect 135880 49920 136040 50080
rect 135880 50080 136040 50240
rect 135880 50240 136040 50400
rect 135880 50400 136040 50560
rect 135880 50560 136040 50720
rect 135880 50720 136040 50880
rect 135880 50880 136040 51040
rect 135880 51040 136040 51200
rect 135880 51200 136040 51360
rect 135880 51360 136040 51520
rect 135880 51520 136040 51680
rect 135880 51680 136040 51840
rect 135880 51840 136040 52000
rect 135880 52000 136040 52160
rect 135880 52160 136040 52320
rect 135880 52320 136040 52480
rect 135880 52480 136040 52640
rect 135880 52640 136040 52800
rect 135880 52800 136040 52960
rect 135880 52960 136040 53120
rect 135880 53120 136040 53280
rect 136040 27040 136200 27200
rect 136040 27200 136200 27360
rect 136040 27360 136200 27520
rect 136040 27520 136200 27680
rect 136040 27680 136200 27840
rect 136040 27840 136200 28000
rect 136040 28000 136200 28160
rect 136040 28160 136200 28320
rect 136040 28320 136200 28480
rect 136040 28480 136200 28640
rect 136040 28640 136200 28800
rect 136040 28800 136200 28960
rect 136040 28960 136200 29120
rect 136040 29120 136200 29280
rect 136040 29280 136200 29440
rect 136040 29440 136200 29600
rect 136040 29600 136200 29760
rect 136040 29760 136200 29920
rect 136040 29920 136200 30080
rect 136040 30080 136200 30240
rect 136040 30240 136200 30400
rect 136040 30400 136200 30560
rect 136040 30560 136200 30720
rect 136040 49760 136200 49920
rect 136040 49920 136200 50080
rect 136040 50080 136200 50240
rect 136040 50240 136200 50400
rect 136040 50400 136200 50560
rect 136040 50560 136200 50720
rect 136040 50720 136200 50880
rect 136040 50880 136200 51040
rect 136040 51040 136200 51200
rect 136040 51200 136200 51360
rect 136040 51360 136200 51520
rect 136040 51520 136200 51680
rect 136040 51680 136200 51840
rect 136040 51840 136200 52000
rect 136040 52000 136200 52160
rect 136040 52160 136200 52320
rect 136040 52320 136200 52480
rect 136040 52480 136200 52640
rect 136040 52640 136200 52800
rect 136040 52800 136200 52960
rect 136040 52960 136200 53120
rect 136040 53120 136200 53280
rect 136200 27040 136360 27200
rect 136200 27200 136360 27360
rect 136200 27360 136360 27520
rect 136200 27520 136360 27680
rect 136200 27680 136360 27840
rect 136200 27840 136360 28000
rect 136200 28000 136360 28160
rect 136200 28160 136360 28320
rect 136200 28320 136360 28480
rect 136200 28480 136360 28640
rect 136200 28640 136360 28800
rect 136200 28800 136360 28960
rect 136200 28960 136360 29120
rect 136200 29120 136360 29280
rect 136200 29280 136360 29440
rect 136200 29440 136360 29600
rect 136200 29600 136360 29760
rect 136200 29760 136360 29920
rect 136200 29920 136360 30080
rect 136200 30080 136360 30240
rect 136200 30240 136360 30400
rect 136200 30400 136360 30560
rect 136200 30560 136360 30720
rect 136200 30720 136360 30880
rect 136200 49760 136360 49920
rect 136200 49920 136360 50080
rect 136200 50080 136360 50240
rect 136200 50240 136360 50400
rect 136200 50400 136360 50560
rect 136200 50560 136360 50720
rect 136200 50720 136360 50880
rect 136200 50880 136360 51040
rect 136200 51040 136360 51200
rect 136200 51200 136360 51360
rect 136200 51360 136360 51520
rect 136200 51520 136360 51680
rect 136200 51680 136360 51840
rect 136200 51840 136360 52000
rect 136200 52000 136360 52160
rect 136200 52160 136360 52320
rect 136200 52320 136360 52480
rect 136200 52480 136360 52640
rect 136200 52640 136360 52800
rect 136200 52800 136360 52960
rect 136200 52960 136360 53120
rect 136200 53120 136360 53280
rect 136360 27200 136520 27360
rect 136360 27360 136520 27520
rect 136360 27520 136520 27680
rect 136360 27680 136520 27840
rect 136360 27840 136520 28000
rect 136360 28000 136520 28160
rect 136360 28160 136520 28320
rect 136360 28320 136520 28480
rect 136360 28480 136520 28640
rect 136360 28640 136520 28800
rect 136360 28800 136520 28960
rect 136360 28960 136520 29120
rect 136360 29120 136520 29280
rect 136360 29280 136520 29440
rect 136360 29440 136520 29600
rect 136360 29600 136520 29760
rect 136360 29760 136520 29920
rect 136360 29920 136520 30080
rect 136360 30080 136520 30240
rect 136360 30240 136520 30400
rect 136360 30400 136520 30560
rect 136360 30560 136520 30720
rect 136360 30720 136520 30880
rect 136360 30880 136520 31040
rect 136360 49760 136520 49920
rect 136360 49920 136520 50080
rect 136360 50080 136520 50240
rect 136360 50240 136520 50400
rect 136360 50400 136520 50560
rect 136360 50560 136520 50720
rect 136360 50720 136520 50880
rect 136360 50880 136520 51040
rect 136360 51040 136520 51200
rect 136360 51200 136520 51360
rect 136360 51360 136520 51520
rect 136360 51520 136520 51680
rect 136360 51680 136520 51840
rect 136360 51840 136520 52000
rect 136360 52000 136520 52160
rect 136360 52160 136520 52320
rect 136360 52320 136520 52480
rect 136360 52480 136520 52640
rect 136360 52640 136520 52800
rect 136360 52800 136520 52960
rect 136360 52960 136520 53120
rect 136360 53120 136520 53280
rect 136520 27200 136680 27360
rect 136520 27360 136680 27520
rect 136520 27520 136680 27680
rect 136520 27680 136680 27840
rect 136520 27840 136680 28000
rect 136520 28000 136680 28160
rect 136520 28160 136680 28320
rect 136520 28320 136680 28480
rect 136520 28480 136680 28640
rect 136520 28640 136680 28800
rect 136520 28800 136680 28960
rect 136520 28960 136680 29120
rect 136520 29120 136680 29280
rect 136520 29280 136680 29440
rect 136520 29440 136680 29600
rect 136520 29600 136680 29760
rect 136520 29760 136680 29920
rect 136520 29920 136680 30080
rect 136520 30080 136680 30240
rect 136520 30240 136680 30400
rect 136520 30400 136680 30560
rect 136520 30560 136680 30720
rect 136520 30720 136680 30880
rect 136520 30880 136680 31040
rect 136520 49760 136680 49920
rect 136520 49920 136680 50080
rect 136520 50080 136680 50240
rect 136520 50240 136680 50400
rect 136520 50400 136680 50560
rect 136520 50560 136680 50720
rect 136520 50720 136680 50880
rect 136520 50880 136680 51040
rect 136520 51040 136680 51200
rect 136520 51200 136680 51360
rect 136520 51360 136680 51520
rect 136520 51520 136680 51680
rect 136520 51680 136680 51840
rect 136520 51840 136680 52000
rect 136520 52000 136680 52160
rect 136520 52160 136680 52320
rect 136520 52320 136680 52480
rect 136520 52480 136680 52640
rect 136520 52640 136680 52800
rect 136520 52800 136680 52960
rect 136520 52960 136680 53120
rect 136520 53120 136680 53280
rect 136680 27200 136840 27360
rect 136680 27360 136840 27520
rect 136680 27520 136840 27680
rect 136680 27680 136840 27840
rect 136680 27840 136840 28000
rect 136680 28000 136840 28160
rect 136680 28160 136840 28320
rect 136680 28320 136840 28480
rect 136680 28480 136840 28640
rect 136680 28640 136840 28800
rect 136680 28800 136840 28960
rect 136680 28960 136840 29120
rect 136680 29120 136840 29280
rect 136680 29280 136840 29440
rect 136680 29440 136840 29600
rect 136680 29600 136840 29760
rect 136680 29760 136840 29920
rect 136680 29920 136840 30080
rect 136680 30080 136840 30240
rect 136680 30240 136840 30400
rect 136680 30400 136840 30560
rect 136680 30560 136840 30720
rect 136680 30720 136840 30880
rect 136680 30880 136840 31040
rect 136680 31040 136840 31200
rect 136680 49600 136840 49760
rect 136680 49760 136840 49920
rect 136680 49920 136840 50080
rect 136680 50080 136840 50240
rect 136680 50240 136840 50400
rect 136680 50400 136840 50560
rect 136680 50560 136840 50720
rect 136680 50720 136840 50880
rect 136680 50880 136840 51040
rect 136680 51040 136840 51200
rect 136680 51200 136840 51360
rect 136680 51360 136840 51520
rect 136680 51520 136840 51680
rect 136680 51680 136840 51840
rect 136680 51840 136840 52000
rect 136680 52000 136840 52160
rect 136680 52160 136840 52320
rect 136680 52320 136840 52480
rect 136680 52480 136840 52640
rect 136680 52640 136840 52800
rect 136680 52800 136840 52960
rect 136680 52960 136840 53120
rect 136680 53120 136840 53280
rect 136840 27360 137000 27520
rect 136840 27520 137000 27680
rect 136840 27680 137000 27840
rect 136840 27840 137000 28000
rect 136840 28000 137000 28160
rect 136840 28160 137000 28320
rect 136840 28320 137000 28480
rect 136840 28480 137000 28640
rect 136840 28640 137000 28800
rect 136840 28800 137000 28960
rect 136840 28960 137000 29120
rect 136840 29120 137000 29280
rect 136840 29280 137000 29440
rect 136840 29440 137000 29600
rect 136840 29600 137000 29760
rect 136840 29760 137000 29920
rect 136840 29920 137000 30080
rect 136840 30080 137000 30240
rect 136840 30240 137000 30400
rect 136840 30400 137000 30560
rect 136840 30560 137000 30720
rect 136840 30720 137000 30880
rect 136840 30880 137000 31040
rect 136840 31040 137000 31200
rect 136840 31200 137000 31360
rect 136840 49600 137000 49760
rect 136840 49760 137000 49920
rect 136840 49920 137000 50080
rect 136840 50080 137000 50240
rect 136840 50240 137000 50400
rect 136840 50400 137000 50560
rect 136840 50560 137000 50720
rect 136840 50720 137000 50880
rect 136840 50880 137000 51040
rect 136840 51040 137000 51200
rect 136840 51200 137000 51360
rect 136840 51360 137000 51520
rect 136840 51520 137000 51680
rect 136840 51680 137000 51840
rect 136840 51840 137000 52000
rect 136840 52000 137000 52160
rect 136840 52160 137000 52320
rect 136840 52320 137000 52480
rect 136840 52480 137000 52640
rect 136840 52640 137000 52800
rect 136840 52800 137000 52960
rect 136840 52960 137000 53120
rect 137000 27360 137160 27520
rect 137000 27520 137160 27680
rect 137000 27680 137160 27840
rect 137000 27840 137160 28000
rect 137000 28000 137160 28160
rect 137000 28160 137160 28320
rect 137000 28320 137160 28480
rect 137000 28480 137160 28640
rect 137000 28640 137160 28800
rect 137000 28800 137160 28960
rect 137000 28960 137160 29120
rect 137000 29120 137160 29280
rect 137000 29280 137160 29440
rect 137000 29440 137160 29600
rect 137000 29600 137160 29760
rect 137000 29760 137160 29920
rect 137000 29920 137160 30080
rect 137000 30080 137160 30240
rect 137000 30240 137160 30400
rect 137000 30400 137160 30560
rect 137000 30560 137160 30720
rect 137000 30720 137160 30880
rect 137000 30880 137160 31040
rect 137000 31040 137160 31200
rect 137000 31200 137160 31360
rect 137000 49600 137160 49760
rect 137000 49760 137160 49920
rect 137000 49920 137160 50080
rect 137000 50080 137160 50240
rect 137000 50240 137160 50400
rect 137000 50400 137160 50560
rect 137000 50560 137160 50720
rect 137000 50720 137160 50880
rect 137000 50880 137160 51040
rect 137000 51040 137160 51200
rect 137000 51200 137160 51360
rect 137000 51360 137160 51520
rect 137000 51520 137160 51680
rect 137000 51680 137160 51840
rect 137000 51840 137160 52000
rect 137000 52000 137160 52160
rect 137000 52160 137160 52320
rect 137000 52320 137160 52480
rect 137000 52480 137160 52640
rect 137000 52640 137160 52800
rect 137000 52800 137160 52960
rect 137000 52960 137160 53120
rect 137160 27520 137320 27680
rect 137160 27680 137320 27840
rect 137160 27840 137320 28000
rect 137160 28000 137320 28160
rect 137160 28160 137320 28320
rect 137160 28320 137320 28480
rect 137160 28480 137320 28640
rect 137160 28640 137320 28800
rect 137160 28800 137320 28960
rect 137160 28960 137320 29120
rect 137160 29120 137320 29280
rect 137160 29280 137320 29440
rect 137160 29440 137320 29600
rect 137160 29600 137320 29760
rect 137160 29760 137320 29920
rect 137160 29920 137320 30080
rect 137160 30080 137320 30240
rect 137160 30240 137320 30400
rect 137160 30400 137320 30560
rect 137160 30560 137320 30720
rect 137160 30720 137320 30880
rect 137160 30880 137320 31040
rect 137160 31040 137320 31200
rect 137160 31200 137320 31360
rect 137160 31360 137320 31520
rect 137160 49600 137320 49760
rect 137160 49760 137320 49920
rect 137160 49920 137320 50080
rect 137160 50080 137320 50240
rect 137160 50240 137320 50400
rect 137160 50400 137320 50560
rect 137160 50560 137320 50720
rect 137160 50720 137320 50880
rect 137160 50880 137320 51040
rect 137160 51040 137320 51200
rect 137160 51200 137320 51360
rect 137160 51360 137320 51520
rect 137160 51520 137320 51680
rect 137160 51680 137320 51840
rect 137160 51840 137320 52000
rect 137160 52000 137320 52160
rect 137160 52160 137320 52320
rect 137160 52320 137320 52480
rect 137160 52480 137320 52640
rect 137160 52640 137320 52800
rect 137160 52800 137320 52960
rect 137160 52960 137320 53120
rect 137320 27520 137480 27680
rect 137320 27680 137480 27840
rect 137320 27840 137480 28000
rect 137320 28000 137480 28160
rect 137320 28160 137480 28320
rect 137320 28320 137480 28480
rect 137320 28480 137480 28640
rect 137320 28640 137480 28800
rect 137320 28800 137480 28960
rect 137320 28960 137480 29120
rect 137320 29120 137480 29280
rect 137320 29280 137480 29440
rect 137320 29440 137480 29600
rect 137320 29600 137480 29760
rect 137320 29760 137480 29920
rect 137320 29920 137480 30080
rect 137320 30080 137480 30240
rect 137320 30240 137480 30400
rect 137320 30400 137480 30560
rect 137320 30560 137480 30720
rect 137320 30720 137480 30880
rect 137320 30880 137480 31040
rect 137320 31040 137480 31200
rect 137320 31200 137480 31360
rect 137320 31360 137480 31520
rect 137320 31520 137480 31680
rect 137320 49440 137480 49600
rect 137320 49600 137480 49760
rect 137320 49760 137480 49920
rect 137320 49920 137480 50080
rect 137320 50080 137480 50240
rect 137320 50240 137480 50400
rect 137320 50400 137480 50560
rect 137320 50560 137480 50720
rect 137320 50720 137480 50880
rect 137320 50880 137480 51040
rect 137320 51040 137480 51200
rect 137320 51200 137480 51360
rect 137320 51360 137480 51520
rect 137320 51520 137480 51680
rect 137320 51680 137480 51840
rect 137320 51840 137480 52000
rect 137320 52000 137480 52160
rect 137320 52160 137480 52320
rect 137320 52320 137480 52480
rect 137320 52480 137480 52640
rect 137320 52640 137480 52800
rect 137320 52800 137480 52960
rect 137320 52960 137480 53120
rect 137480 27680 137640 27840
rect 137480 27840 137640 28000
rect 137480 28000 137640 28160
rect 137480 28160 137640 28320
rect 137480 28320 137640 28480
rect 137480 28480 137640 28640
rect 137480 28640 137640 28800
rect 137480 28800 137640 28960
rect 137480 28960 137640 29120
rect 137480 29120 137640 29280
rect 137480 29280 137640 29440
rect 137480 29440 137640 29600
rect 137480 29600 137640 29760
rect 137480 29760 137640 29920
rect 137480 29920 137640 30080
rect 137480 30080 137640 30240
rect 137480 30240 137640 30400
rect 137480 30400 137640 30560
rect 137480 30560 137640 30720
rect 137480 30720 137640 30880
rect 137480 30880 137640 31040
rect 137480 31040 137640 31200
rect 137480 31200 137640 31360
rect 137480 31360 137640 31520
rect 137480 31520 137640 31680
rect 137480 31680 137640 31840
rect 137480 49440 137640 49600
rect 137480 49600 137640 49760
rect 137480 49760 137640 49920
rect 137480 49920 137640 50080
rect 137480 50080 137640 50240
rect 137480 50240 137640 50400
rect 137480 50400 137640 50560
rect 137480 50560 137640 50720
rect 137480 50720 137640 50880
rect 137480 50880 137640 51040
rect 137480 51040 137640 51200
rect 137480 51200 137640 51360
rect 137480 51360 137640 51520
rect 137480 51520 137640 51680
rect 137480 51680 137640 51840
rect 137480 51840 137640 52000
rect 137480 52000 137640 52160
rect 137480 52160 137640 52320
rect 137480 52320 137640 52480
rect 137480 52480 137640 52640
rect 137480 52640 137640 52800
rect 137480 52800 137640 52960
rect 137480 52960 137640 53120
rect 137640 27680 137800 27840
rect 137640 27840 137800 28000
rect 137640 28000 137800 28160
rect 137640 28160 137800 28320
rect 137640 28320 137800 28480
rect 137640 28480 137800 28640
rect 137640 28640 137800 28800
rect 137640 28800 137800 28960
rect 137640 28960 137800 29120
rect 137640 29120 137800 29280
rect 137640 29280 137800 29440
rect 137640 29440 137800 29600
rect 137640 29600 137800 29760
rect 137640 29760 137800 29920
rect 137640 29920 137800 30080
rect 137640 30080 137800 30240
rect 137640 30240 137800 30400
rect 137640 30400 137800 30560
rect 137640 30560 137800 30720
rect 137640 30720 137800 30880
rect 137640 30880 137800 31040
rect 137640 31040 137800 31200
rect 137640 31200 137800 31360
rect 137640 31360 137800 31520
rect 137640 31520 137800 31680
rect 137640 31680 137800 31840
rect 137640 31840 137800 32000
rect 137640 49440 137800 49600
rect 137640 49600 137800 49760
rect 137640 49760 137800 49920
rect 137640 49920 137800 50080
rect 137640 50080 137800 50240
rect 137640 50240 137800 50400
rect 137640 50400 137800 50560
rect 137640 50560 137800 50720
rect 137640 50720 137800 50880
rect 137640 50880 137800 51040
rect 137640 51040 137800 51200
rect 137640 51200 137800 51360
rect 137640 51360 137800 51520
rect 137640 51520 137800 51680
rect 137640 51680 137800 51840
rect 137640 51840 137800 52000
rect 137640 52000 137800 52160
rect 137640 52160 137800 52320
rect 137640 52320 137800 52480
rect 137640 52480 137800 52640
rect 137640 52640 137800 52800
rect 137640 52800 137800 52960
rect 137640 52960 137800 53120
rect 137800 27840 137960 28000
rect 137800 28000 137960 28160
rect 137800 28160 137960 28320
rect 137800 28320 137960 28480
rect 137800 28480 137960 28640
rect 137800 28640 137960 28800
rect 137800 28800 137960 28960
rect 137800 28960 137960 29120
rect 137800 29120 137960 29280
rect 137800 29280 137960 29440
rect 137800 29440 137960 29600
rect 137800 29600 137960 29760
rect 137800 29760 137960 29920
rect 137800 29920 137960 30080
rect 137800 30080 137960 30240
rect 137800 30240 137960 30400
rect 137800 30400 137960 30560
rect 137800 30560 137960 30720
rect 137800 30720 137960 30880
rect 137800 30880 137960 31040
rect 137800 31040 137960 31200
rect 137800 31200 137960 31360
rect 137800 31360 137960 31520
rect 137800 31520 137960 31680
rect 137800 31680 137960 31840
rect 137800 31840 137960 32000
rect 137800 32000 137960 32160
rect 137800 49280 137960 49440
rect 137800 49440 137960 49600
rect 137800 49600 137960 49760
rect 137800 49760 137960 49920
rect 137800 49920 137960 50080
rect 137800 50080 137960 50240
rect 137800 50240 137960 50400
rect 137800 50400 137960 50560
rect 137800 50560 137960 50720
rect 137800 50720 137960 50880
rect 137800 50880 137960 51040
rect 137800 51040 137960 51200
rect 137800 51200 137960 51360
rect 137800 51360 137960 51520
rect 137800 51520 137960 51680
rect 137800 51680 137960 51840
rect 137800 51840 137960 52000
rect 137800 52000 137960 52160
rect 137800 52160 137960 52320
rect 137800 52320 137960 52480
rect 137800 52480 137960 52640
rect 137800 52640 137960 52800
rect 137800 52800 137960 52960
rect 137960 27840 138120 28000
rect 137960 28000 138120 28160
rect 137960 28160 138120 28320
rect 137960 28320 138120 28480
rect 137960 28480 138120 28640
rect 137960 28640 138120 28800
rect 137960 28800 138120 28960
rect 137960 28960 138120 29120
rect 137960 29120 138120 29280
rect 137960 29280 138120 29440
rect 137960 29440 138120 29600
rect 137960 29600 138120 29760
rect 137960 29760 138120 29920
rect 137960 29920 138120 30080
rect 137960 30080 138120 30240
rect 137960 30240 138120 30400
rect 137960 30400 138120 30560
rect 137960 30560 138120 30720
rect 137960 30720 138120 30880
rect 137960 30880 138120 31040
rect 137960 31040 138120 31200
rect 137960 31200 138120 31360
rect 137960 31360 138120 31520
rect 137960 31520 138120 31680
rect 137960 31680 138120 31840
rect 137960 31840 138120 32000
rect 137960 32000 138120 32160
rect 137960 32160 138120 32320
rect 137960 49280 138120 49440
rect 137960 49440 138120 49600
rect 137960 49600 138120 49760
rect 137960 49760 138120 49920
rect 137960 49920 138120 50080
rect 137960 50080 138120 50240
rect 137960 50240 138120 50400
rect 137960 50400 138120 50560
rect 137960 50560 138120 50720
rect 137960 50720 138120 50880
rect 137960 50880 138120 51040
rect 137960 51040 138120 51200
rect 137960 51200 138120 51360
rect 137960 51360 138120 51520
rect 137960 51520 138120 51680
rect 137960 51680 138120 51840
rect 137960 51840 138120 52000
rect 137960 52000 138120 52160
rect 137960 52160 138120 52320
rect 137960 52320 138120 52480
rect 137960 52480 138120 52640
rect 137960 52640 138120 52800
rect 137960 52800 138120 52960
rect 138120 28000 138280 28160
rect 138120 28160 138280 28320
rect 138120 28320 138280 28480
rect 138120 28480 138280 28640
rect 138120 28640 138280 28800
rect 138120 28800 138280 28960
rect 138120 28960 138280 29120
rect 138120 29120 138280 29280
rect 138120 29280 138280 29440
rect 138120 29440 138280 29600
rect 138120 29600 138280 29760
rect 138120 29760 138280 29920
rect 138120 29920 138280 30080
rect 138120 30080 138280 30240
rect 138120 30240 138280 30400
rect 138120 30400 138280 30560
rect 138120 30560 138280 30720
rect 138120 30720 138280 30880
rect 138120 30880 138280 31040
rect 138120 31040 138280 31200
rect 138120 31200 138280 31360
rect 138120 31360 138280 31520
rect 138120 31520 138280 31680
rect 138120 31680 138280 31840
rect 138120 31840 138280 32000
rect 138120 32000 138280 32160
rect 138120 32160 138280 32320
rect 138120 32320 138280 32480
rect 138120 49120 138280 49280
rect 138120 49280 138280 49440
rect 138120 49440 138280 49600
rect 138120 49600 138280 49760
rect 138120 49760 138280 49920
rect 138120 49920 138280 50080
rect 138120 50080 138280 50240
rect 138120 50240 138280 50400
rect 138120 50400 138280 50560
rect 138120 50560 138280 50720
rect 138120 50720 138280 50880
rect 138120 50880 138280 51040
rect 138120 51040 138280 51200
rect 138120 51200 138280 51360
rect 138120 51360 138280 51520
rect 138120 51520 138280 51680
rect 138120 51680 138280 51840
rect 138120 51840 138280 52000
rect 138120 52000 138280 52160
rect 138120 52160 138280 52320
rect 138120 52320 138280 52480
rect 138120 52480 138280 52640
rect 138120 52640 138280 52800
rect 138120 52800 138280 52960
rect 138280 28160 138440 28320
rect 138280 28320 138440 28480
rect 138280 28480 138440 28640
rect 138280 28640 138440 28800
rect 138280 28800 138440 28960
rect 138280 28960 138440 29120
rect 138280 29120 138440 29280
rect 138280 29280 138440 29440
rect 138280 29440 138440 29600
rect 138280 29600 138440 29760
rect 138280 29760 138440 29920
rect 138280 29920 138440 30080
rect 138280 30080 138440 30240
rect 138280 30240 138440 30400
rect 138280 30400 138440 30560
rect 138280 30560 138440 30720
rect 138280 30720 138440 30880
rect 138280 30880 138440 31040
rect 138280 31040 138440 31200
rect 138280 31200 138440 31360
rect 138280 31360 138440 31520
rect 138280 31520 138440 31680
rect 138280 31680 138440 31840
rect 138280 31840 138440 32000
rect 138280 32000 138440 32160
rect 138280 32160 138440 32320
rect 138280 32320 138440 32480
rect 138280 32480 138440 32640
rect 138280 48960 138440 49120
rect 138280 49120 138440 49280
rect 138280 49280 138440 49440
rect 138280 49440 138440 49600
rect 138280 49600 138440 49760
rect 138280 49760 138440 49920
rect 138280 49920 138440 50080
rect 138280 50080 138440 50240
rect 138280 50240 138440 50400
rect 138280 50400 138440 50560
rect 138280 50560 138440 50720
rect 138280 50720 138440 50880
rect 138280 50880 138440 51040
rect 138280 51040 138440 51200
rect 138280 51200 138440 51360
rect 138280 51360 138440 51520
rect 138280 51520 138440 51680
rect 138280 51680 138440 51840
rect 138280 51840 138440 52000
rect 138280 52000 138440 52160
rect 138280 52160 138440 52320
rect 138280 52320 138440 52480
rect 138280 52480 138440 52640
rect 138280 52640 138440 52800
rect 138440 28160 138600 28320
rect 138440 28320 138600 28480
rect 138440 28480 138600 28640
rect 138440 28640 138600 28800
rect 138440 28800 138600 28960
rect 138440 28960 138600 29120
rect 138440 29120 138600 29280
rect 138440 29280 138600 29440
rect 138440 29440 138600 29600
rect 138440 29600 138600 29760
rect 138440 29760 138600 29920
rect 138440 29920 138600 30080
rect 138440 30080 138600 30240
rect 138440 30240 138600 30400
rect 138440 30400 138600 30560
rect 138440 30560 138600 30720
rect 138440 30720 138600 30880
rect 138440 30880 138600 31040
rect 138440 31040 138600 31200
rect 138440 31200 138600 31360
rect 138440 31360 138600 31520
rect 138440 31520 138600 31680
rect 138440 31680 138600 31840
rect 138440 31840 138600 32000
rect 138440 32000 138600 32160
rect 138440 32160 138600 32320
rect 138440 32320 138600 32480
rect 138440 32480 138600 32640
rect 138440 32640 138600 32800
rect 138440 32800 138600 32960
rect 138440 48960 138600 49120
rect 138440 49120 138600 49280
rect 138440 49280 138600 49440
rect 138440 49440 138600 49600
rect 138440 49600 138600 49760
rect 138440 49760 138600 49920
rect 138440 49920 138600 50080
rect 138440 50080 138600 50240
rect 138440 50240 138600 50400
rect 138440 50400 138600 50560
rect 138440 50560 138600 50720
rect 138440 50720 138600 50880
rect 138440 50880 138600 51040
rect 138440 51040 138600 51200
rect 138440 51200 138600 51360
rect 138440 51360 138600 51520
rect 138440 51520 138600 51680
rect 138440 51680 138600 51840
rect 138440 51840 138600 52000
rect 138440 52000 138600 52160
rect 138440 52160 138600 52320
rect 138440 52320 138600 52480
rect 138440 52480 138600 52640
rect 138440 52640 138600 52800
rect 138600 28320 138760 28480
rect 138600 28480 138760 28640
rect 138600 28640 138760 28800
rect 138600 28800 138760 28960
rect 138600 28960 138760 29120
rect 138600 29120 138760 29280
rect 138600 29280 138760 29440
rect 138600 29440 138760 29600
rect 138600 29600 138760 29760
rect 138600 29760 138760 29920
rect 138600 29920 138760 30080
rect 138600 30080 138760 30240
rect 138600 30240 138760 30400
rect 138600 30400 138760 30560
rect 138600 30560 138760 30720
rect 138600 30720 138760 30880
rect 138600 30880 138760 31040
rect 138600 31040 138760 31200
rect 138600 31200 138760 31360
rect 138600 31360 138760 31520
rect 138600 31520 138760 31680
rect 138600 31680 138760 31840
rect 138600 31840 138760 32000
rect 138600 32000 138760 32160
rect 138600 32160 138760 32320
rect 138600 32320 138760 32480
rect 138600 32480 138760 32640
rect 138600 32640 138760 32800
rect 138600 32800 138760 32960
rect 138600 32960 138760 33120
rect 138600 48800 138760 48960
rect 138600 48960 138760 49120
rect 138600 49120 138760 49280
rect 138600 49280 138760 49440
rect 138600 49440 138760 49600
rect 138600 49600 138760 49760
rect 138600 49760 138760 49920
rect 138600 49920 138760 50080
rect 138600 50080 138760 50240
rect 138600 50240 138760 50400
rect 138600 50400 138760 50560
rect 138600 50560 138760 50720
rect 138600 50720 138760 50880
rect 138600 50880 138760 51040
rect 138600 51040 138760 51200
rect 138600 51200 138760 51360
rect 138600 51360 138760 51520
rect 138600 51520 138760 51680
rect 138600 51680 138760 51840
rect 138600 51840 138760 52000
rect 138600 52000 138760 52160
rect 138600 52160 138760 52320
rect 138600 52320 138760 52480
rect 138600 52480 138760 52640
rect 138600 52640 138760 52800
rect 138760 28480 138920 28640
rect 138760 28640 138920 28800
rect 138760 28800 138920 28960
rect 138760 28960 138920 29120
rect 138760 29120 138920 29280
rect 138760 29280 138920 29440
rect 138760 29440 138920 29600
rect 138760 29600 138920 29760
rect 138760 29760 138920 29920
rect 138760 29920 138920 30080
rect 138760 30080 138920 30240
rect 138760 30240 138920 30400
rect 138760 30400 138920 30560
rect 138760 30560 138920 30720
rect 138760 30720 138920 30880
rect 138760 30880 138920 31040
rect 138760 31040 138920 31200
rect 138760 31200 138920 31360
rect 138760 31360 138920 31520
rect 138760 31520 138920 31680
rect 138760 31680 138920 31840
rect 138760 31840 138920 32000
rect 138760 32000 138920 32160
rect 138760 32160 138920 32320
rect 138760 32320 138920 32480
rect 138760 32480 138920 32640
rect 138760 32640 138920 32800
rect 138760 32800 138920 32960
rect 138760 32960 138920 33120
rect 138760 33120 138920 33280
rect 138760 33280 138920 33440
rect 138760 48640 138920 48800
rect 138760 48800 138920 48960
rect 138760 48960 138920 49120
rect 138760 49120 138920 49280
rect 138760 49280 138920 49440
rect 138760 49440 138920 49600
rect 138760 49600 138920 49760
rect 138760 49760 138920 49920
rect 138760 49920 138920 50080
rect 138760 50080 138920 50240
rect 138760 50240 138920 50400
rect 138760 50400 138920 50560
rect 138760 50560 138920 50720
rect 138760 50720 138920 50880
rect 138760 50880 138920 51040
rect 138760 51040 138920 51200
rect 138760 51200 138920 51360
rect 138760 51360 138920 51520
rect 138760 51520 138920 51680
rect 138760 51680 138920 51840
rect 138760 51840 138920 52000
rect 138760 52000 138920 52160
rect 138760 52160 138920 52320
rect 138760 52320 138920 52480
rect 138760 52480 138920 52640
rect 138920 28640 139080 28800
rect 138920 28800 139080 28960
rect 138920 28960 139080 29120
rect 138920 29120 139080 29280
rect 138920 29280 139080 29440
rect 138920 29440 139080 29600
rect 138920 29600 139080 29760
rect 138920 29760 139080 29920
rect 138920 29920 139080 30080
rect 138920 30080 139080 30240
rect 138920 30240 139080 30400
rect 138920 30400 139080 30560
rect 138920 30560 139080 30720
rect 138920 30720 139080 30880
rect 138920 30880 139080 31040
rect 138920 31040 139080 31200
rect 138920 31200 139080 31360
rect 138920 31360 139080 31520
rect 138920 31520 139080 31680
rect 138920 31680 139080 31840
rect 138920 31840 139080 32000
rect 138920 32000 139080 32160
rect 138920 32160 139080 32320
rect 138920 32320 139080 32480
rect 138920 32480 139080 32640
rect 138920 32640 139080 32800
rect 138920 32800 139080 32960
rect 138920 32960 139080 33120
rect 138920 33120 139080 33280
rect 138920 33280 139080 33440
rect 138920 33440 139080 33600
rect 138920 48480 139080 48640
rect 138920 48640 139080 48800
rect 138920 48800 139080 48960
rect 138920 48960 139080 49120
rect 138920 49120 139080 49280
rect 138920 49280 139080 49440
rect 138920 49440 139080 49600
rect 138920 49600 139080 49760
rect 138920 49760 139080 49920
rect 138920 49920 139080 50080
rect 138920 50080 139080 50240
rect 138920 50240 139080 50400
rect 138920 50400 139080 50560
rect 138920 50560 139080 50720
rect 138920 50720 139080 50880
rect 138920 50880 139080 51040
rect 138920 51040 139080 51200
rect 138920 51200 139080 51360
rect 138920 51360 139080 51520
rect 138920 51520 139080 51680
rect 138920 51680 139080 51840
rect 138920 51840 139080 52000
rect 138920 52000 139080 52160
rect 138920 52160 139080 52320
rect 138920 52320 139080 52480
rect 138920 52480 139080 52640
rect 139080 28640 139240 28800
rect 139080 28800 139240 28960
rect 139080 28960 139240 29120
rect 139080 29120 139240 29280
rect 139080 29280 139240 29440
rect 139080 29440 139240 29600
rect 139080 29600 139240 29760
rect 139080 29760 139240 29920
rect 139080 29920 139240 30080
rect 139080 30080 139240 30240
rect 139080 30240 139240 30400
rect 139080 30400 139240 30560
rect 139080 30560 139240 30720
rect 139080 30720 139240 30880
rect 139080 30880 139240 31040
rect 139080 31040 139240 31200
rect 139080 31200 139240 31360
rect 139080 31360 139240 31520
rect 139080 31520 139240 31680
rect 139080 31680 139240 31840
rect 139080 31840 139240 32000
rect 139080 32000 139240 32160
rect 139080 32160 139240 32320
rect 139080 32320 139240 32480
rect 139080 32480 139240 32640
rect 139080 32640 139240 32800
rect 139080 32800 139240 32960
rect 139080 32960 139240 33120
rect 139080 33120 139240 33280
rect 139080 33280 139240 33440
rect 139080 33440 139240 33600
rect 139080 33600 139240 33760
rect 139080 33760 139240 33920
rect 139080 48320 139240 48480
rect 139080 48480 139240 48640
rect 139080 48640 139240 48800
rect 139080 48800 139240 48960
rect 139080 48960 139240 49120
rect 139080 49120 139240 49280
rect 139080 49280 139240 49440
rect 139080 49440 139240 49600
rect 139080 49600 139240 49760
rect 139080 49760 139240 49920
rect 139080 49920 139240 50080
rect 139080 50080 139240 50240
rect 139080 50240 139240 50400
rect 139080 50400 139240 50560
rect 139080 50560 139240 50720
rect 139080 50720 139240 50880
rect 139080 50880 139240 51040
rect 139080 51040 139240 51200
rect 139080 51200 139240 51360
rect 139080 51360 139240 51520
rect 139080 51520 139240 51680
rect 139080 51680 139240 51840
rect 139080 51840 139240 52000
rect 139080 52000 139240 52160
rect 139080 52160 139240 52320
rect 139080 52320 139240 52480
rect 139240 28800 139400 28960
rect 139240 28960 139400 29120
rect 139240 29120 139400 29280
rect 139240 29280 139400 29440
rect 139240 29440 139400 29600
rect 139240 29600 139400 29760
rect 139240 29760 139400 29920
rect 139240 29920 139400 30080
rect 139240 30080 139400 30240
rect 139240 30240 139400 30400
rect 139240 30400 139400 30560
rect 139240 30560 139400 30720
rect 139240 30720 139400 30880
rect 139240 30880 139400 31040
rect 139240 31040 139400 31200
rect 139240 31200 139400 31360
rect 139240 31360 139400 31520
rect 139240 31520 139400 31680
rect 139240 31680 139400 31840
rect 139240 31840 139400 32000
rect 139240 32000 139400 32160
rect 139240 32160 139400 32320
rect 139240 32320 139400 32480
rect 139240 32480 139400 32640
rect 139240 32640 139400 32800
rect 139240 32800 139400 32960
rect 139240 32960 139400 33120
rect 139240 33120 139400 33280
rect 139240 33280 139400 33440
rect 139240 33440 139400 33600
rect 139240 33600 139400 33760
rect 139240 33760 139400 33920
rect 139240 33920 139400 34080
rect 139240 34080 139400 34240
rect 139240 48160 139400 48320
rect 139240 48320 139400 48480
rect 139240 48480 139400 48640
rect 139240 48640 139400 48800
rect 139240 48800 139400 48960
rect 139240 48960 139400 49120
rect 139240 49120 139400 49280
rect 139240 49280 139400 49440
rect 139240 49440 139400 49600
rect 139240 49600 139400 49760
rect 139240 49760 139400 49920
rect 139240 49920 139400 50080
rect 139240 50080 139400 50240
rect 139240 50240 139400 50400
rect 139240 50400 139400 50560
rect 139240 50560 139400 50720
rect 139240 50720 139400 50880
rect 139240 50880 139400 51040
rect 139240 51040 139400 51200
rect 139240 51200 139400 51360
rect 139240 51360 139400 51520
rect 139240 51520 139400 51680
rect 139240 51680 139400 51840
rect 139240 51840 139400 52000
rect 139240 52000 139400 52160
rect 139240 52160 139400 52320
rect 139240 52320 139400 52480
rect 139400 28960 139560 29120
rect 139400 29120 139560 29280
rect 139400 29280 139560 29440
rect 139400 29440 139560 29600
rect 139400 29600 139560 29760
rect 139400 29760 139560 29920
rect 139400 29920 139560 30080
rect 139400 30080 139560 30240
rect 139400 30240 139560 30400
rect 139400 30400 139560 30560
rect 139400 30560 139560 30720
rect 139400 30720 139560 30880
rect 139400 30880 139560 31040
rect 139400 31040 139560 31200
rect 139400 31200 139560 31360
rect 139400 31360 139560 31520
rect 139400 31520 139560 31680
rect 139400 31680 139560 31840
rect 139400 31840 139560 32000
rect 139400 32000 139560 32160
rect 139400 32160 139560 32320
rect 139400 32320 139560 32480
rect 139400 32480 139560 32640
rect 139400 32640 139560 32800
rect 139400 32800 139560 32960
rect 139400 32960 139560 33120
rect 139400 33120 139560 33280
rect 139400 33280 139560 33440
rect 139400 33440 139560 33600
rect 139400 33600 139560 33760
rect 139400 33760 139560 33920
rect 139400 33920 139560 34080
rect 139400 34080 139560 34240
rect 139400 34240 139560 34400
rect 139400 34400 139560 34560
rect 139400 47840 139560 48000
rect 139400 48000 139560 48160
rect 139400 48160 139560 48320
rect 139400 48320 139560 48480
rect 139400 48480 139560 48640
rect 139400 48640 139560 48800
rect 139400 48800 139560 48960
rect 139400 48960 139560 49120
rect 139400 49120 139560 49280
rect 139400 49280 139560 49440
rect 139400 49440 139560 49600
rect 139400 49600 139560 49760
rect 139400 49760 139560 49920
rect 139400 49920 139560 50080
rect 139400 50080 139560 50240
rect 139400 50240 139560 50400
rect 139400 50400 139560 50560
rect 139400 50560 139560 50720
rect 139400 50720 139560 50880
rect 139400 50880 139560 51040
rect 139400 51040 139560 51200
rect 139400 51200 139560 51360
rect 139400 51360 139560 51520
rect 139400 51520 139560 51680
rect 139400 51680 139560 51840
rect 139400 51840 139560 52000
rect 139400 52000 139560 52160
rect 139400 52160 139560 52320
rect 139560 29120 139720 29280
rect 139560 29280 139720 29440
rect 139560 29440 139720 29600
rect 139560 29600 139720 29760
rect 139560 29760 139720 29920
rect 139560 29920 139720 30080
rect 139560 30080 139720 30240
rect 139560 30240 139720 30400
rect 139560 30400 139720 30560
rect 139560 30560 139720 30720
rect 139560 30720 139720 30880
rect 139560 30880 139720 31040
rect 139560 31040 139720 31200
rect 139560 31200 139720 31360
rect 139560 31360 139720 31520
rect 139560 31520 139720 31680
rect 139560 31680 139720 31840
rect 139560 31840 139720 32000
rect 139560 32000 139720 32160
rect 139560 32160 139720 32320
rect 139560 32320 139720 32480
rect 139560 32480 139720 32640
rect 139560 32640 139720 32800
rect 139560 32800 139720 32960
rect 139560 32960 139720 33120
rect 139560 33120 139720 33280
rect 139560 33280 139720 33440
rect 139560 33440 139720 33600
rect 139560 33600 139720 33760
rect 139560 33760 139720 33920
rect 139560 33920 139720 34080
rect 139560 34080 139720 34240
rect 139560 34240 139720 34400
rect 139560 34400 139720 34560
rect 139560 34560 139720 34720
rect 139560 34720 139720 34880
rect 139560 47680 139720 47840
rect 139560 47840 139720 48000
rect 139560 48000 139720 48160
rect 139560 48160 139720 48320
rect 139560 48320 139720 48480
rect 139560 48480 139720 48640
rect 139560 48640 139720 48800
rect 139560 48800 139720 48960
rect 139560 48960 139720 49120
rect 139560 49120 139720 49280
rect 139560 49280 139720 49440
rect 139560 49440 139720 49600
rect 139560 49600 139720 49760
rect 139560 49760 139720 49920
rect 139560 49920 139720 50080
rect 139560 50080 139720 50240
rect 139560 50240 139720 50400
rect 139560 50400 139720 50560
rect 139560 50560 139720 50720
rect 139560 50720 139720 50880
rect 139560 50880 139720 51040
rect 139560 51040 139720 51200
rect 139560 51200 139720 51360
rect 139560 51360 139720 51520
rect 139560 51520 139720 51680
rect 139560 51680 139720 51840
rect 139560 51840 139720 52000
rect 139560 52000 139720 52160
rect 139560 52160 139720 52320
rect 139720 29280 139880 29440
rect 139720 29440 139880 29600
rect 139720 29600 139880 29760
rect 139720 29760 139880 29920
rect 139720 29920 139880 30080
rect 139720 30080 139880 30240
rect 139720 30240 139880 30400
rect 139720 30400 139880 30560
rect 139720 30560 139880 30720
rect 139720 30720 139880 30880
rect 139720 30880 139880 31040
rect 139720 31040 139880 31200
rect 139720 31200 139880 31360
rect 139720 31360 139880 31520
rect 139720 31520 139880 31680
rect 139720 31680 139880 31840
rect 139720 31840 139880 32000
rect 139720 32000 139880 32160
rect 139720 32160 139880 32320
rect 139720 32320 139880 32480
rect 139720 32480 139880 32640
rect 139720 32640 139880 32800
rect 139720 32800 139880 32960
rect 139720 32960 139880 33120
rect 139720 33120 139880 33280
rect 139720 33280 139880 33440
rect 139720 33440 139880 33600
rect 139720 33600 139880 33760
rect 139720 33760 139880 33920
rect 139720 33920 139880 34080
rect 139720 34080 139880 34240
rect 139720 34240 139880 34400
rect 139720 34400 139880 34560
rect 139720 34560 139880 34720
rect 139720 34720 139880 34880
rect 139720 34880 139880 35040
rect 139720 35040 139880 35200
rect 139720 47360 139880 47520
rect 139720 47520 139880 47680
rect 139720 47680 139880 47840
rect 139720 47840 139880 48000
rect 139720 48000 139880 48160
rect 139720 48160 139880 48320
rect 139720 48320 139880 48480
rect 139720 48480 139880 48640
rect 139720 48640 139880 48800
rect 139720 48800 139880 48960
rect 139720 48960 139880 49120
rect 139720 49120 139880 49280
rect 139720 49280 139880 49440
rect 139720 49440 139880 49600
rect 139720 49600 139880 49760
rect 139720 49760 139880 49920
rect 139720 49920 139880 50080
rect 139720 50080 139880 50240
rect 139720 50240 139880 50400
rect 139720 50400 139880 50560
rect 139720 50560 139880 50720
rect 139720 50720 139880 50880
rect 139720 50880 139880 51040
rect 139720 51040 139880 51200
rect 139720 51200 139880 51360
rect 139720 51360 139880 51520
rect 139720 51520 139880 51680
rect 139720 51680 139880 51840
rect 139720 51840 139880 52000
rect 139720 52000 139880 52160
rect 139880 29440 140040 29600
rect 139880 29600 140040 29760
rect 139880 29760 140040 29920
rect 139880 29920 140040 30080
rect 139880 30080 140040 30240
rect 139880 30240 140040 30400
rect 139880 30400 140040 30560
rect 139880 30560 140040 30720
rect 139880 30720 140040 30880
rect 139880 30880 140040 31040
rect 139880 31040 140040 31200
rect 139880 31200 140040 31360
rect 139880 31360 140040 31520
rect 139880 31520 140040 31680
rect 139880 31680 140040 31840
rect 139880 31840 140040 32000
rect 139880 32000 140040 32160
rect 139880 32160 140040 32320
rect 139880 32320 140040 32480
rect 139880 32480 140040 32640
rect 139880 32640 140040 32800
rect 139880 32800 140040 32960
rect 139880 32960 140040 33120
rect 139880 33120 140040 33280
rect 139880 33280 140040 33440
rect 139880 33440 140040 33600
rect 139880 33600 140040 33760
rect 139880 33760 140040 33920
rect 139880 33920 140040 34080
rect 139880 34080 140040 34240
rect 139880 34240 140040 34400
rect 139880 34400 140040 34560
rect 139880 34560 140040 34720
rect 139880 34720 140040 34880
rect 139880 34880 140040 35040
rect 139880 35040 140040 35200
rect 139880 35200 140040 35360
rect 139880 35360 140040 35520
rect 139880 35520 140040 35680
rect 139880 47040 140040 47200
rect 139880 47200 140040 47360
rect 139880 47360 140040 47520
rect 139880 47520 140040 47680
rect 139880 47680 140040 47840
rect 139880 47840 140040 48000
rect 139880 48000 140040 48160
rect 139880 48160 140040 48320
rect 139880 48320 140040 48480
rect 139880 48480 140040 48640
rect 139880 48640 140040 48800
rect 139880 48800 140040 48960
rect 139880 48960 140040 49120
rect 139880 49120 140040 49280
rect 139880 49280 140040 49440
rect 139880 49440 140040 49600
rect 139880 49600 140040 49760
rect 139880 49760 140040 49920
rect 139880 49920 140040 50080
rect 139880 50080 140040 50240
rect 139880 50240 140040 50400
rect 139880 50400 140040 50560
rect 139880 50560 140040 50720
rect 139880 50720 140040 50880
rect 139880 50880 140040 51040
rect 139880 51040 140040 51200
rect 139880 51200 140040 51360
rect 139880 51360 140040 51520
rect 139880 51520 140040 51680
rect 139880 51680 140040 51840
rect 139880 51840 140040 52000
rect 139880 52000 140040 52160
rect 140040 29600 140200 29760
rect 140040 29760 140200 29920
rect 140040 29920 140200 30080
rect 140040 30080 140200 30240
rect 140040 30240 140200 30400
rect 140040 30400 140200 30560
rect 140040 30560 140200 30720
rect 140040 30720 140200 30880
rect 140040 30880 140200 31040
rect 140040 31040 140200 31200
rect 140040 31200 140200 31360
rect 140040 31360 140200 31520
rect 140040 31520 140200 31680
rect 140040 31680 140200 31840
rect 140040 31840 140200 32000
rect 140040 32000 140200 32160
rect 140040 32160 140200 32320
rect 140040 32320 140200 32480
rect 140040 32480 140200 32640
rect 140040 32640 140200 32800
rect 140040 32800 140200 32960
rect 140040 32960 140200 33120
rect 140040 33120 140200 33280
rect 140040 33280 140200 33440
rect 140040 33440 140200 33600
rect 140040 33600 140200 33760
rect 140040 33760 140200 33920
rect 140040 33920 140200 34080
rect 140040 34080 140200 34240
rect 140040 34240 140200 34400
rect 140040 34400 140200 34560
rect 140040 34560 140200 34720
rect 140040 34720 140200 34880
rect 140040 34880 140200 35040
rect 140040 35040 140200 35200
rect 140040 35200 140200 35360
rect 140040 35360 140200 35520
rect 140040 35520 140200 35680
rect 140040 35680 140200 35840
rect 140040 35840 140200 36000
rect 140040 36000 140200 36160
rect 140040 46560 140200 46720
rect 140040 46720 140200 46880
rect 140040 46880 140200 47040
rect 140040 47040 140200 47200
rect 140040 47200 140200 47360
rect 140040 47360 140200 47520
rect 140040 47520 140200 47680
rect 140040 47680 140200 47840
rect 140040 47840 140200 48000
rect 140040 48000 140200 48160
rect 140040 48160 140200 48320
rect 140040 48320 140200 48480
rect 140040 48480 140200 48640
rect 140040 48640 140200 48800
rect 140040 48800 140200 48960
rect 140040 48960 140200 49120
rect 140040 49120 140200 49280
rect 140040 49280 140200 49440
rect 140040 49440 140200 49600
rect 140040 49600 140200 49760
rect 140040 49760 140200 49920
rect 140040 49920 140200 50080
rect 140040 50080 140200 50240
rect 140040 50240 140200 50400
rect 140040 50400 140200 50560
rect 140040 50560 140200 50720
rect 140040 50720 140200 50880
rect 140040 50880 140200 51040
rect 140040 51040 140200 51200
rect 140040 51200 140200 51360
rect 140040 51360 140200 51520
rect 140040 51520 140200 51680
rect 140040 51680 140200 51840
rect 140040 51840 140200 52000
rect 140200 29760 140360 29920
rect 140200 29920 140360 30080
rect 140200 30080 140360 30240
rect 140200 30240 140360 30400
rect 140200 30400 140360 30560
rect 140200 30560 140360 30720
rect 140200 30720 140360 30880
rect 140200 30880 140360 31040
rect 140200 31040 140360 31200
rect 140200 31200 140360 31360
rect 140200 31360 140360 31520
rect 140200 31520 140360 31680
rect 140200 31680 140360 31840
rect 140200 31840 140360 32000
rect 140200 32000 140360 32160
rect 140200 32160 140360 32320
rect 140200 32320 140360 32480
rect 140200 32480 140360 32640
rect 140200 32640 140360 32800
rect 140200 32800 140360 32960
rect 140200 32960 140360 33120
rect 140200 33120 140360 33280
rect 140200 33280 140360 33440
rect 140200 33440 140360 33600
rect 140200 33600 140360 33760
rect 140200 33760 140360 33920
rect 140200 33920 140360 34080
rect 140200 34080 140360 34240
rect 140200 34240 140360 34400
rect 140200 34400 140360 34560
rect 140200 34560 140360 34720
rect 140200 34720 140360 34880
rect 140200 34880 140360 35040
rect 140200 35040 140360 35200
rect 140200 35200 140360 35360
rect 140200 35360 140360 35520
rect 140200 35520 140360 35680
rect 140200 35680 140360 35840
rect 140200 35840 140360 36000
rect 140200 36000 140360 36160
rect 140200 36160 140360 36320
rect 140200 36320 140360 36480
rect 140200 36480 140360 36640
rect 140200 46240 140360 46400
rect 140200 46400 140360 46560
rect 140200 46560 140360 46720
rect 140200 46720 140360 46880
rect 140200 46880 140360 47040
rect 140200 47040 140360 47200
rect 140200 47200 140360 47360
rect 140200 47360 140360 47520
rect 140200 47520 140360 47680
rect 140200 47680 140360 47840
rect 140200 47840 140360 48000
rect 140200 48000 140360 48160
rect 140200 48160 140360 48320
rect 140200 48320 140360 48480
rect 140200 48480 140360 48640
rect 140200 48640 140360 48800
rect 140200 48800 140360 48960
rect 140200 48960 140360 49120
rect 140200 49120 140360 49280
rect 140200 49280 140360 49440
rect 140200 49440 140360 49600
rect 140200 49600 140360 49760
rect 140200 49760 140360 49920
rect 140200 49920 140360 50080
rect 140200 50080 140360 50240
rect 140200 50240 140360 50400
rect 140200 50400 140360 50560
rect 140200 50560 140360 50720
rect 140200 50720 140360 50880
rect 140200 50880 140360 51040
rect 140200 51040 140360 51200
rect 140200 51200 140360 51360
rect 140200 51360 140360 51520
rect 140200 51520 140360 51680
rect 140200 51680 140360 51840
rect 140360 29920 140520 30080
rect 140360 30080 140520 30240
rect 140360 30240 140520 30400
rect 140360 30400 140520 30560
rect 140360 30560 140520 30720
rect 140360 30720 140520 30880
rect 140360 30880 140520 31040
rect 140360 31040 140520 31200
rect 140360 31200 140520 31360
rect 140360 31360 140520 31520
rect 140360 31520 140520 31680
rect 140360 31680 140520 31840
rect 140360 31840 140520 32000
rect 140360 32000 140520 32160
rect 140360 32160 140520 32320
rect 140360 32320 140520 32480
rect 140360 32480 140520 32640
rect 140360 32640 140520 32800
rect 140360 32800 140520 32960
rect 140360 32960 140520 33120
rect 140360 33120 140520 33280
rect 140360 33280 140520 33440
rect 140360 33440 140520 33600
rect 140360 33600 140520 33760
rect 140360 33760 140520 33920
rect 140360 33920 140520 34080
rect 140360 34080 140520 34240
rect 140360 34240 140520 34400
rect 140360 34400 140520 34560
rect 140360 34560 140520 34720
rect 140360 34720 140520 34880
rect 140360 34880 140520 35040
rect 140360 35040 140520 35200
rect 140360 35200 140520 35360
rect 140360 35360 140520 35520
rect 140360 35520 140520 35680
rect 140360 35680 140520 35840
rect 140360 35840 140520 36000
rect 140360 36000 140520 36160
rect 140360 36160 140520 36320
rect 140360 36320 140520 36480
rect 140360 36480 140520 36640
rect 140360 36640 140520 36800
rect 140360 36800 140520 36960
rect 140360 36960 140520 37120
rect 140360 45600 140520 45760
rect 140360 45760 140520 45920
rect 140360 45920 140520 46080
rect 140360 46080 140520 46240
rect 140360 46240 140520 46400
rect 140360 46400 140520 46560
rect 140360 46560 140520 46720
rect 140360 46720 140520 46880
rect 140360 46880 140520 47040
rect 140360 47040 140520 47200
rect 140360 47200 140520 47360
rect 140360 47360 140520 47520
rect 140360 47520 140520 47680
rect 140360 47680 140520 47840
rect 140360 47840 140520 48000
rect 140360 48000 140520 48160
rect 140360 48160 140520 48320
rect 140360 48320 140520 48480
rect 140360 48480 140520 48640
rect 140360 48640 140520 48800
rect 140360 48800 140520 48960
rect 140360 48960 140520 49120
rect 140360 49120 140520 49280
rect 140360 49280 140520 49440
rect 140360 49440 140520 49600
rect 140360 49600 140520 49760
rect 140360 49760 140520 49920
rect 140360 49920 140520 50080
rect 140360 50080 140520 50240
rect 140360 50240 140520 50400
rect 140360 50400 140520 50560
rect 140360 50560 140520 50720
rect 140360 50720 140520 50880
rect 140360 50880 140520 51040
rect 140360 51040 140520 51200
rect 140360 51200 140520 51360
rect 140360 51360 140520 51520
rect 140360 51520 140520 51680
rect 140360 51680 140520 51840
rect 140520 30240 140680 30400
rect 140520 30400 140680 30560
rect 140520 30560 140680 30720
rect 140520 30720 140680 30880
rect 140520 30880 140680 31040
rect 140520 31040 140680 31200
rect 140520 31200 140680 31360
rect 140520 31360 140680 31520
rect 140520 31520 140680 31680
rect 140520 31680 140680 31840
rect 140520 31840 140680 32000
rect 140520 32000 140680 32160
rect 140520 32160 140680 32320
rect 140520 32320 140680 32480
rect 140520 32480 140680 32640
rect 140520 32640 140680 32800
rect 140520 32800 140680 32960
rect 140520 32960 140680 33120
rect 140520 33120 140680 33280
rect 140520 33280 140680 33440
rect 140520 33440 140680 33600
rect 140520 33600 140680 33760
rect 140520 33760 140680 33920
rect 140520 33920 140680 34080
rect 140520 34080 140680 34240
rect 140520 34240 140680 34400
rect 140520 34400 140680 34560
rect 140520 34560 140680 34720
rect 140520 34720 140680 34880
rect 140520 34880 140680 35040
rect 140520 35040 140680 35200
rect 140520 35200 140680 35360
rect 140520 35360 140680 35520
rect 140520 35520 140680 35680
rect 140520 35680 140680 35840
rect 140520 35840 140680 36000
rect 140520 36000 140680 36160
rect 140520 36160 140680 36320
rect 140520 36320 140680 36480
rect 140520 36480 140680 36640
rect 140520 36640 140680 36800
rect 140520 36800 140680 36960
rect 140520 36960 140680 37120
rect 140520 37120 140680 37280
rect 140520 37280 140680 37440
rect 140520 37440 140680 37600
rect 140520 37600 140680 37760
rect 140520 44960 140680 45120
rect 140520 45120 140680 45280
rect 140520 45280 140680 45440
rect 140520 45440 140680 45600
rect 140520 45600 140680 45760
rect 140520 45760 140680 45920
rect 140520 45920 140680 46080
rect 140520 46080 140680 46240
rect 140520 46240 140680 46400
rect 140520 46400 140680 46560
rect 140520 46560 140680 46720
rect 140520 46720 140680 46880
rect 140520 46880 140680 47040
rect 140520 47040 140680 47200
rect 140520 47200 140680 47360
rect 140520 47360 140680 47520
rect 140520 47520 140680 47680
rect 140520 47680 140680 47840
rect 140520 47840 140680 48000
rect 140520 48000 140680 48160
rect 140520 48160 140680 48320
rect 140520 48320 140680 48480
rect 140520 48480 140680 48640
rect 140520 48640 140680 48800
rect 140520 48800 140680 48960
rect 140520 48960 140680 49120
rect 140520 49120 140680 49280
rect 140520 49280 140680 49440
rect 140520 49440 140680 49600
rect 140520 49600 140680 49760
rect 140520 49760 140680 49920
rect 140520 49920 140680 50080
rect 140520 50080 140680 50240
rect 140520 50240 140680 50400
rect 140520 50400 140680 50560
rect 140520 50560 140680 50720
rect 140520 50720 140680 50880
rect 140520 50880 140680 51040
rect 140520 51040 140680 51200
rect 140520 51200 140680 51360
rect 140520 51360 140680 51520
rect 140520 51520 140680 51680
rect 140680 30400 140840 30560
rect 140680 30560 140840 30720
rect 140680 30720 140840 30880
rect 140680 30880 140840 31040
rect 140680 31040 140840 31200
rect 140680 31200 140840 31360
rect 140680 31360 140840 31520
rect 140680 31520 140840 31680
rect 140680 31680 140840 31840
rect 140680 31840 140840 32000
rect 140680 32000 140840 32160
rect 140680 32160 140840 32320
rect 140680 32320 140840 32480
rect 140680 32480 140840 32640
rect 140680 32640 140840 32800
rect 140680 32800 140840 32960
rect 140680 32960 140840 33120
rect 140680 33120 140840 33280
rect 140680 33280 140840 33440
rect 140680 33440 140840 33600
rect 140680 33600 140840 33760
rect 140680 33760 140840 33920
rect 140680 33920 140840 34080
rect 140680 34080 140840 34240
rect 140680 34240 140840 34400
rect 140680 34400 140840 34560
rect 140680 34560 140840 34720
rect 140680 34720 140840 34880
rect 140680 34880 140840 35040
rect 140680 35040 140840 35200
rect 140680 35200 140840 35360
rect 140680 35360 140840 35520
rect 140680 35520 140840 35680
rect 140680 35680 140840 35840
rect 140680 35840 140840 36000
rect 140680 36000 140840 36160
rect 140680 36160 140840 36320
rect 140680 36320 140840 36480
rect 140680 36480 140840 36640
rect 140680 36640 140840 36800
rect 140680 36800 140840 36960
rect 140680 36960 140840 37120
rect 140680 37120 140840 37280
rect 140680 37280 140840 37440
rect 140680 37440 140840 37600
rect 140680 37600 140840 37760
rect 140680 37760 140840 37920
rect 140680 37920 140840 38080
rect 140680 38080 140840 38240
rect 140680 38240 140840 38400
rect 140680 38400 140840 38560
rect 140680 44160 140840 44320
rect 140680 44320 140840 44480
rect 140680 44480 140840 44640
rect 140680 44640 140840 44800
rect 140680 44800 140840 44960
rect 140680 44960 140840 45120
rect 140680 45120 140840 45280
rect 140680 45280 140840 45440
rect 140680 45440 140840 45600
rect 140680 45600 140840 45760
rect 140680 45760 140840 45920
rect 140680 45920 140840 46080
rect 140680 46080 140840 46240
rect 140680 46240 140840 46400
rect 140680 46400 140840 46560
rect 140680 46560 140840 46720
rect 140680 46720 140840 46880
rect 140680 46880 140840 47040
rect 140680 47040 140840 47200
rect 140680 47200 140840 47360
rect 140680 47360 140840 47520
rect 140680 47520 140840 47680
rect 140680 47680 140840 47840
rect 140680 47840 140840 48000
rect 140680 48000 140840 48160
rect 140680 48160 140840 48320
rect 140680 48320 140840 48480
rect 140680 48480 140840 48640
rect 140680 48640 140840 48800
rect 140680 48800 140840 48960
rect 140680 48960 140840 49120
rect 140680 49120 140840 49280
rect 140680 49280 140840 49440
rect 140680 49440 140840 49600
rect 140680 49600 140840 49760
rect 140680 49760 140840 49920
rect 140680 49920 140840 50080
rect 140680 50080 140840 50240
rect 140680 50240 140840 50400
rect 140680 50400 140840 50560
rect 140680 50560 140840 50720
rect 140680 50720 140840 50880
rect 140680 50880 140840 51040
rect 140680 51040 140840 51200
rect 140680 51200 140840 51360
rect 140680 51360 140840 51520
rect 140840 30560 141000 30720
rect 140840 30720 141000 30880
rect 140840 30880 141000 31040
rect 140840 31040 141000 31200
rect 140840 31200 141000 31360
rect 140840 31360 141000 31520
rect 140840 31520 141000 31680
rect 140840 31680 141000 31840
rect 140840 31840 141000 32000
rect 140840 32000 141000 32160
rect 140840 32160 141000 32320
rect 140840 32320 141000 32480
rect 140840 32480 141000 32640
rect 140840 32640 141000 32800
rect 140840 32800 141000 32960
rect 140840 32960 141000 33120
rect 140840 33120 141000 33280
rect 140840 33280 141000 33440
rect 140840 33440 141000 33600
rect 140840 33600 141000 33760
rect 140840 33760 141000 33920
rect 140840 33920 141000 34080
rect 140840 34080 141000 34240
rect 140840 34240 141000 34400
rect 140840 34400 141000 34560
rect 140840 34560 141000 34720
rect 140840 34720 141000 34880
rect 140840 34880 141000 35040
rect 140840 35040 141000 35200
rect 140840 35200 141000 35360
rect 140840 35360 141000 35520
rect 140840 35520 141000 35680
rect 140840 35680 141000 35840
rect 140840 35840 141000 36000
rect 140840 36000 141000 36160
rect 140840 36160 141000 36320
rect 140840 36320 141000 36480
rect 140840 36480 141000 36640
rect 140840 36640 141000 36800
rect 140840 36800 141000 36960
rect 140840 36960 141000 37120
rect 140840 37120 141000 37280
rect 140840 37280 141000 37440
rect 140840 37440 141000 37600
rect 140840 37600 141000 37760
rect 140840 37760 141000 37920
rect 140840 37920 141000 38080
rect 140840 38080 141000 38240
rect 140840 38240 141000 38400
rect 140840 38400 141000 38560
rect 140840 38560 141000 38720
rect 140840 38720 141000 38880
rect 140840 38880 141000 39040
rect 140840 39040 141000 39200
rect 140840 39200 141000 39360
rect 140840 39360 141000 39520
rect 140840 39520 141000 39680
rect 140840 42880 141000 43040
rect 140840 43040 141000 43200
rect 140840 43200 141000 43360
rect 140840 43360 141000 43520
rect 140840 43520 141000 43680
rect 140840 43680 141000 43840
rect 140840 43840 141000 44000
rect 140840 44000 141000 44160
rect 140840 44160 141000 44320
rect 140840 44320 141000 44480
rect 140840 44480 141000 44640
rect 140840 44640 141000 44800
rect 140840 44800 141000 44960
rect 140840 44960 141000 45120
rect 140840 45120 141000 45280
rect 140840 45280 141000 45440
rect 140840 45440 141000 45600
rect 140840 45600 141000 45760
rect 140840 45760 141000 45920
rect 140840 45920 141000 46080
rect 140840 46080 141000 46240
rect 140840 46240 141000 46400
rect 140840 46400 141000 46560
rect 140840 46560 141000 46720
rect 140840 46720 141000 46880
rect 140840 46880 141000 47040
rect 140840 47040 141000 47200
rect 140840 47200 141000 47360
rect 140840 47360 141000 47520
rect 140840 47520 141000 47680
rect 140840 47680 141000 47840
rect 140840 47840 141000 48000
rect 140840 48000 141000 48160
rect 140840 48160 141000 48320
rect 140840 48320 141000 48480
rect 140840 48480 141000 48640
rect 140840 48640 141000 48800
rect 140840 48800 141000 48960
rect 140840 48960 141000 49120
rect 140840 49120 141000 49280
rect 140840 49280 141000 49440
rect 140840 49440 141000 49600
rect 140840 49600 141000 49760
rect 140840 49760 141000 49920
rect 140840 49920 141000 50080
rect 140840 50080 141000 50240
rect 140840 50240 141000 50400
rect 140840 50400 141000 50560
rect 140840 50560 141000 50720
rect 140840 50720 141000 50880
rect 140840 50880 141000 51040
rect 140840 51040 141000 51200
rect 140840 51200 141000 51360
rect 141000 30720 141160 30880
rect 141000 30880 141160 31040
rect 141000 31040 141160 31200
rect 141000 31200 141160 31360
rect 141000 31360 141160 31520
rect 141000 31520 141160 31680
rect 141000 31680 141160 31840
rect 141000 31840 141160 32000
rect 141000 32000 141160 32160
rect 141000 32160 141160 32320
rect 141000 32320 141160 32480
rect 141000 32480 141160 32640
rect 141000 32640 141160 32800
rect 141000 32800 141160 32960
rect 141000 32960 141160 33120
rect 141000 33120 141160 33280
rect 141000 33280 141160 33440
rect 141000 33440 141160 33600
rect 141000 33600 141160 33760
rect 141000 33760 141160 33920
rect 141000 33920 141160 34080
rect 141000 34080 141160 34240
rect 141000 34240 141160 34400
rect 141000 34400 141160 34560
rect 141000 34560 141160 34720
rect 141000 34720 141160 34880
rect 141000 34880 141160 35040
rect 141000 35040 141160 35200
rect 141000 35200 141160 35360
rect 141000 35360 141160 35520
rect 141000 35520 141160 35680
rect 141000 35680 141160 35840
rect 141000 35840 141160 36000
rect 141000 36000 141160 36160
rect 141000 36160 141160 36320
rect 141000 36320 141160 36480
rect 141000 36480 141160 36640
rect 141000 36640 141160 36800
rect 141000 36800 141160 36960
rect 141000 36960 141160 37120
rect 141000 37120 141160 37280
rect 141000 37280 141160 37440
rect 141000 37440 141160 37600
rect 141000 37600 141160 37760
rect 141000 37760 141160 37920
rect 141000 37920 141160 38080
rect 141000 38080 141160 38240
rect 141000 38240 141160 38400
rect 141000 38400 141160 38560
rect 141000 38560 141160 38720
rect 141000 38720 141160 38880
rect 141000 38880 141160 39040
rect 141000 39040 141160 39200
rect 141000 39200 141160 39360
rect 141000 39360 141160 39520
rect 141000 39520 141160 39680
rect 141000 39680 141160 39840
rect 141000 39840 141160 40000
rect 141000 40000 141160 40160
rect 141000 40160 141160 40320
rect 141000 40320 141160 40480
rect 141000 40480 141160 40640
rect 141000 40640 141160 40800
rect 141000 40800 141160 40960
rect 141000 40960 141160 41120
rect 141000 41120 141160 41280
rect 141000 41280 141160 41440
rect 141000 41440 141160 41600
rect 141000 41600 141160 41760
rect 141000 41760 141160 41920
rect 141000 41920 141160 42080
rect 141000 42080 141160 42240
rect 141000 42240 141160 42400
rect 141000 42400 141160 42560
rect 141000 42560 141160 42720
rect 141000 42720 141160 42880
rect 141000 42880 141160 43040
rect 141000 43040 141160 43200
rect 141000 43200 141160 43360
rect 141000 43360 141160 43520
rect 141000 43520 141160 43680
rect 141000 43680 141160 43840
rect 141000 43840 141160 44000
rect 141000 44000 141160 44160
rect 141000 44160 141160 44320
rect 141000 44320 141160 44480
rect 141000 44480 141160 44640
rect 141000 44640 141160 44800
rect 141000 44800 141160 44960
rect 141000 44960 141160 45120
rect 141000 45120 141160 45280
rect 141000 45280 141160 45440
rect 141000 45440 141160 45600
rect 141000 45600 141160 45760
rect 141000 45760 141160 45920
rect 141000 45920 141160 46080
rect 141000 46080 141160 46240
rect 141000 46240 141160 46400
rect 141000 46400 141160 46560
rect 141000 46560 141160 46720
rect 141000 46720 141160 46880
rect 141000 46880 141160 47040
rect 141000 47040 141160 47200
rect 141000 47200 141160 47360
rect 141000 47360 141160 47520
rect 141000 47520 141160 47680
rect 141000 47680 141160 47840
rect 141000 47840 141160 48000
rect 141000 48000 141160 48160
rect 141000 48160 141160 48320
rect 141000 48320 141160 48480
rect 141000 48480 141160 48640
rect 141000 48640 141160 48800
rect 141000 48800 141160 48960
rect 141000 48960 141160 49120
rect 141000 49120 141160 49280
rect 141000 49280 141160 49440
rect 141000 49440 141160 49600
rect 141000 49600 141160 49760
rect 141000 49760 141160 49920
rect 141000 49920 141160 50080
rect 141000 50080 141160 50240
rect 141000 50240 141160 50400
rect 141000 50400 141160 50560
rect 141000 50560 141160 50720
rect 141000 50720 141160 50880
rect 141000 50880 141160 51040
rect 141000 51040 141160 51200
rect 141160 31040 141320 31200
rect 141160 31200 141320 31360
rect 141160 31360 141320 31520
rect 141160 31520 141320 31680
rect 141160 31680 141320 31840
rect 141160 31840 141320 32000
rect 141160 32000 141320 32160
rect 141160 32160 141320 32320
rect 141160 32320 141320 32480
rect 141160 32480 141320 32640
rect 141160 32640 141320 32800
rect 141160 32800 141320 32960
rect 141160 32960 141320 33120
rect 141160 33120 141320 33280
rect 141160 33280 141320 33440
rect 141160 33440 141320 33600
rect 141160 33600 141320 33760
rect 141160 33760 141320 33920
rect 141160 33920 141320 34080
rect 141160 34080 141320 34240
rect 141160 34240 141320 34400
rect 141160 34400 141320 34560
rect 141160 34560 141320 34720
rect 141160 34720 141320 34880
rect 141160 34880 141320 35040
rect 141160 35040 141320 35200
rect 141160 35200 141320 35360
rect 141160 35360 141320 35520
rect 141160 35520 141320 35680
rect 141160 35680 141320 35840
rect 141160 35840 141320 36000
rect 141160 36000 141320 36160
rect 141160 36160 141320 36320
rect 141160 36320 141320 36480
rect 141160 36480 141320 36640
rect 141160 36640 141320 36800
rect 141160 36800 141320 36960
rect 141160 36960 141320 37120
rect 141160 37120 141320 37280
rect 141160 37280 141320 37440
rect 141160 37440 141320 37600
rect 141160 37600 141320 37760
rect 141160 37760 141320 37920
rect 141160 37920 141320 38080
rect 141160 38080 141320 38240
rect 141160 38240 141320 38400
rect 141160 38400 141320 38560
rect 141160 38560 141320 38720
rect 141160 38720 141320 38880
rect 141160 38880 141320 39040
rect 141160 39040 141320 39200
rect 141160 39200 141320 39360
rect 141160 39360 141320 39520
rect 141160 39520 141320 39680
rect 141160 39680 141320 39840
rect 141160 39840 141320 40000
rect 141160 40000 141320 40160
rect 141160 40160 141320 40320
rect 141160 40320 141320 40480
rect 141160 40480 141320 40640
rect 141160 40640 141320 40800
rect 141160 40800 141320 40960
rect 141160 40960 141320 41120
rect 141160 41120 141320 41280
rect 141160 41280 141320 41440
rect 141160 41440 141320 41600
rect 141160 41600 141320 41760
rect 141160 41760 141320 41920
rect 141160 41920 141320 42080
rect 141160 42080 141320 42240
rect 141160 42240 141320 42400
rect 141160 42400 141320 42560
rect 141160 42560 141320 42720
rect 141160 42720 141320 42880
rect 141160 42880 141320 43040
rect 141160 43040 141320 43200
rect 141160 43200 141320 43360
rect 141160 43360 141320 43520
rect 141160 43520 141320 43680
rect 141160 43680 141320 43840
rect 141160 43840 141320 44000
rect 141160 44000 141320 44160
rect 141160 44160 141320 44320
rect 141160 44320 141320 44480
rect 141160 44480 141320 44640
rect 141160 44640 141320 44800
rect 141160 44800 141320 44960
rect 141160 44960 141320 45120
rect 141160 45120 141320 45280
rect 141160 45280 141320 45440
rect 141160 45440 141320 45600
rect 141160 45600 141320 45760
rect 141160 45760 141320 45920
rect 141160 45920 141320 46080
rect 141160 46080 141320 46240
rect 141160 46240 141320 46400
rect 141160 46400 141320 46560
rect 141160 46560 141320 46720
rect 141160 46720 141320 46880
rect 141160 46880 141320 47040
rect 141160 47040 141320 47200
rect 141160 47200 141320 47360
rect 141160 47360 141320 47520
rect 141160 47520 141320 47680
rect 141160 47680 141320 47840
rect 141160 47840 141320 48000
rect 141160 48000 141320 48160
rect 141160 48160 141320 48320
rect 141160 48320 141320 48480
rect 141160 48480 141320 48640
rect 141160 48640 141320 48800
rect 141160 48800 141320 48960
rect 141160 48960 141320 49120
rect 141160 49120 141320 49280
rect 141160 49280 141320 49440
rect 141160 49440 141320 49600
rect 141160 49600 141320 49760
rect 141160 49760 141320 49920
rect 141160 49920 141320 50080
rect 141160 50080 141320 50240
rect 141160 50240 141320 50400
rect 141160 50400 141320 50560
rect 141160 50560 141320 50720
rect 141160 50720 141320 50880
rect 141160 50880 141320 51040
rect 141320 31200 141480 31360
rect 141320 31360 141480 31520
rect 141320 31520 141480 31680
rect 141320 31680 141480 31840
rect 141320 31840 141480 32000
rect 141320 32000 141480 32160
rect 141320 32160 141480 32320
rect 141320 32320 141480 32480
rect 141320 32480 141480 32640
rect 141320 32640 141480 32800
rect 141320 32800 141480 32960
rect 141320 32960 141480 33120
rect 141320 33120 141480 33280
rect 141320 33280 141480 33440
rect 141320 33440 141480 33600
rect 141320 33600 141480 33760
rect 141320 33760 141480 33920
rect 141320 33920 141480 34080
rect 141320 34080 141480 34240
rect 141320 34240 141480 34400
rect 141320 34400 141480 34560
rect 141320 34560 141480 34720
rect 141320 34720 141480 34880
rect 141320 34880 141480 35040
rect 141320 35040 141480 35200
rect 141320 35200 141480 35360
rect 141320 35360 141480 35520
rect 141320 35520 141480 35680
rect 141320 35680 141480 35840
rect 141320 35840 141480 36000
rect 141320 36000 141480 36160
rect 141320 36160 141480 36320
rect 141320 36320 141480 36480
rect 141320 36480 141480 36640
rect 141320 36640 141480 36800
rect 141320 36800 141480 36960
rect 141320 36960 141480 37120
rect 141320 37120 141480 37280
rect 141320 37280 141480 37440
rect 141320 37440 141480 37600
rect 141320 37600 141480 37760
rect 141320 37760 141480 37920
rect 141320 37920 141480 38080
rect 141320 38080 141480 38240
rect 141320 38240 141480 38400
rect 141320 38400 141480 38560
rect 141320 38560 141480 38720
rect 141320 38720 141480 38880
rect 141320 38880 141480 39040
rect 141320 39040 141480 39200
rect 141320 39200 141480 39360
rect 141320 39360 141480 39520
rect 141320 39520 141480 39680
rect 141320 39680 141480 39840
rect 141320 39840 141480 40000
rect 141320 40000 141480 40160
rect 141320 40160 141480 40320
rect 141320 40320 141480 40480
rect 141320 40480 141480 40640
rect 141320 40640 141480 40800
rect 141320 40800 141480 40960
rect 141320 40960 141480 41120
rect 141320 41120 141480 41280
rect 141320 41280 141480 41440
rect 141320 41440 141480 41600
rect 141320 41600 141480 41760
rect 141320 41760 141480 41920
rect 141320 41920 141480 42080
rect 141320 42080 141480 42240
rect 141320 42240 141480 42400
rect 141320 42400 141480 42560
rect 141320 42560 141480 42720
rect 141320 42720 141480 42880
rect 141320 42880 141480 43040
rect 141320 43040 141480 43200
rect 141320 43200 141480 43360
rect 141320 43360 141480 43520
rect 141320 43520 141480 43680
rect 141320 43680 141480 43840
rect 141320 43840 141480 44000
rect 141320 44000 141480 44160
rect 141320 44160 141480 44320
rect 141320 44320 141480 44480
rect 141320 44480 141480 44640
rect 141320 44640 141480 44800
rect 141320 44800 141480 44960
rect 141320 44960 141480 45120
rect 141320 45120 141480 45280
rect 141320 45280 141480 45440
rect 141320 45440 141480 45600
rect 141320 45600 141480 45760
rect 141320 45760 141480 45920
rect 141320 45920 141480 46080
rect 141320 46080 141480 46240
rect 141320 46240 141480 46400
rect 141320 46400 141480 46560
rect 141320 46560 141480 46720
rect 141320 46720 141480 46880
rect 141320 46880 141480 47040
rect 141320 47040 141480 47200
rect 141320 47200 141480 47360
rect 141320 47360 141480 47520
rect 141320 47520 141480 47680
rect 141320 47680 141480 47840
rect 141320 47840 141480 48000
rect 141320 48000 141480 48160
rect 141320 48160 141480 48320
rect 141320 48320 141480 48480
rect 141320 48480 141480 48640
rect 141320 48640 141480 48800
rect 141320 48800 141480 48960
rect 141320 48960 141480 49120
rect 141320 49120 141480 49280
rect 141320 49280 141480 49440
rect 141320 49440 141480 49600
rect 141320 49600 141480 49760
rect 141320 49760 141480 49920
rect 141320 49920 141480 50080
rect 141320 50080 141480 50240
rect 141320 50240 141480 50400
rect 141320 50400 141480 50560
rect 141320 50560 141480 50720
rect 141320 50720 141480 50880
rect 141480 31520 141640 31680
rect 141480 31680 141640 31840
rect 141480 31840 141640 32000
rect 141480 32000 141640 32160
rect 141480 32160 141640 32320
rect 141480 32320 141640 32480
rect 141480 32480 141640 32640
rect 141480 32640 141640 32800
rect 141480 32800 141640 32960
rect 141480 32960 141640 33120
rect 141480 33120 141640 33280
rect 141480 33280 141640 33440
rect 141480 33440 141640 33600
rect 141480 33600 141640 33760
rect 141480 33760 141640 33920
rect 141480 33920 141640 34080
rect 141480 34080 141640 34240
rect 141480 34240 141640 34400
rect 141480 34400 141640 34560
rect 141480 34560 141640 34720
rect 141480 34720 141640 34880
rect 141480 34880 141640 35040
rect 141480 35040 141640 35200
rect 141480 35200 141640 35360
rect 141480 35360 141640 35520
rect 141480 35520 141640 35680
rect 141480 35680 141640 35840
rect 141480 35840 141640 36000
rect 141480 36000 141640 36160
rect 141480 36160 141640 36320
rect 141480 36320 141640 36480
rect 141480 36480 141640 36640
rect 141480 36640 141640 36800
rect 141480 36800 141640 36960
rect 141480 36960 141640 37120
rect 141480 37120 141640 37280
rect 141480 37280 141640 37440
rect 141480 37440 141640 37600
rect 141480 37600 141640 37760
rect 141480 37760 141640 37920
rect 141480 37920 141640 38080
rect 141480 38080 141640 38240
rect 141480 38240 141640 38400
rect 141480 38400 141640 38560
rect 141480 38560 141640 38720
rect 141480 38720 141640 38880
rect 141480 38880 141640 39040
rect 141480 39040 141640 39200
rect 141480 39200 141640 39360
rect 141480 39360 141640 39520
rect 141480 39520 141640 39680
rect 141480 39680 141640 39840
rect 141480 39840 141640 40000
rect 141480 40000 141640 40160
rect 141480 40160 141640 40320
rect 141480 40320 141640 40480
rect 141480 40480 141640 40640
rect 141480 40640 141640 40800
rect 141480 40800 141640 40960
rect 141480 40960 141640 41120
rect 141480 41120 141640 41280
rect 141480 41280 141640 41440
rect 141480 41440 141640 41600
rect 141480 41600 141640 41760
rect 141480 41760 141640 41920
rect 141480 41920 141640 42080
rect 141480 42080 141640 42240
rect 141480 42240 141640 42400
rect 141480 42400 141640 42560
rect 141480 42560 141640 42720
rect 141480 42720 141640 42880
rect 141480 42880 141640 43040
rect 141480 43040 141640 43200
rect 141480 43200 141640 43360
rect 141480 43360 141640 43520
rect 141480 43520 141640 43680
rect 141480 43680 141640 43840
rect 141480 43840 141640 44000
rect 141480 44000 141640 44160
rect 141480 44160 141640 44320
rect 141480 44320 141640 44480
rect 141480 44480 141640 44640
rect 141480 44640 141640 44800
rect 141480 44800 141640 44960
rect 141480 44960 141640 45120
rect 141480 45120 141640 45280
rect 141480 45280 141640 45440
rect 141480 45440 141640 45600
rect 141480 45600 141640 45760
rect 141480 45760 141640 45920
rect 141480 45920 141640 46080
rect 141480 46080 141640 46240
rect 141480 46240 141640 46400
rect 141480 46400 141640 46560
rect 141480 46560 141640 46720
rect 141480 46720 141640 46880
rect 141480 46880 141640 47040
rect 141480 47040 141640 47200
rect 141480 47200 141640 47360
rect 141480 47360 141640 47520
rect 141480 47520 141640 47680
rect 141480 47680 141640 47840
rect 141480 47840 141640 48000
rect 141480 48000 141640 48160
rect 141480 48160 141640 48320
rect 141480 48320 141640 48480
rect 141480 48480 141640 48640
rect 141480 48640 141640 48800
rect 141480 48800 141640 48960
rect 141480 48960 141640 49120
rect 141480 49120 141640 49280
rect 141480 49280 141640 49440
rect 141480 49440 141640 49600
rect 141480 49600 141640 49760
rect 141480 49760 141640 49920
rect 141480 49920 141640 50080
rect 141480 50080 141640 50240
rect 141480 50240 141640 50400
rect 141480 50400 141640 50560
rect 141480 50560 141640 50720
rect 141640 31840 141800 32000
rect 141640 32000 141800 32160
rect 141640 32160 141800 32320
rect 141640 32320 141800 32480
rect 141640 32480 141800 32640
rect 141640 32640 141800 32800
rect 141640 32800 141800 32960
rect 141640 32960 141800 33120
rect 141640 33120 141800 33280
rect 141640 33280 141800 33440
rect 141640 33440 141800 33600
rect 141640 33600 141800 33760
rect 141640 33760 141800 33920
rect 141640 33920 141800 34080
rect 141640 34080 141800 34240
rect 141640 34240 141800 34400
rect 141640 34400 141800 34560
rect 141640 34560 141800 34720
rect 141640 34720 141800 34880
rect 141640 34880 141800 35040
rect 141640 35040 141800 35200
rect 141640 35200 141800 35360
rect 141640 35360 141800 35520
rect 141640 35520 141800 35680
rect 141640 35680 141800 35840
rect 141640 35840 141800 36000
rect 141640 36000 141800 36160
rect 141640 36160 141800 36320
rect 141640 36320 141800 36480
rect 141640 36480 141800 36640
rect 141640 36640 141800 36800
rect 141640 36800 141800 36960
rect 141640 36960 141800 37120
rect 141640 37120 141800 37280
rect 141640 37280 141800 37440
rect 141640 37440 141800 37600
rect 141640 37600 141800 37760
rect 141640 37760 141800 37920
rect 141640 37920 141800 38080
rect 141640 38080 141800 38240
rect 141640 38240 141800 38400
rect 141640 38400 141800 38560
rect 141640 38560 141800 38720
rect 141640 38720 141800 38880
rect 141640 38880 141800 39040
rect 141640 39040 141800 39200
rect 141640 39200 141800 39360
rect 141640 39360 141800 39520
rect 141640 39520 141800 39680
rect 141640 39680 141800 39840
rect 141640 39840 141800 40000
rect 141640 40000 141800 40160
rect 141640 40160 141800 40320
rect 141640 40320 141800 40480
rect 141640 40480 141800 40640
rect 141640 40640 141800 40800
rect 141640 40800 141800 40960
rect 141640 40960 141800 41120
rect 141640 41120 141800 41280
rect 141640 41280 141800 41440
rect 141640 41440 141800 41600
rect 141640 41600 141800 41760
rect 141640 41760 141800 41920
rect 141640 41920 141800 42080
rect 141640 42080 141800 42240
rect 141640 42240 141800 42400
rect 141640 42400 141800 42560
rect 141640 42560 141800 42720
rect 141640 42720 141800 42880
rect 141640 42880 141800 43040
rect 141640 43040 141800 43200
rect 141640 43200 141800 43360
rect 141640 43360 141800 43520
rect 141640 43520 141800 43680
rect 141640 43680 141800 43840
rect 141640 43840 141800 44000
rect 141640 44000 141800 44160
rect 141640 44160 141800 44320
rect 141640 44320 141800 44480
rect 141640 44480 141800 44640
rect 141640 44640 141800 44800
rect 141640 44800 141800 44960
rect 141640 44960 141800 45120
rect 141640 45120 141800 45280
rect 141640 45280 141800 45440
rect 141640 45440 141800 45600
rect 141640 45600 141800 45760
rect 141640 45760 141800 45920
rect 141640 45920 141800 46080
rect 141640 46080 141800 46240
rect 141640 46240 141800 46400
rect 141640 46400 141800 46560
rect 141640 46560 141800 46720
rect 141640 46720 141800 46880
rect 141640 46880 141800 47040
rect 141640 47040 141800 47200
rect 141640 47200 141800 47360
rect 141640 47360 141800 47520
rect 141640 47520 141800 47680
rect 141640 47680 141800 47840
rect 141640 47840 141800 48000
rect 141640 48000 141800 48160
rect 141640 48160 141800 48320
rect 141640 48320 141800 48480
rect 141640 48480 141800 48640
rect 141640 48640 141800 48800
rect 141640 48800 141800 48960
rect 141640 48960 141800 49120
rect 141640 49120 141800 49280
rect 141640 49280 141800 49440
rect 141640 49440 141800 49600
rect 141640 49600 141800 49760
rect 141640 49760 141800 49920
rect 141640 49920 141800 50080
rect 141640 50080 141800 50240
rect 141640 50240 141800 50400
rect 141640 50400 141800 50560
rect 141800 32000 141960 32160
rect 141800 32160 141960 32320
rect 141800 32320 141960 32480
rect 141800 32480 141960 32640
rect 141800 32640 141960 32800
rect 141800 32800 141960 32960
rect 141800 32960 141960 33120
rect 141800 33120 141960 33280
rect 141800 33280 141960 33440
rect 141800 33440 141960 33600
rect 141800 33600 141960 33760
rect 141800 33760 141960 33920
rect 141800 33920 141960 34080
rect 141800 34080 141960 34240
rect 141800 34240 141960 34400
rect 141800 34400 141960 34560
rect 141800 34560 141960 34720
rect 141800 34720 141960 34880
rect 141800 34880 141960 35040
rect 141800 35040 141960 35200
rect 141800 35200 141960 35360
rect 141800 35360 141960 35520
rect 141800 35520 141960 35680
rect 141800 35680 141960 35840
rect 141800 35840 141960 36000
rect 141800 36000 141960 36160
rect 141800 36160 141960 36320
rect 141800 36320 141960 36480
rect 141800 36480 141960 36640
rect 141800 36640 141960 36800
rect 141800 36800 141960 36960
rect 141800 36960 141960 37120
rect 141800 37120 141960 37280
rect 141800 37280 141960 37440
rect 141800 37440 141960 37600
rect 141800 37600 141960 37760
rect 141800 37760 141960 37920
rect 141800 37920 141960 38080
rect 141800 38080 141960 38240
rect 141800 38240 141960 38400
rect 141800 38400 141960 38560
rect 141800 38560 141960 38720
rect 141800 38720 141960 38880
rect 141800 38880 141960 39040
rect 141800 39040 141960 39200
rect 141800 39200 141960 39360
rect 141800 39360 141960 39520
rect 141800 39520 141960 39680
rect 141800 39680 141960 39840
rect 141800 39840 141960 40000
rect 141800 40000 141960 40160
rect 141800 40160 141960 40320
rect 141800 40320 141960 40480
rect 141800 40480 141960 40640
rect 141800 40640 141960 40800
rect 141800 40800 141960 40960
rect 141800 40960 141960 41120
rect 141800 41120 141960 41280
rect 141800 41280 141960 41440
rect 141800 41440 141960 41600
rect 141800 41600 141960 41760
rect 141800 41760 141960 41920
rect 141800 41920 141960 42080
rect 141800 42080 141960 42240
rect 141800 42240 141960 42400
rect 141800 42400 141960 42560
rect 141800 42560 141960 42720
rect 141800 42720 141960 42880
rect 141800 42880 141960 43040
rect 141800 43040 141960 43200
rect 141800 43200 141960 43360
rect 141800 43360 141960 43520
rect 141800 43520 141960 43680
rect 141800 43680 141960 43840
rect 141800 43840 141960 44000
rect 141800 44000 141960 44160
rect 141800 44160 141960 44320
rect 141800 44320 141960 44480
rect 141800 44480 141960 44640
rect 141800 44640 141960 44800
rect 141800 44800 141960 44960
rect 141800 44960 141960 45120
rect 141800 45120 141960 45280
rect 141800 45280 141960 45440
rect 141800 45440 141960 45600
rect 141800 45600 141960 45760
rect 141800 45760 141960 45920
rect 141800 45920 141960 46080
rect 141800 46080 141960 46240
rect 141800 46240 141960 46400
rect 141800 46400 141960 46560
rect 141800 46560 141960 46720
rect 141800 46720 141960 46880
rect 141800 46880 141960 47040
rect 141800 47040 141960 47200
rect 141800 47200 141960 47360
rect 141800 47360 141960 47520
rect 141800 47520 141960 47680
rect 141800 47680 141960 47840
rect 141800 47840 141960 48000
rect 141800 48000 141960 48160
rect 141800 48160 141960 48320
rect 141800 48320 141960 48480
rect 141800 48480 141960 48640
rect 141800 48640 141960 48800
rect 141800 48800 141960 48960
rect 141800 48960 141960 49120
rect 141800 49120 141960 49280
rect 141800 49280 141960 49440
rect 141800 49440 141960 49600
rect 141800 49600 141960 49760
rect 141800 49760 141960 49920
rect 141800 49920 141960 50080
rect 141800 50080 141960 50240
rect 141960 32320 142120 32480
rect 141960 32480 142120 32640
rect 141960 32640 142120 32800
rect 141960 32800 142120 32960
rect 141960 32960 142120 33120
rect 141960 33120 142120 33280
rect 141960 33280 142120 33440
rect 141960 33440 142120 33600
rect 141960 33600 142120 33760
rect 141960 33760 142120 33920
rect 141960 33920 142120 34080
rect 141960 34080 142120 34240
rect 141960 34240 142120 34400
rect 141960 34400 142120 34560
rect 141960 34560 142120 34720
rect 141960 34720 142120 34880
rect 141960 34880 142120 35040
rect 141960 35040 142120 35200
rect 141960 35200 142120 35360
rect 141960 35360 142120 35520
rect 141960 35520 142120 35680
rect 141960 35680 142120 35840
rect 141960 35840 142120 36000
rect 141960 36000 142120 36160
rect 141960 36160 142120 36320
rect 141960 36320 142120 36480
rect 141960 36480 142120 36640
rect 141960 36640 142120 36800
rect 141960 36800 142120 36960
rect 141960 36960 142120 37120
rect 141960 37120 142120 37280
rect 141960 37280 142120 37440
rect 141960 37440 142120 37600
rect 141960 37600 142120 37760
rect 141960 37760 142120 37920
rect 141960 37920 142120 38080
rect 141960 38080 142120 38240
rect 141960 38240 142120 38400
rect 141960 38400 142120 38560
rect 141960 38560 142120 38720
rect 141960 38720 142120 38880
rect 141960 38880 142120 39040
rect 141960 39040 142120 39200
rect 141960 39200 142120 39360
rect 141960 39360 142120 39520
rect 141960 39520 142120 39680
rect 141960 39680 142120 39840
rect 141960 39840 142120 40000
rect 141960 40000 142120 40160
rect 141960 40160 142120 40320
rect 141960 40320 142120 40480
rect 141960 40480 142120 40640
rect 141960 40640 142120 40800
rect 141960 40800 142120 40960
rect 141960 40960 142120 41120
rect 141960 41120 142120 41280
rect 141960 41280 142120 41440
rect 141960 41440 142120 41600
rect 141960 41600 142120 41760
rect 141960 41760 142120 41920
rect 141960 41920 142120 42080
rect 141960 42080 142120 42240
rect 141960 42240 142120 42400
rect 141960 42400 142120 42560
rect 141960 42560 142120 42720
rect 141960 42720 142120 42880
rect 141960 42880 142120 43040
rect 141960 43040 142120 43200
rect 141960 43200 142120 43360
rect 141960 43360 142120 43520
rect 141960 43520 142120 43680
rect 141960 43680 142120 43840
rect 141960 43840 142120 44000
rect 141960 44000 142120 44160
rect 141960 44160 142120 44320
rect 141960 44320 142120 44480
rect 141960 44480 142120 44640
rect 141960 44640 142120 44800
rect 141960 44800 142120 44960
rect 141960 44960 142120 45120
rect 141960 45120 142120 45280
rect 141960 45280 142120 45440
rect 141960 45440 142120 45600
rect 141960 45600 142120 45760
rect 141960 45760 142120 45920
rect 141960 45920 142120 46080
rect 141960 46080 142120 46240
rect 141960 46240 142120 46400
rect 141960 46400 142120 46560
rect 141960 46560 142120 46720
rect 141960 46720 142120 46880
rect 141960 46880 142120 47040
rect 141960 47040 142120 47200
rect 141960 47200 142120 47360
rect 141960 47360 142120 47520
rect 141960 47520 142120 47680
rect 141960 47680 142120 47840
rect 141960 47840 142120 48000
rect 141960 48000 142120 48160
rect 141960 48160 142120 48320
rect 141960 48320 142120 48480
rect 141960 48480 142120 48640
rect 141960 48640 142120 48800
rect 141960 48800 142120 48960
rect 141960 48960 142120 49120
rect 141960 49120 142120 49280
rect 141960 49280 142120 49440
rect 141960 49440 142120 49600
rect 141960 49600 142120 49760
rect 141960 49760 142120 49920
rect 141960 49920 142120 50080
rect 142120 32640 142280 32800
rect 142120 32800 142280 32960
rect 142120 32960 142280 33120
rect 142120 33120 142280 33280
rect 142120 33280 142280 33440
rect 142120 33440 142280 33600
rect 142120 33600 142280 33760
rect 142120 33760 142280 33920
rect 142120 33920 142280 34080
rect 142120 34080 142280 34240
rect 142120 34240 142280 34400
rect 142120 34400 142280 34560
rect 142120 34560 142280 34720
rect 142120 34720 142280 34880
rect 142120 34880 142280 35040
rect 142120 35040 142280 35200
rect 142120 35200 142280 35360
rect 142120 35360 142280 35520
rect 142120 35520 142280 35680
rect 142120 35680 142280 35840
rect 142120 35840 142280 36000
rect 142120 36000 142280 36160
rect 142120 36160 142280 36320
rect 142120 36320 142280 36480
rect 142120 36480 142280 36640
rect 142120 36640 142280 36800
rect 142120 36800 142280 36960
rect 142120 36960 142280 37120
rect 142120 37120 142280 37280
rect 142120 37280 142280 37440
rect 142120 37440 142280 37600
rect 142120 37600 142280 37760
rect 142120 37760 142280 37920
rect 142120 37920 142280 38080
rect 142120 38080 142280 38240
rect 142120 38240 142280 38400
rect 142120 38400 142280 38560
rect 142120 38560 142280 38720
rect 142120 38720 142280 38880
rect 142120 38880 142280 39040
rect 142120 39040 142280 39200
rect 142120 39200 142280 39360
rect 142120 39360 142280 39520
rect 142120 39520 142280 39680
rect 142120 39680 142280 39840
rect 142120 39840 142280 40000
rect 142120 40000 142280 40160
rect 142120 40160 142280 40320
rect 142120 40320 142280 40480
rect 142120 40480 142280 40640
rect 142120 40640 142280 40800
rect 142120 40800 142280 40960
rect 142120 40960 142280 41120
rect 142120 41120 142280 41280
rect 142120 41280 142280 41440
rect 142120 41440 142280 41600
rect 142120 41600 142280 41760
rect 142120 41760 142280 41920
rect 142120 41920 142280 42080
rect 142120 42080 142280 42240
rect 142120 42240 142280 42400
rect 142120 42400 142280 42560
rect 142120 42560 142280 42720
rect 142120 42720 142280 42880
rect 142120 42880 142280 43040
rect 142120 43040 142280 43200
rect 142120 43200 142280 43360
rect 142120 43360 142280 43520
rect 142120 43520 142280 43680
rect 142120 43680 142280 43840
rect 142120 43840 142280 44000
rect 142120 44000 142280 44160
rect 142120 44160 142280 44320
rect 142120 44320 142280 44480
rect 142120 44480 142280 44640
rect 142120 44640 142280 44800
rect 142120 44800 142280 44960
rect 142120 44960 142280 45120
rect 142120 45120 142280 45280
rect 142120 45280 142280 45440
rect 142120 45440 142280 45600
rect 142120 45600 142280 45760
rect 142120 45760 142280 45920
rect 142120 45920 142280 46080
rect 142120 46080 142280 46240
rect 142120 46240 142280 46400
rect 142120 46400 142280 46560
rect 142120 46560 142280 46720
rect 142120 46720 142280 46880
rect 142120 46880 142280 47040
rect 142120 47040 142280 47200
rect 142120 47200 142280 47360
rect 142120 47360 142280 47520
rect 142120 47520 142280 47680
rect 142120 47680 142280 47840
rect 142120 47840 142280 48000
rect 142120 48000 142280 48160
rect 142120 48160 142280 48320
rect 142120 48320 142280 48480
rect 142120 48480 142280 48640
rect 142120 48640 142280 48800
rect 142120 48800 142280 48960
rect 142120 48960 142280 49120
rect 142120 49120 142280 49280
rect 142120 49280 142280 49440
rect 142120 49440 142280 49600
rect 142120 49600 142280 49760
rect 142280 32960 142440 33120
rect 142280 33120 142440 33280
rect 142280 33280 142440 33440
rect 142280 33440 142440 33600
rect 142280 33600 142440 33760
rect 142280 33760 142440 33920
rect 142280 33920 142440 34080
rect 142280 34080 142440 34240
rect 142280 34240 142440 34400
rect 142280 34400 142440 34560
rect 142280 34560 142440 34720
rect 142280 34720 142440 34880
rect 142280 34880 142440 35040
rect 142280 35040 142440 35200
rect 142280 35200 142440 35360
rect 142280 35360 142440 35520
rect 142280 35520 142440 35680
rect 142280 35680 142440 35840
rect 142280 35840 142440 36000
rect 142280 36000 142440 36160
rect 142280 36160 142440 36320
rect 142280 36320 142440 36480
rect 142280 36480 142440 36640
rect 142280 36640 142440 36800
rect 142280 36800 142440 36960
rect 142280 36960 142440 37120
rect 142280 37120 142440 37280
rect 142280 37280 142440 37440
rect 142280 37440 142440 37600
rect 142280 37600 142440 37760
rect 142280 37760 142440 37920
rect 142280 37920 142440 38080
rect 142280 38080 142440 38240
rect 142280 38240 142440 38400
rect 142280 38400 142440 38560
rect 142280 38560 142440 38720
rect 142280 38720 142440 38880
rect 142280 38880 142440 39040
rect 142280 39040 142440 39200
rect 142280 39200 142440 39360
rect 142280 39360 142440 39520
rect 142280 39520 142440 39680
rect 142280 39680 142440 39840
rect 142280 39840 142440 40000
rect 142280 40000 142440 40160
rect 142280 40160 142440 40320
rect 142280 40320 142440 40480
rect 142280 40480 142440 40640
rect 142280 40640 142440 40800
rect 142280 40800 142440 40960
rect 142280 40960 142440 41120
rect 142280 41120 142440 41280
rect 142280 41280 142440 41440
rect 142280 41440 142440 41600
rect 142280 41600 142440 41760
rect 142280 41760 142440 41920
rect 142280 41920 142440 42080
rect 142280 42080 142440 42240
rect 142280 42240 142440 42400
rect 142280 42400 142440 42560
rect 142280 42560 142440 42720
rect 142280 42720 142440 42880
rect 142280 42880 142440 43040
rect 142280 43040 142440 43200
rect 142280 43200 142440 43360
rect 142280 43360 142440 43520
rect 142280 43520 142440 43680
rect 142280 43680 142440 43840
rect 142280 43840 142440 44000
rect 142280 44000 142440 44160
rect 142280 44160 142440 44320
rect 142280 44320 142440 44480
rect 142280 44480 142440 44640
rect 142280 44640 142440 44800
rect 142280 44800 142440 44960
rect 142280 44960 142440 45120
rect 142280 45120 142440 45280
rect 142280 45280 142440 45440
rect 142280 45440 142440 45600
rect 142280 45600 142440 45760
rect 142280 45760 142440 45920
rect 142280 45920 142440 46080
rect 142280 46080 142440 46240
rect 142280 46240 142440 46400
rect 142280 46400 142440 46560
rect 142280 46560 142440 46720
rect 142280 46720 142440 46880
rect 142280 46880 142440 47040
rect 142280 47040 142440 47200
rect 142280 47200 142440 47360
rect 142280 47360 142440 47520
rect 142280 47520 142440 47680
rect 142280 47680 142440 47840
rect 142280 47840 142440 48000
rect 142280 48000 142440 48160
rect 142280 48160 142440 48320
rect 142280 48320 142440 48480
rect 142280 48480 142440 48640
rect 142280 48640 142440 48800
rect 142280 48800 142440 48960
rect 142280 48960 142440 49120
rect 142280 49120 142440 49280
rect 142280 49280 142440 49440
rect 142280 49440 142440 49600
rect 142440 33280 142600 33440
rect 142440 33440 142600 33600
rect 142440 33600 142600 33760
rect 142440 33760 142600 33920
rect 142440 33920 142600 34080
rect 142440 34080 142600 34240
rect 142440 34240 142600 34400
rect 142440 34400 142600 34560
rect 142440 34560 142600 34720
rect 142440 34720 142600 34880
rect 142440 34880 142600 35040
rect 142440 35040 142600 35200
rect 142440 35200 142600 35360
rect 142440 35360 142600 35520
rect 142440 35520 142600 35680
rect 142440 35680 142600 35840
rect 142440 35840 142600 36000
rect 142440 36000 142600 36160
rect 142440 36160 142600 36320
rect 142440 36320 142600 36480
rect 142440 36480 142600 36640
rect 142440 36640 142600 36800
rect 142440 36800 142600 36960
rect 142440 36960 142600 37120
rect 142440 37120 142600 37280
rect 142440 37280 142600 37440
rect 142440 37440 142600 37600
rect 142440 37600 142600 37760
rect 142440 37760 142600 37920
rect 142440 37920 142600 38080
rect 142440 38080 142600 38240
rect 142440 38240 142600 38400
rect 142440 38400 142600 38560
rect 142440 38560 142600 38720
rect 142440 38720 142600 38880
rect 142440 38880 142600 39040
rect 142440 39040 142600 39200
rect 142440 39200 142600 39360
rect 142440 39360 142600 39520
rect 142440 39520 142600 39680
rect 142440 39680 142600 39840
rect 142440 39840 142600 40000
rect 142440 40000 142600 40160
rect 142440 40160 142600 40320
rect 142440 40320 142600 40480
rect 142440 40480 142600 40640
rect 142440 40640 142600 40800
rect 142440 40800 142600 40960
rect 142440 40960 142600 41120
rect 142440 41120 142600 41280
rect 142440 41280 142600 41440
rect 142440 41440 142600 41600
rect 142440 41600 142600 41760
rect 142440 41760 142600 41920
rect 142440 41920 142600 42080
rect 142440 42080 142600 42240
rect 142440 42240 142600 42400
rect 142440 42400 142600 42560
rect 142440 42560 142600 42720
rect 142440 42720 142600 42880
rect 142440 42880 142600 43040
rect 142440 43040 142600 43200
rect 142440 43200 142600 43360
rect 142440 43360 142600 43520
rect 142440 43520 142600 43680
rect 142440 43680 142600 43840
rect 142440 43840 142600 44000
rect 142440 44000 142600 44160
rect 142440 44160 142600 44320
rect 142440 44320 142600 44480
rect 142440 44480 142600 44640
rect 142440 44640 142600 44800
rect 142440 44800 142600 44960
rect 142440 44960 142600 45120
rect 142440 45120 142600 45280
rect 142440 45280 142600 45440
rect 142440 45440 142600 45600
rect 142440 45600 142600 45760
rect 142440 45760 142600 45920
rect 142440 45920 142600 46080
rect 142440 46080 142600 46240
rect 142440 46240 142600 46400
rect 142440 46400 142600 46560
rect 142440 46560 142600 46720
rect 142440 46720 142600 46880
rect 142440 46880 142600 47040
rect 142440 47040 142600 47200
rect 142440 47200 142600 47360
rect 142440 47360 142600 47520
rect 142440 47520 142600 47680
rect 142440 47680 142600 47840
rect 142440 47840 142600 48000
rect 142440 48000 142600 48160
rect 142440 48160 142600 48320
rect 142440 48320 142600 48480
rect 142440 48480 142600 48640
rect 142440 48640 142600 48800
rect 142440 48800 142600 48960
rect 142440 48960 142600 49120
rect 142440 49120 142600 49280
rect 142600 33760 142760 33920
rect 142600 33920 142760 34080
rect 142600 34080 142760 34240
rect 142600 34240 142760 34400
rect 142600 34400 142760 34560
rect 142600 34560 142760 34720
rect 142600 34720 142760 34880
rect 142600 34880 142760 35040
rect 142600 35040 142760 35200
rect 142600 35200 142760 35360
rect 142600 35360 142760 35520
rect 142600 35520 142760 35680
rect 142600 35680 142760 35840
rect 142600 35840 142760 36000
rect 142600 36000 142760 36160
rect 142600 36160 142760 36320
rect 142600 36320 142760 36480
rect 142600 36480 142760 36640
rect 142600 36640 142760 36800
rect 142600 36800 142760 36960
rect 142600 36960 142760 37120
rect 142600 37120 142760 37280
rect 142600 37280 142760 37440
rect 142600 37440 142760 37600
rect 142600 37600 142760 37760
rect 142600 37760 142760 37920
rect 142600 37920 142760 38080
rect 142600 38080 142760 38240
rect 142600 38240 142760 38400
rect 142600 38400 142760 38560
rect 142600 38560 142760 38720
rect 142600 38720 142760 38880
rect 142600 38880 142760 39040
rect 142600 39040 142760 39200
rect 142600 39200 142760 39360
rect 142600 39360 142760 39520
rect 142600 39520 142760 39680
rect 142600 39680 142760 39840
rect 142600 39840 142760 40000
rect 142600 40000 142760 40160
rect 142600 40160 142760 40320
rect 142600 40320 142760 40480
rect 142600 40480 142760 40640
rect 142600 40640 142760 40800
rect 142600 40800 142760 40960
rect 142600 40960 142760 41120
rect 142600 41120 142760 41280
rect 142600 41280 142760 41440
rect 142600 41440 142760 41600
rect 142600 41600 142760 41760
rect 142600 41760 142760 41920
rect 142600 41920 142760 42080
rect 142600 42080 142760 42240
rect 142600 42240 142760 42400
rect 142600 42400 142760 42560
rect 142600 42560 142760 42720
rect 142600 42720 142760 42880
rect 142600 42880 142760 43040
rect 142600 43040 142760 43200
rect 142600 43200 142760 43360
rect 142600 43360 142760 43520
rect 142600 43520 142760 43680
rect 142600 43680 142760 43840
rect 142600 43840 142760 44000
rect 142600 44000 142760 44160
rect 142600 44160 142760 44320
rect 142600 44320 142760 44480
rect 142600 44480 142760 44640
rect 142600 44640 142760 44800
rect 142600 44800 142760 44960
rect 142600 44960 142760 45120
rect 142600 45120 142760 45280
rect 142600 45280 142760 45440
rect 142600 45440 142760 45600
rect 142600 45600 142760 45760
rect 142600 45760 142760 45920
rect 142600 45920 142760 46080
rect 142600 46080 142760 46240
rect 142600 46240 142760 46400
rect 142600 46400 142760 46560
rect 142600 46560 142760 46720
rect 142600 46720 142760 46880
rect 142600 46880 142760 47040
rect 142600 47040 142760 47200
rect 142600 47200 142760 47360
rect 142600 47360 142760 47520
rect 142600 47520 142760 47680
rect 142600 47680 142760 47840
rect 142600 47840 142760 48000
rect 142600 48000 142760 48160
rect 142600 48160 142760 48320
rect 142600 48320 142760 48480
rect 142600 48480 142760 48640
rect 142600 48640 142760 48800
rect 142600 48800 142760 48960
rect 142760 34080 142920 34240
rect 142760 34240 142920 34400
rect 142760 34400 142920 34560
rect 142760 34560 142920 34720
rect 142760 34720 142920 34880
rect 142760 34880 142920 35040
rect 142760 35040 142920 35200
rect 142760 35200 142920 35360
rect 142760 35360 142920 35520
rect 142760 35520 142920 35680
rect 142760 35680 142920 35840
rect 142760 35840 142920 36000
rect 142760 36000 142920 36160
rect 142760 36160 142920 36320
rect 142760 36320 142920 36480
rect 142760 36480 142920 36640
rect 142760 36640 142920 36800
rect 142760 36800 142920 36960
rect 142760 36960 142920 37120
rect 142760 37120 142920 37280
rect 142760 37280 142920 37440
rect 142760 37440 142920 37600
rect 142760 37600 142920 37760
rect 142760 37760 142920 37920
rect 142760 37920 142920 38080
rect 142760 38080 142920 38240
rect 142760 38240 142920 38400
rect 142760 38400 142920 38560
rect 142760 38560 142920 38720
rect 142760 38720 142920 38880
rect 142760 38880 142920 39040
rect 142760 39040 142920 39200
rect 142760 39200 142920 39360
rect 142760 39360 142920 39520
rect 142760 39520 142920 39680
rect 142760 39680 142920 39840
rect 142760 39840 142920 40000
rect 142760 40000 142920 40160
rect 142760 40160 142920 40320
rect 142760 40320 142920 40480
rect 142760 40480 142920 40640
rect 142760 40640 142920 40800
rect 142760 40800 142920 40960
rect 142760 40960 142920 41120
rect 142760 41120 142920 41280
rect 142760 41280 142920 41440
rect 142760 41440 142920 41600
rect 142760 41600 142920 41760
rect 142760 41760 142920 41920
rect 142760 41920 142920 42080
rect 142760 42080 142920 42240
rect 142760 42240 142920 42400
rect 142760 42400 142920 42560
rect 142760 42560 142920 42720
rect 142760 42720 142920 42880
rect 142760 42880 142920 43040
rect 142760 43040 142920 43200
rect 142760 43200 142920 43360
rect 142760 43360 142920 43520
rect 142760 43520 142920 43680
rect 142760 43680 142920 43840
rect 142760 43840 142920 44000
rect 142760 44000 142920 44160
rect 142760 44160 142920 44320
rect 142760 44320 142920 44480
rect 142760 44480 142920 44640
rect 142760 44640 142920 44800
rect 142760 44800 142920 44960
rect 142760 44960 142920 45120
rect 142760 45120 142920 45280
rect 142760 45280 142920 45440
rect 142760 45440 142920 45600
rect 142760 45600 142920 45760
rect 142760 45760 142920 45920
rect 142760 45920 142920 46080
rect 142760 46080 142920 46240
rect 142760 46240 142920 46400
rect 142760 46400 142920 46560
rect 142760 46560 142920 46720
rect 142760 46720 142920 46880
rect 142760 46880 142920 47040
rect 142760 47040 142920 47200
rect 142760 47200 142920 47360
rect 142760 47360 142920 47520
rect 142760 47520 142920 47680
rect 142760 47680 142920 47840
rect 142760 47840 142920 48000
rect 142760 48000 142920 48160
rect 142760 48160 142920 48320
rect 142760 48320 142920 48480
rect 142760 48480 142920 48640
rect 142920 34560 143080 34720
rect 142920 34720 143080 34880
rect 142920 34880 143080 35040
rect 142920 35040 143080 35200
rect 142920 35200 143080 35360
rect 142920 35360 143080 35520
rect 142920 35520 143080 35680
rect 142920 35680 143080 35840
rect 142920 35840 143080 36000
rect 142920 36000 143080 36160
rect 142920 36160 143080 36320
rect 142920 36320 143080 36480
rect 142920 36480 143080 36640
rect 142920 36640 143080 36800
rect 142920 36800 143080 36960
rect 142920 36960 143080 37120
rect 142920 37120 143080 37280
rect 142920 37280 143080 37440
rect 142920 37440 143080 37600
rect 142920 37600 143080 37760
rect 142920 37760 143080 37920
rect 142920 37920 143080 38080
rect 142920 38080 143080 38240
rect 142920 38240 143080 38400
rect 142920 38400 143080 38560
rect 142920 38560 143080 38720
rect 142920 38720 143080 38880
rect 142920 38880 143080 39040
rect 142920 39040 143080 39200
rect 142920 39200 143080 39360
rect 142920 39360 143080 39520
rect 142920 39520 143080 39680
rect 142920 39680 143080 39840
rect 142920 39840 143080 40000
rect 142920 40000 143080 40160
rect 142920 40160 143080 40320
rect 142920 40320 143080 40480
rect 142920 40480 143080 40640
rect 142920 40640 143080 40800
rect 142920 40800 143080 40960
rect 142920 40960 143080 41120
rect 142920 41120 143080 41280
rect 142920 41280 143080 41440
rect 142920 41440 143080 41600
rect 142920 41600 143080 41760
rect 142920 41760 143080 41920
rect 142920 41920 143080 42080
rect 142920 42080 143080 42240
rect 142920 42240 143080 42400
rect 142920 42400 143080 42560
rect 142920 42560 143080 42720
rect 142920 42720 143080 42880
rect 142920 42880 143080 43040
rect 142920 43040 143080 43200
rect 142920 43200 143080 43360
rect 142920 43360 143080 43520
rect 142920 43520 143080 43680
rect 142920 43680 143080 43840
rect 142920 43840 143080 44000
rect 142920 44000 143080 44160
rect 142920 44160 143080 44320
rect 142920 44320 143080 44480
rect 142920 44480 143080 44640
rect 142920 44640 143080 44800
rect 142920 44800 143080 44960
rect 142920 44960 143080 45120
rect 142920 45120 143080 45280
rect 142920 45280 143080 45440
rect 142920 45440 143080 45600
rect 142920 45600 143080 45760
rect 142920 45760 143080 45920
rect 142920 45920 143080 46080
rect 142920 46080 143080 46240
rect 142920 46240 143080 46400
rect 142920 46400 143080 46560
rect 142920 46560 143080 46720
rect 142920 46720 143080 46880
rect 142920 46880 143080 47040
rect 142920 47040 143080 47200
rect 142920 47200 143080 47360
rect 142920 47360 143080 47520
rect 142920 47520 143080 47680
rect 142920 47680 143080 47840
rect 142920 47840 143080 48000
rect 142920 48000 143080 48160
rect 142920 48160 143080 48320
rect 143080 34880 143240 35040
rect 143080 35040 143240 35200
rect 143080 35200 143240 35360
rect 143080 35360 143240 35520
rect 143080 35520 143240 35680
rect 143080 35680 143240 35840
rect 143080 35840 143240 36000
rect 143080 36000 143240 36160
rect 143080 36160 143240 36320
rect 143080 36320 143240 36480
rect 143080 36480 143240 36640
rect 143080 36640 143240 36800
rect 143080 36800 143240 36960
rect 143080 36960 143240 37120
rect 143080 37120 143240 37280
rect 143080 37280 143240 37440
rect 143080 37440 143240 37600
rect 143080 37600 143240 37760
rect 143080 37760 143240 37920
rect 143080 37920 143240 38080
rect 143080 38080 143240 38240
rect 143080 38240 143240 38400
rect 143080 38400 143240 38560
rect 143080 38560 143240 38720
rect 143080 38720 143240 38880
rect 143080 38880 143240 39040
rect 143080 39040 143240 39200
rect 143080 39200 143240 39360
rect 143080 39360 143240 39520
rect 143080 39520 143240 39680
rect 143080 39680 143240 39840
rect 143080 39840 143240 40000
rect 143080 40000 143240 40160
rect 143080 40160 143240 40320
rect 143080 40320 143240 40480
rect 143080 40480 143240 40640
rect 143080 40640 143240 40800
rect 143080 40800 143240 40960
rect 143080 40960 143240 41120
rect 143080 41120 143240 41280
rect 143080 41280 143240 41440
rect 143080 41440 143240 41600
rect 143080 41600 143240 41760
rect 143080 41760 143240 41920
rect 143080 41920 143240 42080
rect 143080 42080 143240 42240
rect 143080 42240 143240 42400
rect 143080 42400 143240 42560
rect 143080 42560 143240 42720
rect 143080 42720 143240 42880
rect 143080 42880 143240 43040
rect 143080 43040 143240 43200
rect 143080 43200 143240 43360
rect 143080 43360 143240 43520
rect 143080 43520 143240 43680
rect 143080 43680 143240 43840
rect 143080 43840 143240 44000
rect 143080 44000 143240 44160
rect 143080 44160 143240 44320
rect 143080 44320 143240 44480
rect 143080 44480 143240 44640
rect 143080 44640 143240 44800
rect 143080 44800 143240 44960
rect 143080 44960 143240 45120
rect 143080 45120 143240 45280
rect 143080 45280 143240 45440
rect 143080 45440 143240 45600
rect 143080 45600 143240 45760
rect 143080 45760 143240 45920
rect 143080 45920 143240 46080
rect 143080 46080 143240 46240
rect 143080 46240 143240 46400
rect 143080 46400 143240 46560
rect 143080 46560 143240 46720
rect 143080 46720 143240 46880
rect 143080 46880 143240 47040
rect 143080 47040 143240 47200
rect 143080 47200 143240 47360
rect 143080 47360 143240 47520
rect 143080 47520 143240 47680
rect 143080 47680 143240 47840
rect 143240 35360 143400 35520
rect 143240 35520 143400 35680
rect 143240 35680 143400 35840
rect 143240 35840 143400 36000
rect 143240 36000 143400 36160
rect 143240 36160 143400 36320
rect 143240 36320 143400 36480
rect 143240 36480 143400 36640
rect 143240 36640 143400 36800
rect 143240 36800 143400 36960
rect 143240 36960 143400 37120
rect 143240 37120 143400 37280
rect 143240 37280 143400 37440
rect 143240 37440 143400 37600
rect 143240 37600 143400 37760
rect 143240 37760 143400 37920
rect 143240 37920 143400 38080
rect 143240 38080 143400 38240
rect 143240 38240 143400 38400
rect 143240 38400 143400 38560
rect 143240 38560 143400 38720
rect 143240 38720 143400 38880
rect 143240 38880 143400 39040
rect 143240 39040 143400 39200
rect 143240 39200 143400 39360
rect 143240 39360 143400 39520
rect 143240 39520 143400 39680
rect 143240 39680 143400 39840
rect 143240 39840 143400 40000
rect 143240 40000 143400 40160
rect 143240 40160 143400 40320
rect 143240 40320 143400 40480
rect 143240 40480 143400 40640
rect 143240 40640 143400 40800
rect 143240 40800 143400 40960
rect 143240 40960 143400 41120
rect 143240 41120 143400 41280
rect 143240 41280 143400 41440
rect 143240 41440 143400 41600
rect 143240 41600 143400 41760
rect 143240 41760 143400 41920
rect 143240 41920 143400 42080
rect 143240 42080 143400 42240
rect 143240 42240 143400 42400
rect 143240 42400 143400 42560
rect 143240 42560 143400 42720
rect 143240 42720 143400 42880
rect 143240 42880 143400 43040
rect 143240 43040 143400 43200
rect 143240 43200 143400 43360
rect 143240 43360 143400 43520
rect 143240 43520 143400 43680
rect 143240 43680 143400 43840
rect 143240 43840 143400 44000
rect 143240 44000 143400 44160
rect 143240 44160 143400 44320
rect 143240 44320 143400 44480
rect 143240 44480 143400 44640
rect 143240 44640 143400 44800
rect 143240 44800 143400 44960
rect 143240 44960 143400 45120
rect 143240 45120 143400 45280
rect 143240 45280 143400 45440
rect 143240 45440 143400 45600
rect 143240 45600 143400 45760
rect 143240 45760 143400 45920
rect 143240 45920 143400 46080
rect 143240 46080 143400 46240
rect 143240 46240 143400 46400
rect 143240 46400 143400 46560
rect 143240 46560 143400 46720
rect 143240 46720 143400 46880
rect 143240 46880 143400 47040
rect 143240 47040 143400 47200
rect 143240 47200 143400 47360
rect 143400 36000 143560 36160
rect 143400 36160 143560 36320
rect 143400 36320 143560 36480
rect 143400 36480 143560 36640
rect 143400 36640 143560 36800
rect 143400 36800 143560 36960
rect 143400 36960 143560 37120
rect 143400 37120 143560 37280
rect 143400 37280 143560 37440
rect 143400 37440 143560 37600
rect 143400 37600 143560 37760
rect 143400 37760 143560 37920
rect 143400 37920 143560 38080
rect 143400 38080 143560 38240
rect 143400 38240 143560 38400
rect 143400 38400 143560 38560
rect 143400 38560 143560 38720
rect 143400 38720 143560 38880
rect 143400 38880 143560 39040
rect 143400 39040 143560 39200
rect 143400 39200 143560 39360
rect 143400 39360 143560 39520
rect 143400 39520 143560 39680
rect 143400 39680 143560 39840
rect 143400 39840 143560 40000
rect 143400 40000 143560 40160
rect 143400 40160 143560 40320
rect 143400 40320 143560 40480
rect 143400 40480 143560 40640
rect 143400 40640 143560 40800
rect 143400 40800 143560 40960
rect 143400 40960 143560 41120
rect 143400 41120 143560 41280
rect 143400 41280 143560 41440
rect 143400 41440 143560 41600
rect 143400 41600 143560 41760
rect 143400 41760 143560 41920
rect 143400 41920 143560 42080
rect 143400 42080 143560 42240
rect 143400 42240 143560 42400
rect 143400 42400 143560 42560
rect 143400 42560 143560 42720
rect 143400 42720 143560 42880
rect 143400 42880 143560 43040
rect 143400 43040 143560 43200
rect 143400 43200 143560 43360
rect 143400 43360 143560 43520
rect 143400 43520 143560 43680
rect 143400 43680 143560 43840
rect 143400 43840 143560 44000
rect 143400 44000 143560 44160
rect 143400 44160 143560 44320
rect 143400 44320 143560 44480
rect 143400 44480 143560 44640
rect 143400 44640 143560 44800
rect 143400 44800 143560 44960
rect 143400 44960 143560 45120
rect 143400 45120 143560 45280
rect 143400 45280 143560 45440
rect 143400 45440 143560 45600
rect 143400 45600 143560 45760
rect 143400 45760 143560 45920
rect 143400 45920 143560 46080
rect 143400 46080 143560 46240
rect 143400 46240 143560 46400
rect 143400 46400 143560 46560
rect 143400 46560 143560 46720
rect 143400 46720 143560 46880
rect 143560 36480 143720 36640
rect 143560 36640 143720 36800
rect 143560 36800 143720 36960
rect 143560 36960 143720 37120
rect 143560 37120 143720 37280
rect 143560 37280 143720 37440
rect 143560 37440 143720 37600
rect 143560 37600 143720 37760
rect 143560 37760 143720 37920
rect 143560 37920 143720 38080
rect 143560 38080 143720 38240
rect 143560 38240 143720 38400
rect 143560 38400 143720 38560
rect 143560 38560 143720 38720
rect 143560 38720 143720 38880
rect 143560 38880 143720 39040
rect 143560 39040 143720 39200
rect 143560 39200 143720 39360
rect 143560 39360 143720 39520
rect 143560 39520 143720 39680
rect 143560 39680 143720 39840
rect 143560 39840 143720 40000
rect 143560 40000 143720 40160
rect 143560 40160 143720 40320
rect 143560 40320 143720 40480
rect 143560 40480 143720 40640
rect 143560 40640 143720 40800
rect 143560 40800 143720 40960
rect 143560 40960 143720 41120
rect 143560 41120 143720 41280
rect 143560 41280 143720 41440
rect 143560 41440 143720 41600
rect 143560 41600 143720 41760
rect 143560 41760 143720 41920
rect 143560 41920 143720 42080
rect 143560 42080 143720 42240
rect 143560 42240 143720 42400
rect 143560 42400 143720 42560
rect 143560 42560 143720 42720
rect 143560 42720 143720 42880
rect 143560 42880 143720 43040
rect 143560 43040 143720 43200
rect 143560 43200 143720 43360
rect 143560 43360 143720 43520
rect 143560 43520 143720 43680
rect 143560 43680 143720 43840
rect 143560 43840 143720 44000
rect 143560 44000 143720 44160
rect 143560 44160 143720 44320
rect 143560 44320 143720 44480
rect 143560 44480 143720 44640
rect 143560 44640 143720 44800
rect 143560 44800 143720 44960
rect 143560 44960 143720 45120
rect 143560 45120 143720 45280
rect 143560 45280 143720 45440
rect 143560 45440 143720 45600
rect 143560 45600 143720 45760
rect 143560 45760 143720 45920
rect 143560 45920 143720 46080
rect 143560 46080 143720 46240
rect 143720 37280 143880 37440
rect 143720 37440 143880 37600
rect 143720 37600 143880 37760
rect 143720 37760 143880 37920
rect 143720 37920 143880 38080
rect 143720 38080 143880 38240
rect 143720 38240 143880 38400
rect 143720 38400 143880 38560
rect 143720 38560 143880 38720
rect 143720 38720 143880 38880
rect 143720 38880 143880 39040
rect 143720 39040 143880 39200
rect 143720 39200 143880 39360
rect 143720 39360 143880 39520
rect 143720 39520 143880 39680
rect 143720 39680 143880 39840
rect 143720 39840 143880 40000
rect 143720 40000 143880 40160
rect 143720 40160 143880 40320
rect 143720 40320 143880 40480
rect 143720 40480 143880 40640
rect 143720 40640 143880 40800
rect 143720 40800 143880 40960
rect 143720 40960 143880 41120
rect 143720 41120 143880 41280
rect 143720 41280 143880 41440
rect 143720 41440 143880 41600
rect 143720 41600 143880 41760
rect 143720 41760 143880 41920
rect 143720 41920 143880 42080
rect 143720 42080 143880 42240
rect 143720 42240 143880 42400
rect 143720 42400 143880 42560
rect 143720 42560 143880 42720
rect 143720 42720 143880 42880
rect 143720 42880 143880 43040
rect 143720 43040 143880 43200
rect 143720 43200 143880 43360
rect 143720 43360 143880 43520
rect 143720 43520 143880 43680
rect 143720 43680 143880 43840
rect 143720 43840 143880 44000
rect 143720 44000 143880 44160
rect 143720 44160 143880 44320
rect 143720 44320 143880 44480
rect 143720 44480 143880 44640
rect 143720 44640 143880 44800
rect 143720 44800 143880 44960
rect 143720 44960 143880 45120
rect 143720 45120 143880 45280
rect 143720 45280 143880 45440
rect 143720 45440 143880 45600
rect 143880 38080 144040 38240
rect 143880 38240 144040 38400
rect 143880 38400 144040 38560
rect 143880 38560 144040 38720
rect 143880 38720 144040 38880
rect 143880 38880 144040 39040
rect 143880 39040 144040 39200
rect 143880 39200 144040 39360
rect 143880 39360 144040 39520
rect 143880 39520 144040 39680
rect 143880 39680 144040 39840
rect 143880 39840 144040 40000
rect 143880 40000 144040 40160
rect 143880 40160 144040 40320
rect 143880 40320 144040 40480
rect 143880 40480 144040 40640
rect 143880 40640 144040 40800
rect 143880 40800 144040 40960
rect 143880 40960 144040 41120
rect 143880 41120 144040 41280
rect 143880 41280 144040 41440
rect 143880 41440 144040 41600
rect 143880 41600 144040 41760
rect 143880 41760 144040 41920
rect 143880 41920 144040 42080
rect 143880 42080 144040 42240
rect 143880 42240 144040 42400
rect 143880 42400 144040 42560
rect 143880 42560 144040 42720
rect 143880 42720 144040 42880
rect 143880 42880 144040 43040
rect 143880 43040 144040 43200
rect 143880 43200 144040 43360
rect 143880 43360 144040 43520
rect 143880 43520 144040 43680
rect 143880 43680 144040 43840
rect 143880 43840 144040 44000
rect 143880 44000 144040 44160
rect 143880 44160 144040 44320
rect 143880 44320 144040 44480
rect 143880 44480 144040 44640
rect 144040 39200 144200 39360
rect 144040 39360 144200 39520
rect 144040 39520 144200 39680
rect 144040 39680 144200 39840
rect 144040 39840 144200 40000
rect 144040 40000 144200 40160
rect 144040 40160 144200 40320
rect 144040 40320 144200 40480
rect 144040 40480 144200 40640
rect 144040 40640 144200 40800
rect 144040 40800 144200 40960
rect 144040 40960 144200 41120
rect 144040 41120 144200 41280
rect 144040 41280 144200 41440
rect 144040 41440 144200 41600
rect 144040 41600 144200 41760
rect 144040 41760 144200 41920
rect 144040 41920 144200 42080
rect 144040 42080 144200 42240
rect 144040 42240 144200 42400
rect 144040 42400 144200 42560
rect 144040 42560 144200 42720
rect 144040 42720 144200 42880
rect 144040 42880 144200 43040
rect 144040 43040 144200 43200
rect 144040 43200 144200 43360
rect 148840 38560 149000 38720
rect 148840 38720 149000 38880
rect 148840 38880 149000 39040
rect 148840 39040 149000 39200
rect 148840 39200 149000 39360
rect 148840 39360 149000 39520
rect 148840 39520 149000 39680
rect 148840 39680 149000 39840
rect 148840 39840 149000 40000
rect 148840 40000 149000 40160
rect 149000 38080 149160 38240
rect 149000 38240 149160 38400
rect 149000 38400 149160 38560
rect 149000 38560 149160 38720
rect 149000 38720 149160 38880
rect 149000 38880 149160 39040
rect 149000 39040 149160 39200
rect 149000 39200 149160 39360
rect 149000 39360 149160 39520
rect 149000 39520 149160 39680
rect 149000 39680 149160 39840
rect 149000 39840 149160 40000
rect 149000 40000 149160 40160
rect 149000 40160 149160 40320
rect 149000 40320 149160 40480
rect 149000 40480 149160 40640
rect 149160 37920 149320 38080
rect 149160 38080 149320 38240
rect 149160 38240 149320 38400
rect 149160 38400 149320 38560
rect 149160 38560 149320 38720
rect 149160 38720 149320 38880
rect 149160 38880 149320 39040
rect 149160 39040 149320 39200
rect 149160 39200 149320 39360
rect 149160 39360 149320 39520
rect 149160 39520 149320 39680
rect 149160 39680 149320 39840
rect 149160 39840 149320 40000
rect 149160 40000 149320 40160
rect 149160 40160 149320 40320
rect 149160 40320 149320 40480
rect 149160 40480 149320 40640
rect 149160 40640 149320 40800
rect 149160 40800 149320 40960
rect 149160 40960 149320 41120
rect 149320 27520 149480 27680
rect 149320 27680 149480 27840
rect 149320 27840 149480 28000
rect 149320 28000 149480 28160
rect 149320 28160 149480 28320
rect 149320 28320 149480 28480
rect 149320 28480 149480 28640
rect 149320 28640 149480 28800
rect 149320 28800 149480 28960
rect 149320 28960 149480 29120
rect 149320 29120 149480 29280
rect 149320 29280 149480 29440
rect 149320 29440 149480 29600
rect 149320 29600 149480 29760
rect 149320 29760 149480 29920
rect 149320 29920 149480 30080
rect 149320 30080 149480 30240
rect 149320 30240 149480 30400
rect 149320 30400 149480 30560
rect 149320 30560 149480 30720
rect 149320 30720 149480 30880
rect 149320 30880 149480 31040
rect 149320 31040 149480 31200
rect 149320 31200 149480 31360
rect 149320 31360 149480 31520
rect 149320 31520 149480 31680
rect 149320 31680 149480 31840
rect 149320 31840 149480 32000
rect 149320 32000 149480 32160
rect 149320 32160 149480 32320
rect 149320 32320 149480 32480
rect 149320 32480 149480 32640
rect 149320 32640 149480 32800
rect 149320 32800 149480 32960
rect 149320 32960 149480 33120
rect 149320 33280 149480 33440
rect 149320 33600 149480 33760
rect 149320 37600 149480 37760
rect 149320 37760 149480 37920
rect 149320 37920 149480 38080
rect 149320 38080 149480 38240
rect 149320 38240 149480 38400
rect 149320 38400 149480 38560
rect 149320 38560 149480 38720
rect 149320 38720 149480 38880
rect 149320 38880 149480 39040
rect 149320 39040 149480 39200
rect 149320 39200 149480 39360
rect 149320 39360 149480 39520
rect 149320 39520 149480 39680
rect 149320 39680 149480 39840
rect 149320 39840 149480 40000
rect 149320 40000 149480 40160
rect 149320 40160 149480 40320
rect 149320 40320 149480 40480
rect 149320 40480 149480 40640
rect 149320 40640 149480 40800
rect 149320 40800 149480 40960
rect 149320 40960 149480 41120
rect 149320 41120 149480 41280
rect 149320 41280 149480 41440
rect 149480 27040 149640 27200
rect 149480 27200 149640 27360
rect 149480 27360 149640 27520
rect 149480 27520 149640 27680
rect 149480 27680 149640 27840
rect 149480 27840 149640 28000
rect 149480 28000 149640 28160
rect 149480 28160 149640 28320
rect 149480 28320 149640 28480
rect 149480 28480 149640 28640
rect 149480 28640 149640 28800
rect 149480 28800 149640 28960
rect 149480 28960 149640 29120
rect 149480 29120 149640 29280
rect 149480 29280 149640 29440
rect 149480 29440 149640 29600
rect 149480 29600 149640 29760
rect 149480 29760 149640 29920
rect 149480 29920 149640 30080
rect 149480 30080 149640 30240
rect 149480 30240 149640 30400
rect 149480 30400 149640 30560
rect 149480 30560 149640 30720
rect 149480 30720 149640 30880
rect 149480 30880 149640 31040
rect 149480 31040 149640 31200
rect 149480 31200 149640 31360
rect 149480 31360 149640 31520
rect 149480 31520 149640 31680
rect 149480 31680 149640 31840
rect 149480 31840 149640 32000
rect 149480 32000 149640 32160
rect 149480 32160 149640 32320
rect 149480 32320 149640 32480
rect 149480 32480 149640 32640
rect 149480 32640 149640 32800
rect 149480 32800 149640 32960
rect 149480 32960 149640 33120
rect 149480 33120 149640 33280
rect 149480 33280 149640 33440
rect 149480 33440 149640 33600
rect 149480 33600 149640 33760
rect 149480 33760 149640 33920
rect 149480 33920 149640 34080
rect 149480 34080 149640 34240
rect 149480 34240 149640 34400
rect 149480 34400 149640 34560
rect 149480 34560 149640 34720
rect 149480 34720 149640 34880
rect 149480 34880 149640 35040
rect 149480 35040 149640 35200
rect 149480 35200 149640 35360
rect 149480 35360 149640 35520
rect 149480 35520 149640 35680
rect 149480 35680 149640 35840
rect 149480 35840 149640 36000
rect 149480 36000 149640 36160
rect 149480 36160 149640 36320
rect 149480 36320 149640 36480
rect 149480 36480 149640 36640
rect 149480 36640 149640 36800
rect 149480 36800 149640 36960
rect 149480 36960 149640 37120
rect 149480 37120 149640 37280
rect 149480 37280 149640 37440
rect 149480 37440 149640 37600
rect 149480 37600 149640 37760
rect 149480 37760 149640 37920
rect 149480 37920 149640 38080
rect 149480 38080 149640 38240
rect 149480 38240 149640 38400
rect 149480 38400 149640 38560
rect 149480 38560 149640 38720
rect 149480 38720 149640 38880
rect 149480 38880 149640 39040
rect 149480 39040 149640 39200
rect 149480 39200 149640 39360
rect 149480 39360 149640 39520
rect 149480 39520 149640 39680
rect 149480 39680 149640 39840
rect 149480 39840 149640 40000
rect 149480 40000 149640 40160
rect 149480 40160 149640 40320
rect 149480 40320 149640 40480
rect 149480 40480 149640 40640
rect 149480 40640 149640 40800
rect 149480 40800 149640 40960
rect 149480 40960 149640 41120
rect 149480 41120 149640 41280
rect 149480 41280 149640 41440
rect 149480 41440 149640 41600
rect 149480 41600 149640 41760
rect 149640 26720 149800 26880
rect 149640 26880 149800 27040
rect 149640 27040 149800 27200
rect 149640 27200 149800 27360
rect 149640 27360 149800 27520
rect 149640 27520 149800 27680
rect 149640 27680 149800 27840
rect 149640 27840 149800 28000
rect 149640 28000 149800 28160
rect 149640 28160 149800 28320
rect 149640 28320 149800 28480
rect 149640 28480 149800 28640
rect 149640 28640 149800 28800
rect 149640 28800 149800 28960
rect 149640 28960 149800 29120
rect 149640 29120 149800 29280
rect 149640 29280 149800 29440
rect 149640 29440 149800 29600
rect 149640 29600 149800 29760
rect 149640 29760 149800 29920
rect 149640 29920 149800 30080
rect 149640 30080 149800 30240
rect 149640 30240 149800 30400
rect 149640 30400 149800 30560
rect 149640 30560 149800 30720
rect 149640 30720 149800 30880
rect 149640 30880 149800 31040
rect 149640 31040 149800 31200
rect 149640 31200 149800 31360
rect 149640 31360 149800 31520
rect 149640 31520 149800 31680
rect 149640 31680 149800 31840
rect 149640 31840 149800 32000
rect 149640 32000 149800 32160
rect 149640 32160 149800 32320
rect 149640 32320 149800 32480
rect 149640 32480 149800 32640
rect 149640 32640 149800 32800
rect 149640 32800 149800 32960
rect 149640 32960 149800 33120
rect 149640 33120 149800 33280
rect 149640 33280 149800 33440
rect 149640 33440 149800 33600
rect 149640 33600 149800 33760
rect 149640 33760 149800 33920
rect 149640 33920 149800 34080
rect 149640 34080 149800 34240
rect 149640 34240 149800 34400
rect 149640 34400 149800 34560
rect 149640 34560 149800 34720
rect 149640 34720 149800 34880
rect 149640 34880 149800 35040
rect 149640 35040 149800 35200
rect 149640 35200 149800 35360
rect 149640 35360 149800 35520
rect 149640 35520 149800 35680
rect 149640 35680 149800 35840
rect 149640 35840 149800 36000
rect 149640 36000 149800 36160
rect 149640 36160 149800 36320
rect 149640 36320 149800 36480
rect 149640 36480 149800 36640
rect 149640 36640 149800 36800
rect 149640 36800 149800 36960
rect 149640 36960 149800 37120
rect 149640 37120 149800 37280
rect 149640 37280 149800 37440
rect 149640 37440 149800 37600
rect 149640 37600 149800 37760
rect 149640 37760 149800 37920
rect 149640 37920 149800 38080
rect 149640 38080 149800 38240
rect 149640 38240 149800 38400
rect 149640 38400 149800 38560
rect 149640 38560 149800 38720
rect 149640 38720 149800 38880
rect 149640 38880 149800 39040
rect 149640 39040 149800 39200
rect 149640 39200 149800 39360
rect 149640 39360 149800 39520
rect 149640 39520 149800 39680
rect 149640 39680 149800 39840
rect 149640 39840 149800 40000
rect 149640 40000 149800 40160
rect 149640 40160 149800 40320
rect 149640 40320 149800 40480
rect 149640 40480 149800 40640
rect 149640 40640 149800 40800
rect 149640 40800 149800 40960
rect 149640 40960 149800 41120
rect 149640 41120 149800 41280
rect 149640 41280 149800 41440
rect 149640 41440 149800 41600
rect 149640 41600 149800 41760
rect 149640 41760 149800 41920
rect 149640 41920 149800 42080
rect 149640 42080 149800 42240
rect 149640 42240 149800 42400
rect 149640 42400 149800 42560
rect 149640 42560 149800 42720
rect 149640 42720 149800 42880
rect 149640 42880 149800 43040
rect 149640 43040 149800 43200
rect 149640 43200 149800 43360
rect 149640 43360 149800 43520
rect 149640 43520 149800 43680
rect 149640 43680 149800 43840
rect 149640 43840 149800 44000
rect 149640 44000 149800 44160
rect 149640 44160 149800 44320
rect 149640 44320 149800 44480
rect 149640 44480 149800 44640
rect 149640 44640 149800 44800
rect 149640 44800 149800 44960
rect 149640 44960 149800 45120
rect 149640 45120 149800 45280
rect 149640 45280 149800 45440
rect 149640 45440 149800 45600
rect 149640 45600 149800 45760
rect 149640 45760 149800 45920
rect 149640 45920 149800 46080
rect 149640 46080 149800 46240
rect 149640 46400 149800 46560
rect 149640 46720 149800 46880
rect 149800 26560 149960 26720
rect 149800 26720 149960 26880
rect 149800 26880 149960 27040
rect 149800 27040 149960 27200
rect 149800 27200 149960 27360
rect 149800 27360 149960 27520
rect 149800 27520 149960 27680
rect 149800 27680 149960 27840
rect 149800 27840 149960 28000
rect 149800 28000 149960 28160
rect 149800 28160 149960 28320
rect 149800 28320 149960 28480
rect 149800 28480 149960 28640
rect 149800 28640 149960 28800
rect 149800 28800 149960 28960
rect 149800 28960 149960 29120
rect 149800 29120 149960 29280
rect 149800 29280 149960 29440
rect 149800 29440 149960 29600
rect 149800 29600 149960 29760
rect 149800 29760 149960 29920
rect 149800 29920 149960 30080
rect 149800 30080 149960 30240
rect 149800 30240 149960 30400
rect 149800 30400 149960 30560
rect 149800 30560 149960 30720
rect 149800 30720 149960 30880
rect 149800 30880 149960 31040
rect 149800 31040 149960 31200
rect 149800 31200 149960 31360
rect 149800 31360 149960 31520
rect 149800 31520 149960 31680
rect 149800 31680 149960 31840
rect 149800 31840 149960 32000
rect 149800 32000 149960 32160
rect 149800 32160 149960 32320
rect 149800 32320 149960 32480
rect 149800 32480 149960 32640
rect 149800 32640 149960 32800
rect 149800 32800 149960 32960
rect 149800 32960 149960 33120
rect 149800 33120 149960 33280
rect 149800 33280 149960 33440
rect 149800 33440 149960 33600
rect 149800 33600 149960 33760
rect 149800 33760 149960 33920
rect 149800 33920 149960 34080
rect 149800 34080 149960 34240
rect 149800 34240 149960 34400
rect 149800 34400 149960 34560
rect 149800 34560 149960 34720
rect 149800 34720 149960 34880
rect 149800 34880 149960 35040
rect 149800 35040 149960 35200
rect 149800 35200 149960 35360
rect 149800 35360 149960 35520
rect 149800 35520 149960 35680
rect 149800 35680 149960 35840
rect 149800 35840 149960 36000
rect 149800 36000 149960 36160
rect 149800 36160 149960 36320
rect 149800 36320 149960 36480
rect 149800 36480 149960 36640
rect 149800 36640 149960 36800
rect 149800 36800 149960 36960
rect 149800 36960 149960 37120
rect 149800 37120 149960 37280
rect 149800 37280 149960 37440
rect 149800 37440 149960 37600
rect 149800 37600 149960 37760
rect 149800 37760 149960 37920
rect 149800 37920 149960 38080
rect 149800 38080 149960 38240
rect 149800 38240 149960 38400
rect 149800 38400 149960 38560
rect 149800 38560 149960 38720
rect 149800 38720 149960 38880
rect 149800 38880 149960 39040
rect 149800 39040 149960 39200
rect 149800 39200 149960 39360
rect 149800 39360 149960 39520
rect 149800 39520 149960 39680
rect 149800 39680 149960 39840
rect 149800 39840 149960 40000
rect 149800 40000 149960 40160
rect 149800 40160 149960 40320
rect 149800 40320 149960 40480
rect 149800 40480 149960 40640
rect 149800 40640 149960 40800
rect 149800 40800 149960 40960
rect 149800 40960 149960 41120
rect 149800 41120 149960 41280
rect 149800 41280 149960 41440
rect 149800 41440 149960 41600
rect 149800 41600 149960 41760
rect 149800 41760 149960 41920
rect 149800 41920 149960 42080
rect 149800 42080 149960 42240
rect 149800 42240 149960 42400
rect 149800 42400 149960 42560
rect 149800 42560 149960 42720
rect 149800 42720 149960 42880
rect 149800 42880 149960 43040
rect 149800 43040 149960 43200
rect 149800 43200 149960 43360
rect 149800 43360 149960 43520
rect 149800 43520 149960 43680
rect 149800 43680 149960 43840
rect 149800 43840 149960 44000
rect 149800 44000 149960 44160
rect 149800 44160 149960 44320
rect 149800 44320 149960 44480
rect 149800 44480 149960 44640
rect 149800 44640 149960 44800
rect 149800 44800 149960 44960
rect 149800 44960 149960 45120
rect 149800 45120 149960 45280
rect 149800 45280 149960 45440
rect 149800 45440 149960 45600
rect 149800 45600 149960 45760
rect 149800 45760 149960 45920
rect 149800 45920 149960 46080
rect 149800 46080 149960 46240
rect 149800 46240 149960 46400
rect 149800 46400 149960 46560
rect 149800 46560 149960 46720
rect 149800 46720 149960 46880
rect 149800 46880 149960 47040
rect 149800 47040 149960 47200
rect 149800 47200 149960 47360
rect 149800 47360 149960 47520
rect 149800 47520 149960 47680
rect 149800 47680 149960 47840
rect 149800 47840 149960 48000
rect 149800 48000 149960 48160
rect 149800 48160 149960 48320
rect 149800 48320 149960 48480
rect 149800 48480 149960 48640
rect 149800 48640 149960 48800
rect 149800 48800 149960 48960
rect 149800 48960 149960 49120
rect 149800 49120 149960 49280
rect 149800 49280 149960 49440
rect 149800 49440 149960 49600
rect 149800 49600 149960 49760
rect 149800 49760 149960 49920
rect 149800 49920 149960 50080
rect 149800 50080 149960 50240
rect 149800 50240 149960 50400
rect 149800 50400 149960 50560
rect 149800 50560 149960 50720
rect 149800 50720 149960 50880
rect 149800 50880 149960 51040
rect 149800 51040 149960 51200
rect 149800 51200 149960 51360
rect 149800 51360 149960 51520
rect 149800 51520 149960 51680
rect 149800 51680 149960 51840
rect 149800 51840 149960 52000
rect 149800 52000 149960 52160
rect 149960 26400 150120 26560
rect 149960 26560 150120 26720
rect 149960 26720 150120 26880
rect 149960 26880 150120 27040
rect 149960 27040 150120 27200
rect 149960 27200 150120 27360
rect 149960 27360 150120 27520
rect 149960 27520 150120 27680
rect 149960 27680 150120 27840
rect 149960 27840 150120 28000
rect 149960 28000 150120 28160
rect 149960 28160 150120 28320
rect 149960 28320 150120 28480
rect 149960 28480 150120 28640
rect 149960 28640 150120 28800
rect 149960 28800 150120 28960
rect 149960 28960 150120 29120
rect 149960 29120 150120 29280
rect 149960 29280 150120 29440
rect 149960 29440 150120 29600
rect 149960 29600 150120 29760
rect 149960 29760 150120 29920
rect 149960 29920 150120 30080
rect 149960 30080 150120 30240
rect 149960 30240 150120 30400
rect 149960 30400 150120 30560
rect 149960 30560 150120 30720
rect 149960 30720 150120 30880
rect 149960 30880 150120 31040
rect 149960 31040 150120 31200
rect 149960 31200 150120 31360
rect 149960 31360 150120 31520
rect 149960 31520 150120 31680
rect 149960 31680 150120 31840
rect 149960 31840 150120 32000
rect 149960 32000 150120 32160
rect 149960 32160 150120 32320
rect 149960 32320 150120 32480
rect 149960 32480 150120 32640
rect 149960 32640 150120 32800
rect 149960 32800 150120 32960
rect 149960 32960 150120 33120
rect 149960 33120 150120 33280
rect 149960 33280 150120 33440
rect 149960 33440 150120 33600
rect 149960 33600 150120 33760
rect 149960 33760 150120 33920
rect 149960 33920 150120 34080
rect 149960 34080 150120 34240
rect 149960 34240 150120 34400
rect 149960 34400 150120 34560
rect 149960 34560 150120 34720
rect 149960 34720 150120 34880
rect 149960 34880 150120 35040
rect 149960 35040 150120 35200
rect 149960 35200 150120 35360
rect 149960 35360 150120 35520
rect 149960 35520 150120 35680
rect 149960 35680 150120 35840
rect 149960 35840 150120 36000
rect 149960 36000 150120 36160
rect 149960 36160 150120 36320
rect 149960 36320 150120 36480
rect 149960 36480 150120 36640
rect 149960 36640 150120 36800
rect 149960 36800 150120 36960
rect 149960 36960 150120 37120
rect 149960 37120 150120 37280
rect 149960 37280 150120 37440
rect 149960 37440 150120 37600
rect 149960 37600 150120 37760
rect 149960 37760 150120 37920
rect 149960 37920 150120 38080
rect 149960 38080 150120 38240
rect 149960 38240 150120 38400
rect 149960 38400 150120 38560
rect 149960 38560 150120 38720
rect 149960 38720 150120 38880
rect 149960 38880 150120 39040
rect 149960 39040 150120 39200
rect 149960 39200 150120 39360
rect 149960 39360 150120 39520
rect 149960 39520 150120 39680
rect 149960 39680 150120 39840
rect 149960 39840 150120 40000
rect 149960 40000 150120 40160
rect 149960 40160 150120 40320
rect 149960 40320 150120 40480
rect 149960 40480 150120 40640
rect 149960 40640 150120 40800
rect 149960 40800 150120 40960
rect 149960 40960 150120 41120
rect 149960 41120 150120 41280
rect 149960 41280 150120 41440
rect 149960 41440 150120 41600
rect 149960 41600 150120 41760
rect 149960 41760 150120 41920
rect 149960 41920 150120 42080
rect 149960 42080 150120 42240
rect 149960 42240 150120 42400
rect 149960 42400 150120 42560
rect 149960 42560 150120 42720
rect 149960 42720 150120 42880
rect 149960 42880 150120 43040
rect 149960 43040 150120 43200
rect 149960 43200 150120 43360
rect 149960 43360 150120 43520
rect 149960 43520 150120 43680
rect 149960 43680 150120 43840
rect 149960 43840 150120 44000
rect 149960 44000 150120 44160
rect 149960 44160 150120 44320
rect 149960 44320 150120 44480
rect 149960 44480 150120 44640
rect 149960 44640 150120 44800
rect 149960 44800 150120 44960
rect 149960 44960 150120 45120
rect 149960 45120 150120 45280
rect 149960 45280 150120 45440
rect 149960 45440 150120 45600
rect 149960 45600 150120 45760
rect 149960 45760 150120 45920
rect 149960 45920 150120 46080
rect 149960 46080 150120 46240
rect 149960 46240 150120 46400
rect 149960 46400 150120 46560
rect 149960 46560 150120 46720
rect 149960 46720 150120 46880
rect 149960 46880 150120 47040
rect 149960 47040 150120 47200
rect 149960 47200 150120 47360
rect 149960 47360 150120 47520
rect 149960 47520 150120 47680
rect 149960 47680 150120 47840
rect 149960 47840 150120 48000
rect 149960 48000 150120 48160
rect 149960 48160 150120 48320
rect 149960 48320 150120 48480
rect 149960 48480 150120 48640
rect 149960 48640 150120 48800
rect 149960 48800 150120 48960
rect 149960 48960 150120 49120
rect 149960 49120 150120 49280
rect 149960 49280 150120 49440
rect 149960 49440 150120 49600
rect 149960 49600 150120 49760
rect 149960 49760 150120 49920
rect 149960 49920 150120 50080
rect 149960 50080 150120 50240
rect 149960 50240 150120 50400
rect 149960 50400 150120 50560
rect 149960 50560 150120 50720
rect 149960 50720 150120 50880
rect 149960 50880 150120 51040
rect 149960 51040 150120 51200
rect 149960 51200 150120 51360
rect 149960 51360 150120 51520
rect 149960 51520 150120 51680
rect 149960 51680 150120 51840
rect 149960 51840 150120 52000
rect 149960 52000 150120 52160
rect 149960 52160 150120 52320
rect 149960 52320 150120 52480
rect 149960 52480 150120 52640
rect 150120 26240 150280 26400
rect 150120 26400 150280 26560
rect 150120 26560 150280 26720
rect 150120 26720 150280 26880
rect 150120 26880 150280 27040
rect 150120 27040 150280 27200
rect 150120 27200 150280 27360
rect 150120 27360 150280 27520
rect 150120 27520 150280 27680
rect 150120 27680 150280 27840
rect 150120 27840 150280 28000
rect 150120 28000 150280 28160
rect 150120 28160 150280 28320
rect 150120 28320 150280 28480
rect 150120 28480 150280 28640
rect 150120 28640 150280 28800
rect 150120 28800 150280 28960
rect 150120 28960 150280 29120
rect 150120 29120 150280 29280
rect 150120 29280 150280 29440
rect 150120 29440 150280 29600
rect 150120 29600 150280 29760
rect 150120 29760 150280 29920
rect 150120 29920 150280 30080
rect 150120 30080 150280 30240
rect 150120 30240 150280 30400
rect 150120 30400 150280 30560
rect 150120 30560 150280 30720
rect 150120 30720 150280 30880
rect 150120 30880 150280 31040
rect 150120 31040 150280 31200
rect 150120 31200 150280 31360
rect 150120 31360 150280 31520
rect 150120 31520 150280 31680
rect 150120 31680 150280 31840
rect 150120 31840 150280 32000
rect 150120 32000 150280 32160
rect 150120 32160 150280 32320
rect 150120 32320 150280 32480
rect 150120 32480 150280 32640
rect 150120 32640 150280 32800
rect 150120 32800 150280 32960
rect 150120 32960 150280 33120
rect 150120 33120 150280 33280
rect 150120 33280 150280 33440
rect 150120 33440 150280 33600
rect 150120 33600 150280 33760
rect 150120 33760 150280 33920
rect 150120 33920 150280 34080
rect 150120 34080 150280 34240
rect 150120 34240 150280 34400
rect 150120 34400 150280 34560
rect 150120 34560 150280 34720
rect 150120 34720 150280 34880
rect 150120 34880 150280 35040
rect 150120 35040 150280 35200
rect 150120 35200 150280 35360
rect 150120 35360 150280 35520
rect 150120 35520 150280 35680
rect 150120 35680 150280 35840
rect 150120 35840 150280 36000
rect 150120 36000 150280 36160
rect 150120 36160 150280 36320
rect 150120 36320 150280 36480
rect 150120 36480 150280 36640
rect 150120 36640 150280 36800
rect 150120 36800 150280 36960
rect 150120 36960 150280 37120
rect 150120 37120 150280 37280
rect 150120 37280 150280 37440
rect 150120 37440 150280 37600
rect 150120 37600 150280 37760
rect 150120 37760 150280 37920
rect 150120 37920 150280 38080
rect 150120 38080 150280 38240
rect 150120 38240 150280 38400
rect 150120 38400 150280 38560
rect 150120 38560 150280 38720
rect 150120 38720 150280 38880
rect 150120 38880 150280 39040
rect 150120 39040 150280 39200
rect 150120 39200 150280 39360
rect 150120 39360 150280 39520
rect 150120 39520 150280 39680
rect 150120 39680 150280 39840
rect 150120 39840 150280 40000
rect 150120 40000 150280 40160
rect 150120 40160 150280 40320
rect 150120 40320 150280 40480
rect 150120 40480 150280 40640
rect 150120 40640 150280 40800
rect 150120 40800 150280 40960
rect 150120 40960 150280 41120
rect 150120 41120 150280 41280
rect 150120 41280 150280 41440
rect 150120 41440 150280 41600
rect 150120 41600 150280 41760
rect 150120 41760 150280 41920
rect 150120 41920 150280 42080
rect 150120 42080 150280 42240
rect 150120 42240 150280 42400
rect 150120 42400 150280 42560
rect 150120 42560 150280 42720
rect 150120 42720 150280 42880
rect 150120 42880 150280 43040
rect 150120 43040 150280 43200
rect 150120 43200 150280 43360
rect 150120 43360 150280 43520
rect 150120 43520 150280 43680
rect 150120 43680 150280 43840
rect 150120 43840 150280 44000
rect 150120 44000 150280 44160
rect 150120 44160 150280 44320
rect 150120 44320 150280 44480
rect 150120 44480 150280 44640
rect 150120 44640 150280 44800
rect 150120 44800 150280 44960
rect 150120 44960 150280 45120
rect 150120 45120 150280 45280
rect 150120 45280 150280 45440
rect 150120 45440 150280 45600
rect 150120 45600 150280 45760
rect 150120 45760 150280 45920
rect 150120 45920 150280 46080
rect 150120 46080 150280 46240
rect 150120 46240 150280 46400
rect 150120 46400 150280 46560
rect 150120 46560 150280 46720
rect 150120 46720 150280 46880
rect 150120 46880 150280 47040
rect 150120 47040 150280 47200
rect 150120 47200 150280 47360
rect 150120 47360 150280 47520
rect 150120 47520 150280 47680
rect 150120 47680 150280 47840
rect 150120 47840 150280 48000
rect 150120 48000 150280 48160
rect 150120 48160 150280 48320
rect 150120 48320 150280 48480
rect 150120 48480 150280 48640
rect 150120 48640 150280 48800
rect 150120 48800 150280 48960
rect 150120 48960 150280 49120
rect 150120 49120 150280 49280
rect 150120 49280 150280 49440
rect 150120 49440 150280 49600
rect 150120 49600 150280 49760
rect 150120 49760 150280 49920
rect 150120 49920 150280 50080
rect 150120 50080 150280 50240
rect 150120 50240 150280 50400
rect 150120 50400 150280 50560
rect 150120 50560 150280 50720
rect 150120 50720 150280 50880
rect 150120 50880 150280 51040
rect 150120 51040 150280 51200
rect 150120 51200 150280 51360
rect 150120 51360 150280 51520
rect 150120 51520 150280 51680
rect 150120 51680 150280 51840
rect 150120 51840 150280 52000
rect 150120 52000 150280 52160
rect 150120 52160 150280 52320
rect 150120 52320 150280 52480
rect 150120 52480 150280 52640
rect 150120 52640 150280 52800
rect 150280 26080 150440 26240
rect 150280 26240 150440 26400
rect 150280 26400 150440 26560
rect 150280 26560 150440 26720
rect 150280 26720 150440 26880
rect 150280 26880 150440 27040
rect 150280 27040 150440 27200
rect 150280 27200 150440 27360
rect 150280 27360 150440 27520
rect 150280 27520 150440 27680
rect 150280 27680 150440 27840
rect 150280 27840 150440 28000
rect 150280 28000 150440 28160
rect 150280 28160 150440 28320
rect 150280 28320 150440 28480
rect 150280 28480 150440 28640
rect 150280 28640 150440 28800
rect 150280 28800 150440 28960
rect 150280 28960 150440 29120
rect 150280 29120 150440 29280
rect 150280 29280 150440 29440
rect 150280 29440 150440 29600
rect 150280 29600 150440 29760
rect 150280 29760 150440 29920
rect 150280 29920 150440 30080
rect 150280 30080 150440 30240
rect 150280 30240 150440 30400
rect 150280 30400 150440 30560
rect 150280 30560 150440 30720
rect 150280 30720 150440 30880
rect 150280 30880 150440 31040
rect 150280 31040 150440 31200
rect 150280 31200 150440 31360
rect 150280 31360 150440 31520
rect 150280 31520 150440 31680
rect 150280 31680 150440 31840
rect 150280 31840 150440 32000
rect 150280 32000 150440 32160
rect 150280 32160 150440 32320
rect 150280 32320 150440 32480
rect 150280 32480 150440 32640
rect 150280 32640 150440 32800
rect 150280 32800 150440 32960
rect 150280 32960 150440 33120
rect 150280 33120 150440 33280
rect 150280 33280 150440 33440
rect 150280 33440 150440 33600
rect 150280 33600 150440 33760
rect 150280 33760 150440 33920
rect 150280 33920 150440 34080
rect 150280 34080 150440 34240
rect 150280 34240 150440 34400
rect 150280 34400 150440 34560
rect 150280 34560 150440 34720
rect 150280 34720 150440 34880
rect 150280 34880 150440 35040
rect 150280 35040 150440 35200
rect 150280 35200 150440 35360
rect 150280 35360 150440 35520
rect 150280 35520 150440 35680
rect 150280 35680 150440 35840
rect 150280 35840 150440 36000
rect 150280 36000 150440 36160
rect 150280 36160 150440 36320
rect 150280 36320 150440 36480
rect 150280 36480 150440 36640
rect 150280 36640 150440 36800
rect 150280 36800 150440 36960
rect 150280 36960 150440 37120
rect 150280 37120 150440 37280
rect 150280 37280 150440 37440
rect 150280 37440 150440 37600
rect 150280 37600 150440 37760
rect 150280 37760 150440 37920
rect 150280 37920 150440 38080
rect 150280 38080 150440 38240
rect 150280 38240 150440 38400
rect 150280 38400 150440 38560
rect 150280 38560 150440 38720
rect 150280 38720 150440 38880
rect 150280 38880 150440 39040
rect 150280 39040 150440 39200
rect 150280 39200 150440 39360
rect 150280 39360 150440 39520
rect 150280 39520 150440 39680
rect 150280 39680 150440 39840
rect 150280 39840 150440 40000
rect 150280 40000 150440 40160
rect 150280 40160 150440 40320
rect 150280 40320 150440 40480
rect 150280 40480 150440 40640
rect 150280 40640 150440 40800
rect 150280 40800 150440 40960
rect 150280 40960 150440 41120
rect 150280 41120 150440 41280
rect 150280 41280 150440 41440
rect 150280 41440 150440 41600
rect 150280 41600 150440 41760
rect 150280 41760 150440 41920
rect 150280 41920 150440 42080
rect 150280 42080 150440 42240
rect 150280 42240 150440 42400
rect 150280 42400 150440 42560
rect 150280 42560 150440 42720
rect 150280 42720 150440 42880
rect 150280 42880 150440 43040
rect 150280 43040 150440 43200
rect 150280 43200 150440 43360
rect 150280 43360 150440 43520
rect 150280 43520 150440 43680
rect 150280 43680 150440 43840
rect 150280 43840 150440 44000
rect 150280 44000 150440 44160
rect 150280 44160 150440 44320
rect 150280 44320 150440 44480
rect 150280 44480 150440 44640
rect 150280 44640 150440 44800
rect 150280 44800 150440 44960
rect 150280 44960 150440 45120
rect 150280 45120 150440 45280
rect 150280 45280 150440 45440
rect 150280 45440 150440 45600
rect 150280 45600 150440 45760
rect 150280 45760 150440 45920
rect 150280 45920 150440 46080
rect 150280 46080 150440 46240
rect 150280 46240 150440 46400
rect 150280 46400 150440 46560
rect 150280 46560 150440 46720
rect 150280 46720 150440 46880
rect 150280 46880 150440 47040
rect 150280 47040 150440 47200
rect 150280 47200 150440 47360
rect 150280 47360 150440 47520
rect 150280 47520 150440 47680
rect 150280 47680 150440 47840
rect 150280 47840 150440 48000
rect 150280 48000 150440 48160
rect 150280 48160 150440 48320
rect 150280 48320 150440 48480
rect 150280 48480 150440 48640
rect 150280 48640 150440 48800
rect 150280 48800 150440 48960
rect 150280 48960 150440 49120
rect 150280 49120 150440 49280
rect 150280 49280 150440 49440
rect 150280 49440 150440 49600
rect 150280 49600 150440 49760
rect 150280 49760 150440 49920
rect 150280 49920 150440 50080
rect 150280 50080 150440 50240
rect 150280 50240 150440 50400
rect 150280 50400 150440 50560
rect 150280 50560 150440 50720
rect 150280 50720 150440 50880
rect 150280 50880 150440 51040
rect 150280 51040 150440 51200
rect 150280 51200 150440 51360
rect 150280 51360 150440 51520
rect 150280 51520 150440 51680
rect 150280 51680 150440 51840
rect 150280 51840 150440 52000
rect 150280 52000 150440 52160
rect 150280 52160 150440 52320
rect 150280 52320 150440 52480
rect 150280 52480 150440 52640
rect 150280 52640 150440 52800
rect 150280 52800 150440 52960
rect 150440 25920 150600 26080
rect 150440 26080 150600 26240
rect 150440 26240 150600 26400
rect 150440 26400 150600 26560
rect 150440 26560 150600 26720
rect 150440 26720 150600 26880
rect 150440 26880 150600 27040
rect 150440 27040 150600 27200
rect 150440 27200 150600 27360
rect 150440 27360 150600 27520
rect 150440 27520 150600 27680
rect 150440 27680 150600 27840
rect 150440 27840 150600 28000
rect 150440 28000 150600 28160
rect 150440 28160 150600 28320
rect 150440 28320 150600 28480
rect 150440 28480 150600 28640
rect 150440 28640 150600 28800
rect 150440 28800 150600 28960
rect 150440 28960 150600 29120
rect 150440 29120 150600 29280
rect 150440 29280 150600 29440
rect 150440 29440 150600 29600
rect 150440 29600 150600 29760
rect 150440 29760 150600 29920
rect 150440 29920 150600 30080
rect 150440 30080 150600 30240
rect 150440 30240 150600 30400
rect 150440 30400 150600 30560
rect 150440 30560 150600 30720
rect 150440 30720 150600 30880
rect 150440 30880 150600 31040
rect 150440 31040 150600 31200
rect 150440 31200 150600 31360
rect 150440 31360 150600 31520
rect 150440 31520 150600 31680
rect 150440 31680 150600 31840
rect 150440 31840 150600 32000
rect 150440 32000 150600 32160
rect 150440 32160 150600 32320
rect 150440 32320 150600 32480
rect 150440 32480 150600 32640
rect 150440 32640 150600 32800
rect 150440 32800 150600 32960
rect 150440 32960 150600 33120
rect 150440 33120 150600 33280
rect 150440 33280 150600 33440
rect 150440 33440 150600 33600
rect 150440 33600 150600 33760
rect 150440 33760 150600 33920
rect 150440 33920 150600 34080
rect 150440 34080 150600 34240
rect 150440 34240 150600 34400
rect 150440 34400 150600 34560
rect 150440 34560 150600 34720
rect 150440 34720 150600 34880
rect 150440 34880 150600 35040
rect 150440 35040 150600 35200
rect 150440 35200 150600 35360
rect 150440 35360 150600 35520
rect 150440 35520 150600 35680
rect 150440 35680 150600 35840
rect 150440 35840 150600 36000
rect 150440 36000 150600 36160
rect 150440 36160 150600 36320
rect 150440 36320 150600 36480
rect 150440 36480 150600 36640
rect 150440 36640 150600 36800
rect 150440 36800 150600 36960
rect 150440 36960 150600 37120
rect 150440 37120 150600 37280
rect 150440 37280 150600 37440
rect 150440 37440 150600 37600
rect 150440 37600 150600 37760
rect 150440 37760 150600 37920
rect 150440 37920 150600 38080
rect 150440 38080 150600 38240
rect 150440 38240 150600 38400
rect 150440 38400 150600 38560
rect 150440 38560 150600 38720
rect 150440 38720 150600 38880
rect 150440 38880 150600 39040
rect 150440 39040 150600 39200
rect 150440 39200 150600 39360
rect 150440 39360 150600 39520
rect 150440 39520 150600 39680
rect 150440 39680 150600 39840
rect 150440 39840 150600 40000
rect 150440 40000 150600 40160
rect 150440 40160 150600 40320
rect 150440 40320 150600 40480
rect 150440 40480 150600 40640
rect 150440 40640 150600 40800
rect 150440 40800 150600 40960
rect 150440 40960 150600 41120
rect 150440 41120 150600 41280
rect 150440 41280 150600 41440
rect 150440 41440 150600 41600
rect 150440 41600 150600 41760
rect 150440 41760 150600 41920
rect 150440 41920 150600 42080
rect 150440 42080 150600 42240
rect 150440 42240 150600 42400
rect 150440 42400 150600 42560
rect 150440 42560 150600 42720
rect 150440 42720 150600 42880
rect 150440 42880 150600 43040
rect 150440 43040 150600 43200
rect 150440 43200 150600 43360
rect 150440 43360 150600 43520
rect 150440 43520 150600 43680
rect 150440 43680 150600 43840
rect 150440 43840 150600 44000
rect 150440 44000 150600 44160
rect 150440 44160 150600 44320
rect 150440 44320 150600 44480
rect 150440 44480 150600 44640
rect 150440 44640 150600 44800
rect 150440 44800 150600 44960
rect 150440 44960 150600 45120
rect 150440 45120 150600 45280
rect 150440 45280 150600 45440
rect 150440 45440 150600 45600
rect 150440 45600 150600 45760
rect 150440 45760 150600 45920
rect 150440 45920 150600 46080
rect 150440 46080 150600 46240
rect 150440 46240 150600 46400
rect 150440 46400 150600 46560
rect 150440 46560 150600 46720
rect 150440 46720 150600 46880
rect 150440 46880 150600 47040
rect 150440 47040 150600 47200
rect 150440 47200 150600 47360
rect 150440 47360 150600 47520
rect 150440 47520 150600 47680
rect 150440 47680 150600 47840
rect 150440 47840 150600 48000
rect 150440 48000 150600 48160
rect 150440 48160 150600 48320
rect 150440 48320 150600 48480
rect 150440 48480 150600 48640
rect 150440 48640 150600 48800
rect 150440 48800 150600 48960
rect 150440 48960 150600 49120
rect 150440 49120 150600 49280
rect 150440 49280 150600 49440
rect 150440 49440 150600 49600
rect 150440 49600 150600 49760
rect 150440 49760 150600 49920
rect 150440 49920 150600 50080
rect 150440 50080 150600 50240
rect 150440 50240 150600 50400
rect 150440 50400 150600 50560
rect 150440 50560 150600 50720
rect 150440 50720 150600 50880
rect 150440 50880 150600 51040
rect 150440 51040 150600 51200
rect 150440 51200 150600 51360
rect 150440 51360 150600 51520
rect 150440 51520 150600 51680
rect 150440 51680 150600 51840
rect 150440 51840 150600 52000
rect 150440 52000 150600 52160
rect 150440 52160 150600 52320
rect 150440 52320 150600 52480
rect 150440 52480 150600 52640
rect 150440 52640 150600 52800
rect 150440 52800 150600 52960
rect 150440 52960 150600 53120
rect 150600 25920 150760 26080
rect 150600 26080 150760 26240
rect 150600 26240 150760 26400
rect 150600 26400 150760 26560
rect 150600 26560 150760 26720
rect 150600 26720 150760 26880
rect 150600 26880 150760 27040
rect 150600 27040 150760 27200
rect 150600 27200 150760 27360
rect 150600 27360 150760 27520
rect 150600 27520 150760 27680
rect 150600 27680 150760 27840
rect 150600 27840 150760 28000
rect 150600 28000 150760 28160
rect 150600 28160 150760 28320
rect 150600 28320 150760 28480
rect 150600 28480 150760 28640
rect 150600 28640 150760 28800
rect 150600 28800 150760 28960
rect 150600 28960 150760 29120
rect 150600 29120 150760 29280
rect 150600 29280 150760 29440
rect 150600 29440 150760 29600
rect 150600 29600 150760 29760
rect 150600 29760 150760 29920
rect 150600 29920 150760 30080
rect 150600 30080 150760 30240
rect 150600 30240 150760 30400
rect 150600 30400 150760 30560
rect 150600 30560 150760 30720
rect 150600 30720 150760 30880
rect 150600 30880 150760 31040
rect 150600 31040 150760 31200
rect 150600 31200 150760 31360
rect 150600 31360 150760 31520
rect 150600 31520 150760 31680
rect 150600 31680 150760 31840
rect 150600 31840 150760 32000
rect 150600 32000 150760 32160
rect 150600 32160 150760 32320
rect 150600 32320 150760 32480
rect 150600 32480 150760 32640
rect 150600 32640 150760 32800
rect 150600 32800 150760 32960
rect 150600 32960 150760 33120
rect 150600 33120 150760 33280
rect 150600 33280 150760 33440
rect 150600 33440 150760 33600
rect 150600 33600 150760 33760
rect 150600 33760 150760 33920
rect 150600 33920 150760 34080
rect 150600 34080 150760 34240
rect 150600 34240 150760 34400
rect 150600 34400 150760 34560
rect 150600 34560 150760 34720
rect 150600 34720 150760 34880
rect 150600 34880 150760 35040
rect 150600 35040 150760 35200
rect 150600 35200 150760 35360
rect 150600 35360 150760 35520
rect 150600 35520 150760 35680
rect 150600 35680 150760 35840
rect 150600 35840 150760 36000
rect 150600 36000 150760 36160
rect 150600 36160 150760 36320
rect 150600 36320 150760 36480
rect 150600 36480 150760 36640
rect 150600 36640 150760 36800
rect 150600 36800 150760 36960
rect 150600 36960 150760 37120
rect 150600 37120 150760 37280
rect 150600 37280 150760 37440
rect 150600 37440 150760 37600
rect 150600 37600 150760 37760
rect 150600 37760 150760 37920
rect 150600 37920 150760 38080
rect 150600 38080 150760 38240
rect 150600 38240 150760 38400
rect 150600 38400 150760 38560
rect 150600 38560 150760 38720
rect 150600 38720 150760 38880
rect 150600 38880 150760 39040
rect 150600 39040 150760 39200
rect 150600 39200 150760 39360
rect 150600 39360 150760 39520
rect 150600 39520 150760 39680
rect 150600 39680 150760 39840
rect 150600 39840 150760 40000
rect 150600 40000 150760 40160
rect 150600 40160 150760 40320
rect 150600 40320 150760 40480
rect 150600 40480 150760 40640
rect 150600 40640 150760 40800
rect 150600 40800 150760 40960
rect 150600 40960 150760 41120
rect 150600 41120 150760 41280
rect 150600 41280 150760 41440
rect 150600 41440 150760 41600
rect 150600 41600 150760 41760
rect 150600 41760 150760 41920
rect 150600 41920 150760 42080
rect 150600 42080 150760 42240
rect 150600 42240 150760 42400
rect 150600 42400 150760 42560
rect 150600 42560 150760 42720
rect 150600 42720 150760 42880
rect 150600 42880 150760 43040
rect 150600 43040 150760 43200
rect 150600 43200 150760 43360
rect 150600 43360 150760 43520
rect 150600 43520 150760 43680
rect 150600 43680 150760 43840
rect 150600 43840 150760 44000
rect 150600 44000 150760 44160
rect 150600 44160 150760 44320
rect 150600 44320 150760 44480
rect 150600 44480 150760 44640
rect 150600 44640 150760 44800
rect 150600 44800 150760 44960
rect 150600 44960 150760 45120
rect 150600 45120 150760 45280
rect 150600 45280 150760 45440
rect 150600 45440 150760 45600
rect 150600 45600 150760 45760
rect 150600 45760 150760 45920
rect 150600 45920 150760 46080
rect 150600 46080 150760 46240
rect 150600 46240 150760 46400
rect 150600 46400 150760 46560
rect 150600 46560 150760 46720
rect 150600 46720 150760 46880
rect 150600 46880 150760 47040
rect 150600 47040 150760 47200
rect 150600 47200 150760 47360
rect 150600 47360 150760 47520
rect 150600 47520 150760 47680
rect 150600 47680 150760 47840
rect 150600 47840 150760 48000
rect 150600 48000 150760 48160
rect 150600 48160 150760 48320
rect 150600 48320 150760 48480
rect 150600 48480 150760 48640
rect 150600 48640 150760 48800
rect 150600 48800 150760 48960
rect 150600 48960 150760 49120
rect 150600 49120 150760 49280
rect 150600 49280 150760 49440
rect 150600 49440 150760 49600
rect 150600 49600 150760 49760
rect 150600 49760 150760 49920
rect 150600 49920 150760 50080
rect 150600 50080 150760 50240
rect 150600 50240 150760 50400
rect 150600 50400 150760 50560
rect 150600 50560 150760 50720
rect 150600 50720 150760 50880
rect 150600 50880 150760 51040
rect 150600 51040 150760 51200
rect 150600 51200 150760 51360
rect 150600 51360 150760 51520
rect 150600 51520 150760 51680
rect 150600 51680 150760 51840
rect 150600 51840 150760 52000
rect 150600 52000 150760 52160
rect 150600 52160 150760 52320
rect 150600 52320 150760 52480
rect 150600 52480 150760 52640
rect 150600 52640 150760 52800
rect 150600 52800 150760 52960
rect 150600 52960 150760 53120
rect 150760 25920 150920 26080
rect 150760 26080 150920 26240
rect 150760 26240 150920 26400
rect 150760 26400 150920 26560
rect 150760 26560 150920 26720
rect 150760 26720 150920 26880
rect 150760 26880 150920 27040
rect 150760 27040 150920 27200
rect 150760 27200 150920 27360
rect 150760 27360 150920 27520
rect 150760 27520 150920 27680
rect 150760 27680 150920 27840
rect 150760 27840 150920 28000
rect 150760 28000 150920 28160
rect 150760 28160 150920 28320
rect 150760 28320 150920 28480
rect 150760 28480 150920 28640
rect 150760 28640 150920 28800
rect 150760 28800 150920 28960
rect 150760 28960 150920 29120
rect 150760 29120 150920 29280
rect 150760 29280 150920 29440
rect 150760 29440 150920 29600
rect 150760 29600 150920 29760
rect 150760 29760 150920 29920
rect 150760 29920 150920 30080
rect 150760 30080 150920 30240
rect 150760 30240 150920 30400
rect 150760 30400 150920 30560
rect 150760 30560 150920 30720
rect 150760 30720 150920 30880
rect 150760 30880 150920 31040
rect 150760 31040 150920 31200
rect 150760 31200 150920 31360
rect 150760 31360 150920 31520
rect 150760 31520 150920 31680
rect 150760 31680 150920 31840
rect 150760 31840 150920 32000
rect 150760 32000 150920 32160
rect 150760 32160 150920 32320
rect 150760 32320 150920 32480
rect 150760 32480 150920 32640
rect 150760 32640 150920 32800
rect 150760 32800 150920 32960
rect 150760 32960 150920 33120
rect 150760 33120 150920 33280
rect 150760 33280 150920 33440
rect 150760 33440 150920 33600
rect 150760 33600 150920 33760
rect 150760 33760 150920 33920
rect 150760 33920 150920 34080
rect 150760 34080 150920 34240
rect 150760 34240 150920 34400
rect 150760 34400 150920 34560
rect 150760 34560 150920 34720
rect 150760 34720 150920 34880
rect 150760 34880 150920 35040
rect 150760 35040 150920 35200
rect 150760 35200 150920 35360
rect 150760 35360 150920 35520
rect 150760 35520 150920 35680
rect 150760 35680 150920 35840
rect 150760 35840 150920 36000
rect 150760 36000 150920 36160
rect 150760 36160 150920 36320
rect 150760 36320 150920 36480
rect 150760 36480 150920 36640
rect 150760 36640 150920 36800
rect 150760 36800 150920 36960
rect 150760 36960 150920 37120
rect 150760 37120 150920 37280
rect 150760 37280 150920 37440
rect 150760 37440 150920 37600
rect 150760 37600 150920 37760
rect 150760 37760 150920 37920
rect 150760 37920 150920 38080
rect 150760 38080 150920 38240
rect 150760 38240 150920 38400
rect 150760 38400 150920 38560
rect 150760 38560 150920 38720
rect 150760 38720 150920 38880
rect 150760 38880 150920 39040
rect 150760 39040 150920 39200
rect 150760 39200 150920 39360
rect 150760 39360 150920 39520
rect 150760 39520 150920 39680
rect 150760 39680 150920 39840
rect 150760 39840 150920 40000
rect 150760 40000 150920 40160
rect 150760 40160 150920 40320
rect 150760 40320 150920 40480
rect 150760 40480 150920 40640
rect 150760 40640 150920 40800
rect 150760 40800 150920 40960
rect 150760 40960 150920 41120
rect 150760 41120 150920 41280
rect 150760 41280 150920 41440
rect 150760 41440 150920 41600
rect 150760 41600 150920 41760
rect 150760 41760 150920 41920
rect 150760 41920 150920 42080
rect 150760 42080 150920 42240
rect 150760 42240 150920 42400
rect 150760 42400 150920 42560
rect 150760 42560 150920 42720
rect 150760 42720 150920 42880
rect 150760 42880 150920 43040
rect 150760 43040 150920 43200
rect 150760 43200 150920 43360
rect 150760 43360 150920 43520
rect 150760 43520 150920 43680
rect 150760 43680 150920 43840
rect 150760 43840 150920 44000
rect 150760 44000 150920 44160
rect 150760 44160 150920 44320
rect 150760 44320 150920 44480
rect 150760 44480 150920 44640
rect 150760 44640 150920 44800
rect 150760 44800 150920 44960
rect 150760 44960 150920 45120
rect 150760 45120 150920 45280
rect 150760 45280 150920 45440
rect 150760 45440 150920 45600
rect 150760 45600 150920 45760
rect 150760 45760 150920 45920
rect 150760 45920 150920 46080
rect 150760 46080 150920 46240
rect 150760 46240 150920 46400
rect 150760 46400 150920 46560
rect 150760 46560 150920 46720
rect 150760 46720 150920 46880
rect 150760 46880 150920 47040
rect 150760 47040 150920 47200
rect 150760 47200 150920 47360
rect 150760 47360 150920 47520
rect 150760 47520 150920 47680
rect 150760 47680 150920 47840
rect 150760 47840 150920 48000
rect 150760 48000 150920 48160
rect 150760 48160 150920 48320
rect 150760 48320 150920 48480
rect 150760 48480 150920 48640
rect 150760 48640 150920 48800
rect 150760 48800 150920 48960
rect 150760 48960 150920 49120
rect 150760 49120 150920 49280
rect 150760 49280 150920 49440
rect 150760 49440 150920 49600
rect 150760 49600 150920 49760
rect 150760 49760 150920 49920
rect 150760 49920 150920 50080
rect 150760 50080 150920 50240
rect 150760 50240 150920 50400
rect 150760 50400 150920 50560
rect 150760 50560 150920 50720
rect 150760 50720 150920 50880
rect 150760 50880 150920 51040
rect 150760 51040 150920 51200
rect 150760 51200 150920 51360
rect 150760 51360 150920 51520
rect 150760 51520 150920 51680
rect 150760 51680 150920 51840
rect 150760 51840 150920 52000
rect 150760 52000 150920 52160
rect 150760 52160 150920 52320
rect 150760 52320 150920 52480
rect 150760 52480 150920 52640
rect 150760 52640 150920 52800
rect 150760 52800 150920 52960
rect 150760 52960 150920 53120
rect 150760 53120 150920 53280
rect 150920 25920 151080 26080
rect 150920 26080 151080 26240
rect 150920 26240 151080 26400
rect 150920 26400 151080 26560
rect 150920 26560 151080 26720
rect 150920 26720 151080 26880
rect 150920 26880 151080 27040
rect 150920 27040 151080 27200
rect 150920 27200 151080 27360
rect 150920 27360 151080 27520
rect 150920 27520 151080 27680
rect 150920 27680 151080 27840
rect 150920 27840 151080 28000
rect 150920 28000 151080 28160
rect 150920 28160 151080 28320
rect 150920 28320 151080 28480
rect 150920 28480 151080 28640
rect 150920 28640 151080 28800
rect 150920 28800 151080 28960
rect 150920 28960 151080 29120
rect 150920 29120 151080 29280
rect 150920 29280 151080 29440
rect 150920 29440 151080 29600
rect 150920 29600 151080 29760
rect 150920 29760 151080 29920
rect 150920 29920 151080 30080
rect 150920 30080 151080 30240
rect 150920 30240 151080 30400
rect 150920 30400 151080 30560
rect 150920 30560 151080 30720
rect 150920 30720 151080 30880
rect 150920 30880 151080 31040
rect 150920 31040 151080 31200
rect 150920 31200 151080 31360
rect 150920 31360 151080 31520
rect 150920 31520 151080 31680
rect 150920 31680 151080 31840
rect 150920 31840 151080 32000
rect 150920 32000 151080 32160
rect 150920 32160 151080 32320
rect 150920 32320 151080 32480
rect 150920 32480 151080 32640
rect 150920 32640 151080 32800
rect 150920 32800 151080 32960
rect 150920 32960 151080 33120
rect 150920 33120 151080 33280
rect 150920 33280 151080 33440
rect 150920 33440 151080 33600
rect 150920 33600 151080 33760
rect 150920 33760 151080 33920
rect 150920 33920 151080 34080
rect 150920 34080 151080 34240
rect 150920 34240 151080 34400
rect 150920 34400 151080 34560
rect 150920 34560 151080 34720
rect 150920 34720 151080 34880
rect 150920 34880 151080 35040
rect 150920 35040 151080 35200
rect 150920 35200 151080 35360
rect 150920 35360 151080 35520
rect 150920 35520 151080 35680
rect 150920 35680 151080 35840
rect 150920 35840 151080 36000
rect 150920 36000 151080 36160
rect 150920 36160 151080 36320
rect 150920 36320 151080 36480
rect 150920 36480 151080 36640
rect 150920 36640 151080 36800
rect 150920 36800 151080 36960
rect 150920 36960 151080 37120
rect 150920 37120 151080 37280
rect 150920 37280 151080 37440
rect 150920 37440 151080 37600
rect 150920 37600 151080 37760
rect 150920 37760 151080 37920
rect 150920 37920 151080 38080
rect 150920 38080 151080 38240
rect 150920 38240 151080 38400
rect 150920 38400 151080 38560
rect 150920 38560 151080 38720
rect 150920 38720 151080 38880
rect 150920 38880 151080 39040
rect 150920 39040 151080 39200
rect 150920 39200 151080 39360
rect 150920 39360 151080 39520
rect 150920 39520 151080 39680
rect 150920 39680 151080 39840
rect 150920 39840 151080 40000
rect 150920 40000 151080 40160
rect 150920 40160 151080 40320
rect 150920 40320 151080 40480
rect 150920 40480 151080 40640
rect 150920 40640 151080 40800
rect 150920 40800 151080 40960
rect 150920 40960 151080 41120
rect 150920 41120 151080 41280
rect 150920 41280 151080 41440
rect 150920 41440 151080 41600
rect 150920 41600 151080 41760
rect 150920 41760 151080 41920
rect 150920 41920 151080 42080
rect 150920 42080 151080 42240
rect 150920 42240 151080 42400
rect 150920 42400 151080 42560
rect 150920 42560 151080 42720
rect 150920 42720 151080 42880
rect 150920 42880 151080 43040
rect 150920 43040 151080 43200
rect 150920 43200 151080 43360
rect 150920 43360 151080 43520
rect 150920 43520 151080 43680
rect 150920 43680 151080 43840
rect 150920 43840 151080 44000
rect 150920 44000 151080 44160
rect 150920 44160 151080 44320
rect 150920 44320 151080 44480
rect 150920 44480 151080 44640
rect 150920 44640 151080 44800
rect 150920 44800 151080 44960
rect 150920 44960 151080 45120
rect 150920 45120 151080 45280
rect 150920 45280 151080 45440
rect 150920 45440 151080 45600
rect 150920 45600 151080 45760
rect 150920 45760 151080 45920
rect 150920 45920 151080 46080
rect 150920 46080 151080 46240
rect 150920 46240 151080 46400
rect 150920 46400 151080 46560
rect 150920 46560 151080 46720
rect 150920 46720 151080 46880
rect 150920 46880 151080 47040
rect 150920 47040 151080 47200
rect 150920 47200 151080 47360
rect 150920 47360 151080 47520
rect 150920 47520 151080 47680
rect 150920 47680 151080 47840
rect 150920 47840 151080 48000
rect 150920 48000 151080 48160
rect 150920 48160 151080 48320
rect 150920 48320 151080 48480
rect 150920 48480 151080 48640
rect 150920 48640 151080 48800
rect 150920 48800 151080 48960
rect 150920 48960 151080 49120
rect 150920 49120 151080 49280
rect 150920 49280 151080 49440
rect 150920 49440 151080 49600
rect 150920 49600 151080 49760
rect 150920 49760 151080 49920
rect 150920 49920 151080 50080
rect 150920 50080 151080 50240
rect 150920 50240 151080 50400
rect 150920 50400 151080 50560
rect 150920 50560 151080 50720
rect 150920 50720 151080 50880
rect 150920 50880 151080 51040
rect 150920 51040 151080 51200
rect 150920 51200 151080 51360
rect 150920 51360 151080 51520
rect 150920 51520 151080 51680
rect 150920 51680 151080 51840
rect 150920 51840 151080 52000
rect 150920 52000 151080 52160
rect 150920 52160 151080 52320
rect 150920 52320 151080 52480
rect 150920 52480 151080 52640
rect 150920 52640 151080 52800
rect 150920 52800 151080 52960
rect 150920 52960 151080 53120
rect 150920 53120 151080 53280
rect 151080 25760 151240 25920
rect 151080 25920 151240 26080
rect 151080 26080 151240 26240
rect 151080 26240 151240 26400
rect 151080 26400 151240 26560
rect 151080 26560 151240 26720
rect 151080 26720 151240 26880
rect 151080 26880 151240 27040
rect 151080 27040 151240 27200
rect 151080 27200 151240 27360
rect 151080 27360 151240 27520
rect 151080 27520 151240 27680
rect 151080 27680 151240 27840
rect 151080 27840 151240 28000
rect 151080 28000 151240 28160
rect 151080 28160 151240 28320
rect 151080 28320 151240 28480
rect 151080 28480 151240 28640
rect 151080 28640 151240 28800
rect 151080 28800 151240 28960
rect 151080 28960 151240 29120
rect 151080 29120 151240 29280
rect 151080 29280 151240 29440
rect 151080 29440 151240 29600
rect 151080 29600 151240 29760
rect 151080 29760 151240 29920
rect 151080 29920 151240 30080
rect 151080 30080 151240 30240
rect 151080 30240 151240 30400
rect 151080 30400 151240 30560
rect 151080 30560 151240 30720
rect 151080 30720 151240 30880
rect 151080 30880 151240 31040
rect 151080 31040 151240 31200
rect 151080 31200 151240 31360
rect 151080 31360 151240 31520
rect 151080 31520 151240 31680
rect 151080 31680 151240 31840
rect 151080 31840 151240 32000
rect 151080 32000 151240 32160
rect 151080 32160 151240 32320
rect 151080 32320 151240 32480
rect 151080 32480 151240 32640
rect 151080 32640 151240 32800
rect 151080 32800 151240 32960
rect 151080 32960 151240 33120
rect 151080 33120 151240 33280
rect 151080 33280 151240 33440
rect 151080 33440 151240 33600
rect 151080 33600 151240 33760
rect 151080 33760 151240 33920
rect 151080 33920 151240 34080
rect 151080 34080 151240 34240
rect 151080 34240 151240 34400
rect 151080 34400 151240 34560
rect 151080 34560 151240 34720
rect 151080 34720 151240 34880
rect 151080 34880 151240 35040
rect 151080 35040 151240 35200
rect 151080 35200 151240 35360
rect 151080 35360 151240 35520
rect 151080 35520 151240 35680
rect 151080 35680 151240 35840
rect 151080 35840 151240 36000
rect 151080 36000 151240 36160
rect 151080 36160 151240 36320
rect 151080 36320 151240 36480
rect 151080 36480 151240 36640
rect 151080 36640 151240 36800
rect 151080 36800 151240 36960
rect 151080 36960 151240 37120
rect 151080 37120 151240 37280
rect 151080 37280 151240 37440
rect 151080 37440 151240 37600
rect 151080 37600 151240 37760
rect 151080 37760 151240 37920
rect 151080 37920 151240 38080
rect 151080 38080 151240 38240
rect 151080 38240 151240 38400
rect 151080 38400 151240 38560
rect 151080 38560 151240 38720
rect 151080 38720 151240 38880
rect 151080 38880 151240 39040
rect 151080 39040 151240 39200
rect 151080 39200 151240 39360
rect 151080 39360 151240 39520
rect 151080 39520 151240 39680
rect 151080 39680 151240 39840
rect 151080 39840 151240 40000
rect 151080 40000 151240 40160
rect 151080 40160 151240 40320
rect 151080 40320 151240 40480
rect 151080 40480 151240 40640
rect 151080 40640 151240 40800
rect 151080 40800 151240 40960
rect 151080 40960 151240 41120
rect 151080 41120 151240 41280
rect 151080 41280 151240 41440
rect 151080 41440 151240 41600
rect 151080 41600 151240 41760
rect 151080 41760 151240 41920
rect 151080 41920 151240 42080
rect 151080 42080 151240 42240
rect 151080 42240 151240 42400
rect 151080 42400 151240 42560
rect 151080 42560 151240 42720
rect 151080 42720 151240 42880
rect 151080 42880 151240 43040
rect 151080 43040 151240 43200
rect 151080 43200 151240 43360
rect 151080 43360 151240 43520
rect 151080 43520 151240 43680
rect 151080 43680 151240 43840
rect 151080 43840 151240 44000
rect 151080 44000 151240 44160
rect 151080 44160 151240 44320
rect 151080 44320 151240 44480
rect 151080 44480 151240 44640
rect 151080 44640 151240 44800
rect 151080 44800 151240 44960
rect 151080 44960 151240 45120
rect 151080 45120 151240 45280
rect 151080 45280 151240 45440
rect 151080 45440 151240 45600
rect 151080 45600 151240 45760
rect 151080 45760 151240 45920
rect 151080 45920 151240 46080
rect 151080 46080 151240 46240
rect 151080 46240 151240 46400
rect 151080 46400 151240 46560
rect 151080 46560 151240 46720
rect 151080 46720 151240 46880
rect 151080 46880 151240 47040
rect 151080 47040 151240 47200
rect 151080 47200 151240 47360
rect 151080 47360 151240 47520
rect 151080 47520 151240 47680
rect 151080 47680 151240 47840
rect 151080 47840 151240 48000
rect 151080 48000 151240 48160
rect 151080 48160 151240 48320
rect 151080 48320 151240 48480
rect 151080 48480 151240 48640
rect 151080 48640 151240 48800
rect 151080 48800 151240 48960
rect 151080 48960 151240 49120
rect 151080 49120 151240 49280
rect 151080 49280 151240 49440
rect 151080 49440 151240 49600
rect 151080 49600 151240 49760
rect 151080 49760 151240 49920
rect 151080 49920 151240 50080
rect 151080 50080 151240 50240
rect 151080 50240 151240 50400
rect 151080 50400 151240 50560
rect 151080 50560 151240 50720
rect 151080 50720 151240 50880
rect 151080 50880 151240 51040
rect 151080 51040 151240 51200
rect 151080 51200 151240 51360
rect 151080 51360 151240 51520
rect 151080 51520 151240 51680
rect 151080 51680 151240 51840
rect 151080 51840 151240 52000
rect 151080 52000 151240 52160
rect 151080 52160 151240 52320
rect 151080 52320 151240 52480
rect 151080 52480 151240 52640
rect 151080 52640 151240 52800
rect 151080 52800 151240 52960
rect 151080 52960 151240 53120
rect 151080 53120 151240 53280
rect 151240 25760 151400 25920
rect 151240 25920 151400 26080
rect 151240 26080 151400 26240
rect 151240 26240 151400 26400
rect 151240 26400 151400 26560
rect 151240 26560 151400 26720
rect 151240 26720 151400 26880
rect 151240 26880 151400 27040
rect 151240 27040 151400 27200
rect 151240 27200 151400 27360
rect 151240 27360 151400 27520
rect 151240 27520 151400 27680
rect 151240 27680 151400 27840
rect 151240 27840 151400 28000
rect 151240 28000 151400 28160
rect 151240 28160 151400 28320
rect 151240 28320 151400 28480
rect 151240 28480 151400 28640
rect 151240 28640 151400 28800
rect 151240 28800 151400 28960
rect 151240 28960 151400 29120
rect 151240 29120 151400 29280
rect 151240 29280 151400 29440
rect 151240 29440 151400 29600
rect 151240 29600 151400 29760
rect 151240 29760 151400 29920
rect 151240 29920 151400 30080
rect 151240 30080 151400 30240
rect 151240 30240 151400 30400
rect 151240 30400 151400 30560
rect 151240 30560 151400 30720
rect 151240 30720 151400 30880
rect 151240 30880 151400 31040
rect 151240 31040 151400 31200
rect 151240 31200 151400 31360
rect 151240 31360 151400 31520
rect 151240 31520 151400 31680
rect 151240 31680 151400 31840
rect 151240 31840 151400 32000
rect 151240 32000 151400 32160
rect 151240 32160 151400 32320
rect 151240 32320 151400 32480
rect 151240 32480 151400 32640
rect 151240 32640 151400 32800
rect 151240 32800 151400 32960
rect 151240 32960 151400 33120
rect 151240 33120 151400 33280
rect 151240 33280 151400 33440
rect 151240 33440 151400 33600
rect 151240 33600 151400 33760
rect 151240 33760 151400 33920
rect 151240 33920 151400 34080
rect 151240 34080 151400 34240
rect 151240 34240 151400 34400
rect 151240 34400 151400 34560
rect 151240 34560 151400 34720
rect 151240 34720 151400 34880
rect 151240 34880 151400 35040
rect 151240 35040 151400 35200
rect 151240 35200 151400 35360
rect 151240 35360 151400 35520
rect 151240 35520 151400 35680
rect 151240 35680 151400 35840
rect 151240 35840 151400 36000
rect 151240 36000 151400 36160
rect 151240 36160 151400 36320
rect 151240 36320 151400 36480
rect 151240 36480 151400 36640
rect 151240 36640 151400 36800
rect 151240 36800 151400 36960
rect 151240 36960 151400 37120
rect 151240 37120 151400 37280
rect 151240 37280 151400 37440
rect 151240 37440 151400 37600
rect 151240 37600 151400 37760
rect 151240 37760 151400 37920
rect 151240 37920 151400 38080
rect 151240 38080 151400 38240
rect 151240 38240 151400 38400
rect 151240 38400 151400 38560
rect 151240 38560 151400 38720
rect 151240 38720 151400 38880
rect 151240 38880 151400 39040
rect 151240 39040 151400 39200
rect 151240 39200 151400 39360
rect 151240 39360 151400 39520
rect 151240 39520 151400 39680
rect 151240 39680 151400 39840
rect 151240 39840 151400 40000
rect 151240 40000 151400 40160
rect 151240 40160 151400 40320
rect 151240 40320 151400 40480
rect 151240 40480 151400 40640
rect 151240 40640 151400 40800
rect 151240 40800 151400 40960
rect 151240 40960 151400 41120
rect 151240 41120 151400 41280
rect 151240 41280 151400 41440
rect 151240 41440 151400 41600
rect 151240 41600 151400 41760
rect 151240 41760 151400 41920
rect 151240 41920 151400 42080
rect 151240 42080 151400 42240
rect 151240 42240 151400 42400
rect 151240 42400 151400 42560
rect 151240 42560 151400 42720
rect 151240 42720 151400 42880
rect 151240 42880 151400 43040
rect 151240 43040 151400 43200
rect 151240 43200 151400 43360
rect 151240 43360 151400 43520
rect 151240 43520 151400 43680
rect 151240 43680 151400 43840
rect 151240 43840 151400 44000
rect 151240 44000 151400 44160
rect 151240 44160 151400 44320
rect 151240 44320 151400 44480
rect 151240 44480 151400 44640
rect 151240 44640 151400 44800
rect 151240 44800 151400 44960
rect 151240 44960 151400 45120
rect 151240 45120 151400 45280
rect 151240 45280 151400 45440
rect 151240 45440 151400 45600
rect 151240 45600 151400 45760
rect 151240 45760 151400 45920
rect 151240 45920 151400 46080
rect 151240 46080 151400 46240
rect 151240 46240 151400 46400
rect 151240 46400 151400 46560
rect 151240 46560 151400 46720
rect 151240 46720 151400 46880
rect 151240 46880 151400 47040
rect 151240 47040 151400 47200
rect 151240 47200 151400 47360
rect 151240 47360 151400 47520
rect 151240 47520 151400 47680
rect 151240 47680 151400 47840
rect 151240 47840 151400 48000
rect 151240 48000 151400 48160
rect 151240 48160 151400 48320
rect 151240 48320 151400 48480
rect 151240 48480 151400 48640
rect 151240 48640 151400 48800
rect 151240 48800 151400 48960
rect 151240 48960 151400 49120
rect 151240 49120 151400 49280
rect 151240 49280 151400 49440
rect 151240 49440 151400 49600
rect 151240 49600 151400 49760
rect 151240 49760 151400 49920
rect 151240 49920 151400 50080
rect 151240 50080 151400 50240
rect 151240 50240 151400 50400
rect 151240 50400 151400 50560
rect 151240 50560 151400 50720
rect 151240 50720 151400 50880
rect 151240 50880 151400 51040
rect 151240 51040 151400 51200
rect 151240 51200 151400 51360
rect 151240 51360 151400 51520
rect 151240 51520 151400 51680
rect 151240 51680 151400 51840
rect 151240 51840 151400 52000
rect 151240 52000 151400 52160
rect 151240 52160 151400 52320
rect 151240 52320 151400 52480
rect 151240 52480 151400 52640
rect 151240 52640 151400 52800
rect 151240 52800 151400 52960
rect 151240 52960 151400 53120
rect 151240 53120 151400 53280
rect 151400 25760 151560 25920
rect 151400 25920 151560 26080
rect 151400 26080 151560 26240
rect 151400 26240 151560 26400
rect 151400 26400 151560 26560
rect 151400 26560 151560 26720
rect 151400 26720 151560 26880
rect 151400 26880 151560 27040
rect 151400 27040 151560 27200
rect 151400 27200 151560 27360
rect 151400 27360 151560 27520
rect 151400 27520 151560 27680
rect 151400 27680 151560 27840
rect 151400 27840 151560 28000
rect 151400 28000 151560 28160
rect 151400 28160 151560 28320
rect 151400 28320 151560 28480
rect 151400 28480 151560 28640
rect 151400 28640 151560 28800
rect 151400 28800 151560 28960
rect 151400 28960 151560 29120
rect 151400 29120 151560 29280
rect 151400 29280 151560 29440
rect 151400 29440 151560 29600
rect 151400 29600 151560 29760
rect 151400 29760 151560 29920
rect 151400 29920 151560 30080
rect 151400 30080 151560 30240
rect 151400 30240 151560 30400
rect 151400 30400 151560 30560
rect 151400 30560 151560 30720
rect 151400 30720 151560 30880
rect 151400 30880 151560 31040
rect 151400 31040 151560 31200
rect 151400 31200 151560 31360
rect 151400 31360 151560 31520
rect 151400 31520 151560 31680
rect 151400 31680 151560 31840
rect 151400 31840 151560 32000
rect 151400 32000 151560 32160
rect 151400 32160 151560 32320
rect 151400 32320 151560 32480
rect 151400 32480 151560 32640
rect 151400 32640 151560 32800
rect 151400 32800 151560 32960
rect 151400 32960 151560 33120
rect 151400 33120 151560 33280
rect 151400 33280 151560 33440
rect 151400 33440 151560 33600
rect 151400 33600 151560 33760
rect 151400 33760 151560 33920
rect 151400 33920 151560 34080
rect 151400 34080 151560 34240
rect 151400 34240 151560 34400
rect 151400 34400 151560 34560
rect 151400 34560 151560 34720
rect 151400 34720 151560 34880
rect 151400 34880 151560 35040
rect 151400 35040 151560 35200
rect 151400 35200 151560 35360
rect 151400 35360 151560 35520
rect 151400 35520 151560 35680
rect 151400 35680 151560 35840
rect 151400 35840 151560 36000
rect 151400 36000 151560 36160
rect 151400 36160 151560 36320
rect 151400 36320 151560 36480
rect 151400 36480 151560 36640
rect 151400 36640 151560 36800
rect 151400 36800 151560 36960
rect 151400 36960 151560 37120
rect 151400 37120 151560 37280
rect 151400 37280 151560 37440
rect 151400 37440 151560 37600
rect 151400 37600 151560 37760
rect 151400 37760 151560 37920
rect 151400 37920 151560 38080
rect 151400 38080 151560 38240
rect 151400 38240 151560 38400
rect 151400 38400 151560 38560
rect 151400 38560 151560 38720
rect 151400 38720 151560 38880
rect 151400 38880 151560 39040
rect 151400 39040 151560 39200
rect 151400 39840 151560 40000
rect 151400 40000 151560 40160
rect 151400 40160 151560 40320
rect 151400 40320 151560 40480
rect 151400 40480 151560 40640
rect 151400 40640 151560 40800
rect 151400 40800 151560 40960
rect 151400 40960 151560 41120
rect 151400 41120 151560 41280
rect 151400 41280 151560 41440
rect 151400 41440 151560 41600
rect 151400 41600 151560 41760
rect 151400 41760 151560 41920
rect 151400 41920 151560 42080
rect 151400 42080 151560 42240
rect 151400 42240 151560 42400
rect 151400 42400 151560 42560
rect 151400 42560 151560 42720
rect 151400 42720 151560 42880
rect 151400 42880 151560 43040
rect 151400 43040 151560 43200
rect 151400 43200 151560 43360
rect 151400 43360 151560 43520
rect 151400 43520 151560 43680
rect 151400 43680 151560 43840
rect 151400 43840 151560 44000
rect 151400 44000 151560 44160
rect 151400 44160 151560 44320
rect 151400 44320 151560 44480
rect 151400 44480 151560 44640
rect 151400 44640 151560 44800
rect 151400 44800 151560 44960
rect 151400 44960 151560 45120
rect 151400 45120 151560 45280
rect 151400 45280 151560 45440
rect 151400 45440 151560 45600
rect 151400 45600 151560 45760
rect 151400 45760 151560 45920
rect 151400 45920 151560 46080
rect 151400 46080 151560 46240
rect 151400 46240 151560 46400
rect 151400 46400 151560 46560
rect 151400 46560 151560 46720
rect 151400 46720 151560 46880
rect 151400 46880 151560 47040
rect 151400 47040 151560 47200
rect 151400 47200 151560 47360
rect 151400 47360 151560 47520
rect 151400 47520 151560 47680
rect 151400 47680 151560 47840
rect 151400 47840 151560 48000
rect 151400 48000 151560 48160
rect 151400 48160 151560 48320
rect 151400 48320 151560 48480
rect 151400 48480 151560 48640
rect 151400 48640 151560 48800
rect 151400 48800 151560 48960
rect 151400 48960 151560 49120
rect 151400 49120 151560 49280
rect 151400 49280 151560 49440
rect 151400 49440 151560 49600
rect 151400 49600 151560 49760
rect 151400 49760 151560 49920
rect 151400 49920 151560 50080
rect 151400 50080 151560 50240
rect 151400 50240 151560 50400
rect 151400 50400 151560 50560
rect 151400 50560 151560 50720
rect 151400 50720 151560 50880
rect 151400 50880 151560 51040
rect 151400 51040 151560 51200
rect 151400 51200 151560 51360
rect 151400 51360 151560 51520
rect 151400 51520 151560 51680
rect 151400 51680 151560 51840
rect 151400 51840 151560 52000
rect 151400 52000 151560 52160
rect 151400 52160 151560 52320
rect 151400 52320 151560 52480
rect 151400 52480 151560 52640
rect 151400 52640 151560 52800
rect 151400 52800 151560 52960
rect 151400 52960 151560 53120
rect 151400 53120 151560 53280
rect 151400 53280 151560 53440
rect 151560 25920 151720 26080
rect 151560 26080 151720 26240
rect 151560 26240 151720 26400
rect 151560 26400 151720 26560
rect 151560 26560 151720 26720
rect 151560 26720 151720 26880
rect 151560 26880 151720 27040
rect 151560 27040 151720 27200
rect 151560 27200 151720 27360
rect 151560 27360 151720 27520
rect 151560 27520 151720 27680
rect 151560 27680 151720 27840
rect 151560 27840 151720 28000
rect 151560 28000 151720 28160
rect 151560 28160 151720 28320
rect 151560 28320 151720 28480
rect 151560 28480 151720 28640
rect 151560 28640 151720 28800
rect 151560 28800 151720 28960
rect 151560 28960 151720 29120
rect 151560 29120 151720 29280
rect 151560 29280 151720 29440
rect 151560 29440 151720 29600
rect 151560 29600 151720 29760
rect 151560 29760 151720 29920
rect 151560 29920 151720 30080
rect 151560 30080 151720 30240
rect 151560 30240 151720 30400
rect 151560 30400 151720 30560
rect 151560 30560 151720 30720
rect 151560 30720 151720 30880
rect 151560 30880 151720 31040
rect 151560 31040 151720 31200
rect 151560 31200 151720 31360
rect 151560 31360 151720 31520
rect 151560 31520 151720 31680
rect 151560 31680 151720 31840
rect 151560 31840 151720 32000
rect 151560 32000 151720 32160
rect 151560 32160 151720 32320
rect 151560 32320 151720 32480
rect 151560 32480 151720 32640
rect 151560 32640 151720 32800
rect 151560 32800 151720 32960
rect 151560 32960 151720 33120
rect 151560 33120 151720 33280
rect 151560 33280 151720 33440
rect 151560 33440 151720 33600
rect 151560 33600 151720 33760
rect 151560 33760 151720 33920
rect 151560 33920 151720 34080
rect 151560 34080 151720 34240
rect 151560 34240 151720 34400
rect 151560 34400 151720 34560
rect 151560 34560 151720 34720
rect 151560 34720 151720 34880
rect 151560 34880 151720 35040
rect 151560 35040 151720 35200
rect 151560 35200 151720 35360
rect 151560 35360 151720 35520
rect 151560 35520 151720 35680
rect 151560 35680 151720 35840
rect 151560 35840 151720 36000
rect 151560 36000 151720 36160
rect 151560 36160 151720 36320
rect 151560 36320 151720 36480
rect 151560 36480 151720 36640
rect 151560 36640 151720 36800
rect 151560 36800 151720 36960
rect 151560 36960 151720 37120
rect 151560 37120 151720 37280
rect 151560 37280 151720 37440
rect 151560 37440 151720 37600
rect 151560 37600 151720 37760
rect 151560 37760 151720 37920
rect 151560 37920 151720 38080
rect 151560 38080 151720 38240
rect 151560 38240 151720 38400
rect 151560 38400 151720 38560
rect 151560 38560 151720 38720
rect 151560 38720 151720 38880
rect 151560 40160 151720 40320
rect 151560 40320 151720 40480
rect 151560 40480 151720 40640
rect 151560 40640 151720 40800
rect 151560 40800 151720 40960
rect 151560 40960 151720 41120
rect 151560 41120 151720 41280
rect 151560 41280 151720 41440
rect 151560 41440 151720 41600
rect 151560 41600 151720 41760
rect 151560 41760 151720 41920
rect 151560 41920 151720 42080
rect 151560 42080 151720 42240
rect 151560 42240 151720 42400
rect 151560 42400 151720 42560
rect 151560 42560 151720 42720
rect 151560 42720 151720 42880
rect 151560 42880 151720 43040
rect 151560 43040 151720 43200
rect 151560 43200 151720 43360
rect 151560 43360 151720 43520
rect 151560 43520 151720 43680
rect 151560 43680 151720 43840
rect 151560 43840 151720 44000
rect 151560 44000 151720 44160
rect 151560 44160 151720 44320
rect 151560 44320 151720 44480
rect 151560 44480 151720 44640
rect 151560 44640 151720 44800
rect 151560 44800 151720 44960
rect 151560 44960 151720 45120
rect 151560 45120 151720 45280
rect 151560 45280 151720 45440
rect 151560 45440 151720 45600
rect 151560 45600 151720 45760
rect 151560 45760 151720 45920
rect 151560 45920 151720 46080
rect 151560 46080 151720 46240
rect 151560 46240 151720 46400
rect 151560 46400 151720 46560
rect 151560 46560 151720 46720
rect 151560 46720 151720 46880
rect 151560 46880 151720 47040
rect 151560 47040 151720 47200
rect 151560 47200 151720 47360
rect 151560 47360 151720 47520
rect 151560 47520 151720 47680
rect 151560 47680 151720 47840
rect 151560 47840 151720 48000
rect 151560 48000 151720 48160
rect 151560 48160 151720 48320
rect 151560 48320 151720 48480
rect 151560 48480 151720 48640
rect 151560 48640 151720 48800
rect 151560 48800 151720 48960
rect 151560 48960 151720 49120
rect 151560 49120 151720 49280
rect 151560 49280 151720 49440
rect 151560 49440 151720 49600
rect 151560 49600 151720 49760
rect 151560 49760 151720 49920
rect 151560 49920 151720 50080
rect 151560 50080 151720 50240
rect 151560 50240 151720 50400
rect 151560 50400 151720 50560
rect 151560 50560 151720 50720
rect 151560 50720 151720 50880
rect 151560 50880 151720 51040
rect 151560 51040 151720 51200
rect 151560 51200 151720 51360
rect 151560 51360 151720 51520
rect 151560 51520 151720 51680
rect 151560 51680 151720 51840
rect 151560 51840 151720 52000
rect 151560 52000 151720 52160
rect 151560 52160 151720 52320
rect 151560 52320 151720 52480
rect 151560 52480 151720 52640
rect 151560 52640 151720 52800
rect 151560 52800 151720 52960
rect 151560 52960 151720 53120
rect 151560 53120 151720 53280
rect 151720 25920 151880 26080
rect 151720 26080 151880 26240
rect 151720 26240 151880 26400
rect 151720 26400 151880 26560
rect 151720 26560 151880 26720
rect 151720 26720 151880 26880
rect 151720 26880 151880 27040
rect 151720 27040 151880 27200
rect 151720 27200 151880 27360
rect 151720 27360 151880 27520
rect 151720 27520 151880 27680
rect 151720 27680 151880 27840
rect 151720 27840 151880 28000
rect 151720 28000 151880 28160
rect 151720 28160 151880 28320
rect 151720 28320 151880 28480
rect 151720 28480 151880 28640
rect 151720 28640 151880 28800
rect 151720 28800 151880 28960
rect 151720 28960 151880 29120
rect 151720 29120 151880 29280
rect 151720 29280 151880 29440
rect 151720 29440 151880 29600
rect 151720 29600 151880 29760
rect 151720 29760 151880 29920
rect 151720 29920 151880 30080
rect 151720 30080 151880 30240
rect 151720 30240 151880 30400
rect 151720 30400 151880 30560
rect 151720 30560 151880 30720
rect 151720 30720 151880 30880
rect 151720 30880 151880 31040
rect 151720 31040 151880 31200
rect 151720 31200 151880 31360
rect 151720 31360 151880 31520
rect 151720 31520 151880 31680
rect 151720 31680 151880 31840
rect 151720 31840 151880 32000
rect 151720 32000 151880 32160
rect 151720 32160 151880 32320
rect 151720 32320 151880 32480
rect 151720 32480 151880 32640
rect 151720 32640 151880 32800
rect 151720 32800 151880 32960
rect 151720 32960 151880 33120
rect 151720 33120 151880 33280
rect 151720 33280 151880 33440
rect 151720 33440 151880 33600
rect 151720 33600 151880 33760
rect 151720 33760 151880 33920
rect 151720 33920 151880 34080
rect 151720 34080 151880 34240
rect 151720 34240 151880 34400
rect 151720 34400 151880 34560
rect 151720 34560 151880 34720
rect 151720 34720 151880 34880
rect 151720 34880 151880 35040
rect 151720 35040 151880 35200
rect 151720 35200 151880 35360
rect 151720 35360 151880 35520
rect 151720 35520 151880 35680
rect 151720 35680 151880 35840
rect 151720 35840 151880 36000
rect 151720 36000 151880 36160
rect 151720 36160 151880 36320
rect 151720 36320 151880 36480
rect 151720 36480 151880 36640
rect 151720 36640 151880 36800
rect 151720 36800 151880 36960
rect 151720 36960 151880 37120
rect 151720 37120 151880 37280
rect 151720 37280 151880 37440
rect 151720 37440 151880 37600
rect 151720 37600 151880 37760
rect 151720 37760 151880 37920
rect 151720 37920 151880 38080
rect 151720 38080 151880 38240
rect 151720 38240 151880 38400
rect 151720 38400 151880 38560
rect 151720 40480 151880 40640
rect 151720 40640 151880 40800
rect 151720 40800 151880 40960
rect 151720 40960 151880 41120
rect 151720 41120 151880 41280
rect 151720 41280 151880 41440
rect 151720 41440 151880 41600
rect 151720 41600 151880 41760
rect 151720 41760 151880 41920
rect 151720 41920 151880 42080
rect 151720 42080 151880 42240
rect 151720 42240 151880 42400
rect 151720 42400 151880 42560
rect 151720 42560 151880 42720
rect 151720 42720 151880 42880
rect 151720 42880 151880 43040
rect 151720 43040 151880 43200
rect 151720 43200 151880 43360
rect 151720 43360 151880 43520
rect 151720 43520 151880 43680
rect 151720 43680 151880 43840
rect 151720 43840 151880 44000
rect 151720 44000 151880 44160
rect 151720 44160 151880 44320
rect 151720 44320 151880 44480
rect 151720 44480 151880 44640
rect 151720 44640 151880 44800
rect 151720 44800 151880 44960
rect 151720 44960 151880 45120
rect 151720 45120 151880 45280
rect 151720 45280 151880 45440
rect 151720 45440 151880 45600
rect 151720 45600 151880 45760
rect 151720 45760 151880 45920
rect 151720 45920 151880 46080
rect 151720 46080 151880 46240
rect 151720 46240 151880 46400
rect 151720 46400 151880 46560
rect 151720 46560 151880 46720
rect 151720 46720 151880 46880
rect 151720 46880 151880 47040
rect 151720 47040 151880 47200
rect 151720 47200 151880 47360
rect 151720 47360 151880 47520
rect 151720 47520 151880 47680
rect 151720 47680 151880 47840
rect 151720 47840 151880 48000
rect 151720 48000 151880 48160
rect 151720 48160 151880 48320
rect 151720 48320 151880 48480
rect 151720 48480 151880 48640
rect 151720 48640 151880 48800
rect 151720 48800 151880 48960
rect 151720 48960 151880 49120
rect 151720 49120 151880 49280
rect 151720 49280 151880 49440
rect 151720 49440 151880 49600
rect 151720 49600 151880 49760
rect 151720 49760 151880 49920
rect 151720 49920 151880 50080
rect 151720 50080 151880 50240
rect 151720 50240 151880 50400
rect 151720 50400 151880 50560
rect 151720 50560 151880 50720
rect 151720 50720 151880 50880
rect 151720 50880 151880 51040
rect 151720 51040 151880 51200
rect 151720 51200 151880 51360
rect 151720 51360 151880 51520
rect 151720 51520 151880 51680
rect 151720 51680 151880 51840
rect 151720 51840 151880 52000
rect 151720 52000 151880 52160
rect 151720 52160 151880 52320
rect 151720 52320 151880 52480
rect 151720 52480 151880 52640
rect 151720 52640 151880 52800
rect 151720 52800 151880 52960
rect 151720 52960 151880 53120
rect 151720 53120 151880 53280
rect 151880 25920 152040 26080
rect 151880 26080 152040 26240
rect 151880 26240 152040 26400
rect 151880 26400 152040 26560
rect 151880 26560 152040 26720
rect 151880 26720 152040 26880
rect 151880 26880 152040 27040
rect 151880 27040 152040 27200
rect 151880 27200 152040 27360
rect 151880 27360 152040 27520
rect 151880 27520 152040 27680
rect 151880 27680 152040 27840
rect 151880 27840 152040 28000
rect 151880 28000 152040 28160
rect 151880 28160 152040 28320
rect 151880 28320 152040 28480
rect 151880 28480 152040 28640
rect 151880 28640 152040 28800
rect 151880 28800 152040 28960
rect 151880 28960 152040 29120
rect 151880 29120 152040 29280
rect 151880 29280 152040 29440
rect 151880 29440 152040 29600
rect 151880 29600 152040 29760
rect 151880 29760 152040 29920
rect 151880 29920 152040 30080
rect 151880 30080 152040 30240
rect 151880 30240 152040 30400
rect 151880 30400 152040 30560
rect 151880 30560 152040 30720
rect 151880 30720 152040 30880
rect 151880 30880 152040 31040
rect 151880 31040 152040 31200
rect 151880 31200 152040 31360
rect 151880 31360 152040 31520
rect 151880 31520 152040 31680
rect 151880 31680 152040 31840
rect 151880 31840 152040 32000
rect 151880 32000 152040 32160
rect 151880 32160 152040 32320
rect 151880 32320 152040 32480
rect 151880 32480 152040 32640
rect 151880 32640 152040 32800
rect 151880 32800 152040 32960
rect 151880 32960 152040 33120
rect 151880 33120 152040 33280
rect 151880 33280 152040 33440
rect 151880 33440 152040 33600
rect 151880 33600 152040 33760
rect 151880 33760 152040 33920
rect 151880 33920 152040 34080
rect 151880 34080 152040 34240
rect 151880 34240 152040 34400
rect 151880 34400 152040 34560
rect 151880 34560 152040 34720
rect 151880 34720 152040 34880
rect 151880 34880 152040 35040
rect 151880 35040 152040 35200
rect 151880 35200 152040 35360
rect 151880 35360 152040 35520
rect 151880 35520 152040 35680
rect 151880 35680 152040 35840
rect 151880 35840 152040 36000
rect 151880 36000 152040 36160
rect 151880 36160 152040 36320
rect 151880 36320 152040 36480
rect 151880 36480 152040 36640
rect 151880 36640 152040 36800
rect 151880 36800 152040 36960
rect 151880 36960 152040 37120
rect 151880 37120 152040 37280
rect 151880 37280 152040 37440
rect 151880 37440 152040 37600
rect 151880 37600 152040 37760
rect 151880 37760 152040 37920
rect 151880 37920 152040 38080
rect 151880 38080 152040 38240
rect 151880 38240 152040 38400
rect 151880 40640 152040 40800
rect 151880 40800 152040 40960
rect 151880 40960 152040 41120
rect 151880 41120 152040 41280
rect 151880 41280 152040 41440
rect 151880 41440 152040 41600
rect 151880 41600 152040 41760
rect 151880 41760 152040 41920
rect 151880 41920 152040 42080
rect 151880 42080 152040 42240
rect 151880 42240 152040 42400
rect 151880 42400 152040 42560
rect 151880 42560 152040 42720
rect 151880 42720 152040 42880
rect 151880 42880 152040 43040
rect 151880 43040 152040 43200
rect 151880 43200 152040 43360
rect 151880 43360 152040 43520
rect 151880 43520 152040 43680
rect 151880 43680 152040 43840
rect 151880 43840 152040 44000
rect 151880 44000 152040 44160
rect 151880 44160 152040 44320
rect 151880 44320 152040 44480
rect 151880 44480 152040 44640
rect 151880 44640 152040 44800
rect 151880 44800 152040 44960
rect 151880 44960 152040 45120
rect 151880 45120 152040 45280
rect 151880 45280 152040 45440
rect 151880 45440 152040 45600
rect 151880 45600 152040 45760
rect 151880 45760 152040 45920
rect 151880 45920 152040 46080
rect 151880 46080 152040 46240
rect 151880 46240 152040 46400
rect 151880 46400 152040 46560
rect 151880 46560 152040 46720
rect 151880 46720 152040 46880
rect 151880 46880 152040 47040
rect 151880 47040 152040 47200
rect 151880 47200 152040 47360
rect 151880 47360 152040 47520
rect 151880 47520 152040 47680
rect 151880 47680 152040 47840
rect 151880 47840 152040 48000
rect 151880 48000 152040 48160
rect 151880 48160 152040 48320
rect 151880 48320 152040 48480
rect 151880 48480 152040 48640
rect 151880 48640 152040 48800
rect 151880 48800 152040 48960
rect 151880 48960 152040 49120
rect 151880 49120 152040 49280
rect 151880 49280 152040 49440
rect 151880 49440 152040 49600
rect 151880 49600 152040 49760
rect 151880 49760 152040 49920
rect 151880 49920 152040 50080
rect 151880 50080 152040 50240
rect 151880 50240 152040 50400
rect 151880 50400 152040 50560
rect 151880 50560 152040 50720
rect 151880 50720 152040 50880
rect 151880 50880 152040 51040
rect 151880 51040 152040 51200
rect 151880 51200 152040 51360
rect 151880 51360 152040 51520
rect 151880 51520 152040 51680
rect 151880 51680 152040 51840
rect 151880 51840 152040 52000
rect 151880 52000 152040 52160
rect 151880 52160 152040 52320
rect 151880 52320 152040 52480
rect 151880 52480 152040 52640
rect 151880 52640 152040 52800
rect 151880 52800 152040 52960
rect 151880 52960 152040 53120
rect 151880 53120 152040 53280
rect 152040 25920 152200 26080
rect 152040 26080 152200 26240
rect 152040 26240 152200 26400
rect 152040 26400 152200 26560
rect 152040 26560 152200 26720
rect 152040 26720 152200 26880
rect 152040 26880 152200 27040
rect 152040 27040 152200 27200
rect 152040 27200 152200 27360
rect 152040 27360 152200 27520
rect 152040 27520 152200 27680
rect 152040 27680 152200 27840
rect 152040 27840 152200 28000
rect 152040 28000 152200 28160
rect 152040 28160 152200 28320
rect 152040 28320 152200 28480
rect 152040 28480 152200 28640
rect 152040 28640 152200 28800
rect 152040 28800 152200 28960
rect 152040 28960 152200 29120
rect 152040 29120 152200 29280
rect 152040 29280 152200 29440
rect 152040 29440 152200 29600
rect 152040 29600 152200 29760
rect 152040 29760 152200 29920
rect 152040 29920 152200 30080
rect 152040 30080 152200 30240
rect 152040 30240 152200 30400
rect 152040 30400 152200 30560
rect 152040 30560 152200 30720
rect 152040 30720 152200 30880
rect 152040 30880 152200 31040
rect 152040 31040 152200 31200
rect 152040 31200 152200 31360
rect 152040 31360 152200 31520
rect 152040 31520 152200 31680
rect 152040 31680 152200 31840
rect 152040 31840 152200 32000
rect 152040 32000 152200 32160
rect 152040 32160 152200 32320
rect 152040 32320 152200 32480
rect 152040 32480 152200 32640
rect 152040 32640 152200 32800
rect 152040 32800 152200 32960
rect 152040 32960 152200 33120
rect 152040 33120 152200 33280
rect 152040 33280 152200 33440
rect 152040 33440 152200 33600
rect 152040 33600 152200 33760
rect 152040 33760 152200 33920
rect 152040 33920 152200 34080
rect 152040 34080 152200 34240
rect 152040 34240 152200 34400
rect 152040 34400 152200 34560
rect 152040 34560 152200 34720
rect 152040 34720 152200 34880
rect 152040 34880 152200 35040
rect 152040 35040 152200 35200
rect 152040 35200 152200 35360
rect 152040 35360 152200 35520
rect 152040 35520 152200 35680
rect 152040 35680 152200 35840
rect 152040 35840 152200 36000
rect 152040 36000 152200 36160
rect 152040 36160 152200 36320
rect 152040 36320 152200 36480
rect 152040 36480 152200 36640
rect 152040 36640 152200 36800
rect 152040 36800 152200 36960
rect 152040 36960 152200 37120
rect 152040 37120 152200 37280
rect 152040 37280 152200 37440
rect 152040 37440 152200 37600
rect 152040 37600 152200 37760
rect 152040 37760 152200 37920
rect 152040 37920 152200 38080
rect 152040 38080 152200 38240
rect 152040 38240 152200 38400
rect 152040 40640 152200 40800
rect 152040 40800 152200 40960
rect 152040 40960 152200 41120
rect 152040 41120 152200 41280
rect 152040 41280 152200 41440
rect 152040 41440 152200 41600
rect 152040 41600 152200 41760
rect 152040 41760 152200 41920
rect 152040 41920 152200 42080
rect 152040 42080 152200 42240
rect 152040 42240 152200 42400
rect 152040 42400 152200 42560
rect 152040 42560 152200 42720
rect 152040 42720 152200 42880
rect 152040 42880 152200 43040
rect 152040 43040 152200 43200
rect 152040 43200 152200 43360
rect 152040 43360 152200 43520
rect 152040 43520 152200 43680
rect 152040 43680 152200 43840
rect 152040 43840 152200 44000
rect 152040 44000 152200 44160
rect 152040 44160 152200 44320
rect 152040 44320 152200 44480
rect 152040 44480 152200 44640
rect 152040 44640 152200 44800
rect 152040 44800 152200 44960
rect 152040 44960 152200 45120
rect 152040 45120 152200 45280
rect 152040 45280 152200 45440
rect 152040 45440 152200 45600
rect 152040 45600 152200 45760
rect 152040 45760 152200 45920
rect 152040 45920 152200 46080
rect 152040 46080 152200 46240
rect 152040 46240 152200 46400
rect 152040 46400 152200 46560
rect 152040 46560 152200 46720
rect 152040 46720 152200 46880
rect 152040 46880 152200 47040
rect 152040 47040 152200 47200
rect 152040 47200 152200 47360
rect 152040 47360 152200 47520
rect 152040 47520 152200 47680
rect 152040 47680 152200 47840
rect 152040 47840 152200 48000
rect 152040 48000 152200 48160
rect 152040 48160 152200 48320
rect 152040 48320 152200 48480
rect 152040 48480 152200 48640
rect 152040 48640 152200 48800
rect 152040 48800 152200 48960
rect 152040 48960 152200 49120
rect 152040 49120 152200 49280
rect 152040 49280 152200 49440
rect 152040 49440 152200 49600
rect 152040 49600 152200 49760
rect 152040 49760 152200 49920
rect 152040 49920 152200 50080
rect 152040 50080 152200 50240
rect 152040 50240 152200 50400
rect 152040 50400 152200 50560
rect 152040 50560 152200 50720
rect 152040 50720 152200 50880
rect 152040 50880 152200 51040
rect 152040 51040 152200 51200
rect 152040 51200 152200 51360
rect 152040 51360 152200 51520
rect 152040 51520 152200 51680
rect 152040 51680 152200 51840
rect 152040 51840 152200 52000
rect 152040 52000 152200 52160
rect 152040 52160 152200 52320
rect 152040 52320 152200 52480
rect 152040 52480 152200 52640
rect 152040 52640 152200 52800
rect 152040 52800 152200 52960
rect 152040 52960 152200 53120
rect 152040 53120 152200 53280
rect 152200 26080 152360 26240
rect 152200 26240 152360 26400
rect 152200 26400 152360 26560
rect 152200 26560 152360 26720
rect 152200 26720 152360 26880
rect 152200 26880 152360 27040
rect 152200 27040 152360 27200
rect 152200 27200 152360 27360
rect 152200 27360 152360 27520
rect 152200 27520 152360 27680
rect 152200 27680 152360 27840
rect 152200 27840 152360 28000
rect 152200 28000 152360 28160
rect 152200 28160 152360 28320
rect 152200 28320 152360 28480
rect 152200 28480 152360 28640
rect 152200 28640 152360 28800
rect 152200 28800 152360 28960
rect 152200 28960 152360 29120
rect 152200 29120 152360 29280
rect 152200 29280 152360 29440
rect 152200 29440 152360 29600
rect 152200 29600 152360 29760
rect 152200 29760 152360 29920
rect 152200 29920 152360 30080
rect 152200 30080 152360 30240
rect 152200 30240 152360 30400
rect 152200 30400 152360 30560
rect 152200 30560 152360 30720
rect 152200 30720 152360 30880
rect 152200 30880 152360 31040
rect 152200 31040 152360 31200
rect 152200 31200 152360 31360
rect 152200 31360 152360 31520
rect 152200 31520 152360 31680
rect 152200 31680 152360 31840
rect 152200 31840 152360 32000
rect 152200 32000 152360 32160
rect 152200 32160 152360 32320
rect 152200 32320 152360 32480
rect 152200 32480 152360 32640
rect 152200 32640 152360 32800
rect 152200 32800 152360 32960
rect 152200 32960 152360 33120
rect 152200 33120 152360 33280
rect 152200 33280 152360 33440
rect 152200 33440 152360 33600
rect 152200 33600 152360 33760
rect 152200 33760 152360 33920
rect 152200 33920 152360 34080
rect 152200 34080 152360 34240
rect 152200 34240 152360 34400
rect 152200 34400 152360 34560
rect 152200 34560 152360 34720
rect 152200 34720 152360 34880
rect 152200 34880 152360 35040
rect 152200 35040 152360 35200
rect 152200 35200 152360 35360
rect 152200 35360 152360 35520
rect 152200 35520 152360 35680
rect 152200 35680 152360 35840
rect 152200 35840 152360 36000
rect 152200 36000 152360 36160
rect 152200 36160 152360 36320
rect 152200 36320 152360 36480
rect 152200 36480 152360 36640
rect 152200 36640 152360 36800
rect 152200 36800 152360 36960
rect 152200 36960 152360 37120
rect 152200 37120 152360 37280
rect 152200 37280 152360 37440
rect 152200 37440 152360 37600
rect 152200 37600 152360 37760
rect 152200 37760 152360 37920
rect 152200 37920 152360 38080
rect 152200 38080 152360 38240
rect 152200 38240 152360 38400
rect 152200 40800 152360 40960
rect 152200 40960 152360 41120
rect 152200 41120 152360 41280
rect 152200 41280 152360 41440
rect 152200 41440 152360 41600
rect 152200 41600 152360 41760
rect 152200 41760 152360 41920
rect 152200 41920 152360 42080
rect 152200 42080 152360 42240
rect 152200 42240 152360 42400
rect 152200 42400 152360 42560
rect 152200 42560 152360 42720
rect 152200 42720 152360 42880
rect 152200 42880 152360 43040
rect 152200 43040 152360 43200
rect 152200 43200 152360 43360
rect 152200 43360 152360 43520
rect 152200 43520 152360 43680
rect 152200 43680 152360 43840
rect 152200 43840 152360 44000
rect 152200 44000 152360 44160
rect 152200 44160 152360 44320
rect 152200 44320 152360 44480
rect 152200 44480 152360 44640
rect 152200 44640 152360 44800
rect 152200 44800 152360 44960
rect 152200 44960 152360 45120
rect 152200 45120 152360 45280
rect 152200 45280 152360 45440
rect 152200 45440 152360 45600
rect 152200 45600 152360 45760
rect 152200 45760 152360 45920
rect 152200 45920 152360 46080
rect 152200 46080 152360 46240
rect 152200 46240 152360 46400
rect 152200 46400 152360 46560
rect 152200 46560 152360 46720
rect 152200 46720 152360 46880
rect 152200 46880 152360 47040
rect 152200 47040 152360 47200
rect 152200 47200 152360 47360
rect 152200 47360 152360 47520
rect 152200 47520 152360 47680
rect 152200 47680 152360 47840
rect 152200 47840 152360 48000
rect 152200 48000 152360 48160
rect 152200 48160 152360 48320
rect 152200 48320 152360 48480
rect 152200 48480 152360 48640
rect 152200 48640 152360 48800
rect 152200 48800 152360 48960
rect 152200 48960 152360 49120
rect 152200 49120 152360 49280
rect 152200 49280 152360 49440
rect 152200 49440 152360 49600
rect 152200 49600 152360 49760
rect 152200 49760 152360 49920
rect 152200 49920 152360 50080
rect 152200 50080 152360 50240
rect 152200 50240 152360 50400
rect 152200 50400 152360 50560
rect 152200 50560 152360 50720
rect 152200 50720 152360 50880
rect 152200 50880 152360 51040
rect 152200 51040 152360 51200
rect 152200 51200 152360 51360
rect 152200 51360 152360 51520
rect 152200 51520 152360 51680
rect 152200 51680 152360 51840
rect 152200 51840 152360 52000
rect 152200 52000 152360 52160
rect 152200 52160 152360 52320
rect 152200 52320 152360 52480
rect 152200 52480 152360 52640
rect 152200 52640 152360 52800
rect 152200 52800 152360 52960
rect 152200 52960 152360 53120
rect 152360 26240 152520 26400
rect 152360 26400 152520 26560
rect 152360 26560 152520 26720
rect 152360 26720 152520 26880
rect 152360 26880 152520 27040
rect 152360 27040 152520 27200
rect 152360 27200 152520 27360
rect 152360 27360 152520 27520
rect 152360 27520 152520 27680
rect 152360 27680 152520 27840
rect 152360 27840 152520 28000
rect 152360 28000 152520 28160
rect 152360 28160 152520 28320
rect 152360 28320 152520 28480
rect 152360 28480 152520 28640
rect 152360 28640 152520 28800
rect 152360 28800 152520 28960
rect 152360 28960 152520 29120
rect 152360 29120 152520 29280
rect 152360 29280 152520 29440
rect 152360 29440 152520 29600
rect 152360 29600 152520 29760
rect 152360 29760 152520 29920
rect 152360 29920 152520 30080
rect 152360 30080 152520 30240
rect 152360 30240 152520 30400
rect 152360 30400 152520 30560
rect 152360 30560 152520 30720
rect 152360 30720 152520 30880
rect 152360 30880 152520 31040
rect 152360 31040 152520 31200
rect 152360 31200 152520 31360
rect 152360 31360 152520 31520
rect 152360 31520 152520 31680
rect 152360 31680 152520 31840
rect 152360 31840 152520 32000
rect 152360 32000 152520 32160
rect 152360 32160 152520 32320
rect 152360 32320 152520 32480
rect 152360 32480 152520 32640
rect 152360 32640 152520 32800
rect 152360 32800 152520 32960
rect 152360 32960 152520 33120
rect 152360 33120 152520 33280
rect 152360 33280 152520 33440
rect 152360 33440 152520 33600
rect 152360 33600 152520 33760
rect 152360 33760 152520 33920
rect 152360 33920 152520 34080
rect 152360 34080 152520 34240
rect 152360 34240 152520 34400
rect 152360 34400 152520 34560
rect 152360 34560 152520 34720
rect 152360 34720 152520 34880
rect 152360 34880 152520 35040
rect 152360 35040 152520 35200
rect 152360 35200 152520 35360
rect 152360 35360 152520 35520
rect 152360 35520 152520 35680
rect 152360 35680 152520 35840
rect 152360 35840 152520 36000
rect 152360 36000 152520 36160
rect 152360 36160 152520 36320
rect 152360 36320 152520 36480
rect 152360 36480 152520 36640
rect 152360 36640 152520 36800
rect 152360 36800 152520 36960
rect 152360 36960 152520 37120
rect 152360 37120 152520 37280
rect 152360 37280 152520 37440
rect 152360 37440 152520 37600
rect 152360 37600 152520 37760
rect 152360 37760 152520 37920
rect 152360 37920 152520 38080
rect 152360 38080 152520 38240
rect 152360 40800 152520 40960
rect 152360 40960 152520 41120
rect 152360 41120 152520 41280
rect 152360 41280 152520 41440
rect 152360 41440 152520 41600
rect 152360 41600 152520 41760
rect 152360 41760 152520 41920
rect 152360 41920 152520 42080
rect 152360 42080 152520 42240
rect 152360 42240 152520 42400
rect 152360 42400 152520 42560
rect 152360 42560 152520 42720
rect 152360 42720 152520 42880
rect 152360 42880 152520 43040
rect 152360 43040 152520 43200
rect 152360 43200 152520 43360
rect 152360 43360 152520 43520
rect 152360 43520 152520 43680
rect 152360 43680 152520 43840
rect 152360 43840 152520 44000
rect 152360 44000 152520 44160
rect 152360 44160 152520 44320
rect 152360 44320 152520 44480
rect 152360 44480 152520 44640
rect 152360 44640 152520 44800
rect 152360 44800 152520 44960
rect 152360 44960 152520 45120
rect 152360 45120 152520 45280
rect 152360 45280 152520 45440
rect 152360 45440 152520 45600
rect 152360 45600 152520 45760
rect 152360 45760 152520 45920
rect 152360 45920 152520 46080
rect 152360 46080 152520 46240
rect 152360 46240 152520 46400
rect 152360 46400 152520 46560
rect 152360 46560 152520 46720
rect 152360 46720 152520 46880
rect 152360 46880 152520 47040
rect 152360 47040 152520 47200
rect 152360 47200 152520 47360
rect 152360 47360 152520 47520
rect 152360 47520 152520 47680
rect 152360 47680 152520 47840
rect 152360 47840 152520 48000
rect 152360 48000 152520 48160
rect 152360 48160 152520 48320
rect 152360 48320 152520 48480
rect 152360 48480 152520 48640
rect 152360 48640 152520 48800
rect 152360 48800 152520 48960
rect 152360 48960 152520 49120
rect 152360 49120 152520 49280
rect 152360 49280 152520 49440
rect 152360 49440 152520 49600
rect 152360 49600 152520 49760
rect 152360 49760 152520 49920
rect 152360 49920 152520 50080
rect 152360 50080 152520 50240
rect 152360 50240 152520 50400
rect 152360 50400 152520 50560
rect 152360 50560 152520 50720
rect 152360 50720 152520 50880
rect 152360 50880 152520 51040
rect 152360 51040 152520 51200
rect 152360 51200 152520 51360
rect 152360 51360 152520 51520
rect 152360 51520 152520 51680
rect 152360 51680 152520 51840
rect 152360 51840 152520 52000
rect 152360 52000 152520 52160
rect 152360 52160 152520 52320
rect 152360 52320 152520 52480
rect 152360 52480 152520 52640
rect 152360 52640 152520 52800
rect 152360 52800 152520 52960
rect 152360 52960 152520 53120
rect 152520 26560 152680 26720
rect 152520 26720 152680 26880
rect 152520 26880 152680 27040
rect 152520 27040 152680 27200
rect 152520 27200 152680 27360
rect 152520 27360 152680 27520
rect 152520 27520 152680 27680
rect 152520 27680 152680 27840
rect 152520 27840 152680 28000
rect 152520 28000 152680 28160
rect 152520 28160 152680 28320
rect 152520 28320 152680 28480
rect 152520 28480 152680 28640
rect 152520 28640 152680 28800
rect 152520 28800 152680 28960
rect 152520 28960 152680 29120
rect 152520 29120 152680 29280
rect 152520 29280 152680 29440
rect 152520 29440 152680 29600
rect 152520 29600 152680 29760
rect 152520 29760 152680 29920
rect 152520 29920 152680 30080
rect 152520 30080 152680 30240
rect 152520 30240 152680 30400
rect 152520 30400 152680 30560
rect 152520 30560 152680 30720
rect 152520 30720 152680 30880
rect 152520 30880 152680 31040
rect 152520 31040 152680 31200
rect 152520 31200 152680 31360
rect 152520 31360 152680 31520
rect 152520 31520 152680 31680
rect 152520 31680 152680 31840
rect 152520 31840 152680 32000
rect 152520 32000 152680 32160
rect 152520 32160 152680 32320
rect 152520 32320 152680 32480
rect 152520 32480 152680 32640
rect 152520 32640 152680 32800
rect 152520 32800 152680 32960
rect 152520 32960 152680 33120
rect 152520 33120 152680 33280
rect 152520 33280 152680 33440
rect 152520 33440 152680 33600
rect 152520 33600 152680 33760
rect 152520 33760 152680 33920
rect 152520 33920 152680 34080
rect 152520 34080 152680 34240
rect 152520 34240 152680 34400
rect 152520 34400 152680 34560
rect 152520 34560 152680 34720
rect 152520 34720 152680 34880
rect 152520 34880 152680 35040
rect 152520 35040 152680 35200
rect 152520 35200 152680 35360
rect 152520 35360 152680 35520
rect 152520 35520 152680 35680
rect 152520 35680 152680 35840
rect 152520 35840 152680 36000
rect 152520 36000 152680 36160
rect 152520 36160 152680 36320
rect 152520 36320 152680 36480
rect 152520 36480 152680 36640
rect 152520 36640 152680 36800
rect 152520 36800 152680 36960
rect 152520 36960 152680 37120
rect 152520 37120 152680 37280
rect 152520 37280 152680 37440
rect 152520 37440 152680 37600
rect 152520 37600 152680 37760
rect 152520 37760 152680 37920
rect 152520 37920 152680 38080
rect 152520 38080 152680 38240
rect 152520 38240 152680 38400
rect 152520 40960 152680 41120
rect 152520 41120 152680 41280
rect 152520 41280 152680 41440
rect 152520 41440 152680 41600
rect 152520 41600 152680 41760
rect 152520 41760 152680 41920
rect 152520 41920 152680 42080
rect 152520 42080 152680 42240
rect 152520 42240 152680 42400
rect 152520 42400 152680 42560
rect 152520 42560 152680 42720
rect 152520 42720 152680 42880
rect 152520 42880 152680 43040
rect 152520 43040 152680 43200
rect 152520 43200 152680 43360
rect 152520 43360 152680 43520
rect 152520 43520 152680 43680
rect 152520 43680 152680 43840
rect 152520 43840 152680 44000
rect 152520 44000 152680 44160
rect 152520 44160 152680 44320
rect 152520 44320 152680 44480
rect 152520 44480 152680 44640
rect 152520 44640 152680 44800
rect 152520 44800 152680 44960
rect 152520 44960 152680 45120
rect 152520 45120 152680 45280
rect 152520 45280 152680 45440
rect 152520 45440 152680 45600
rect 152520 45600 152680 45760
rect 152520 45760 152680 45920
rect 152520 45920 152680 46080
rect 152520 46080 152680 46240
rect 152520 46240 152680 46400
rect 152520 46400 152680 46560
rect 152520 46560 152680 46720
rect 152520 46720 152680 46880
rect 152520 46880 152680 47040
rect 152520 47040 152680 47200
rect 152520 47200 152680 47360
rect 152520 47360 152680 47520
rect 152520 47520 152680 47680
rect 152520 47680 152680 47840
rect 152520 47840 152680 48000
rect 152520 48000 152680 48160
rect 152520 48160 152680 48320
rect 152520 48320 152680 48480
rect 152520 48480 152680 48640
rect 152520 48640 152680 48800
rect 152520 48800 152680 48960
rect 152520 48960 152680 49120
rect 152520 49120 152680 49280
rect 152520 49280 152680 49440
rect 152520 49440 152680 49600
rect 152520 49600 152680 49760
rect 152520 49760 152680 49920
rect 152520 49920 152680 50080
rect 152520 50080 152680 50240
rect 152520 50240 152680 50400
rect 152520 50400 152680 50560
rect 152520 50560 152680 50720
rect 152520 50720 152680 50880
rect 152520 50880 152680 51040
rect 152520 51040 152680 51200
rect 152520 51200 152680 51360
rect 152520 51360 152680 51520
rect 152520 51520 152680 51680
rect 152520 51680 152680 51840
rect 152520 51840 152680 52000
rect 152520 52000 152680 52160
rect 152520 52160 152680 52320
rect 152520 52320 152680 52480
rect 152520 52480 152680 52640
rect 152520 52640 152680 52800
rect 152520 52800 152680 52960
rect 152680 27040 152840 27200
rect 152680 27200 152840 27360
rect 152680 27360 152840 27520
rect 152680 27520 152840 27680
rect 152680 27680 152840 27840
rect 152680 27840 152840 28000
rect 152680 28000 152840 28160
rect 152680 28160 152840 28320
rect 152680 28320 152840 28480
rect 152680 28480 152840 28640
rect 152680 28640 152840 28800
rect 152680 28800 152840 28960
rect 152680 28960 152840 29120
rect 152680 29120 152840 29280
rect 152680 29280 152840 29440
rect 152680 29440 152840 29600
rect 152680 29600 152840 29760
rect 152680 29760 152840 29920
rect 152680 29920 152840 30080
rect 152680 30080 152840 30240
rect 152680 30240 152840 30400
rect 152680 30400 152840 30560
rect 152680 30560 152840 30720
rect 152680 30720 152840 30880
rect 152680 30880 152840 31040
rect 152680 31040 152840 31200
rect 152680 31200 152840 31360
rect 152680 31360 152840 31520
rect 152680 31520 152840 31680
rect 152680 31680 152840 31840
rect 152680 31840 152840 32000
rect 152680 32000 152840 32160
rect 152680 32160 152840 32320
rect 152680 32320 152840 32480
rect 152680 32480 152840 32640
rect 152680 32640 152840 32800
rect 152680 32800 152840 32960
rect 152680 32960 152840 33120
rect 152680 33120 152840 33280
rect 152680 33280 152840 33440
rect 152680 33440 152840 33600
rect 152680 33600 152840 33760
rect 152680 33760 152840 33920
rect 152680 33920 152840 34080
rect 152680 34080 152840 34240
rect 152680 34240 152840 34400
rect 152680 34400 152840 34560
rect 152680 34560 152840 34720
rect 152680 34720 152840 34880
rect 152680 34880 152840 35040
rect 152680 35040 152840 35200
rect 152680 35200 152840 35360
rect 152680 35360 152840 35520
rect 152680 35520 152840 35680
rect 152680 35680 152840 35840
rect 152680 35840 152840 36000
rect 152680 36000 152840 36160
rect 152680 36160 152840 36320
rect 152680 36320 152840 36480
rect 152680 36480 152840 36640
rect 152680 36640 152840 36800
rect 152680 36800 152840 36960
rect 152680 36960 152840 37120
rect 152680 37120 152840 37280
rect 152680 37280 152840 37440
rect 152680 37440 152840 37600
rect 152680 37600 152840 37760
rect 152680 37760 152840 37920
rect 152680 37920 152840 38080
rect 152680 38080 152840 38240
rect 152680 38240 152840 38400
rect 152680 40960 152840 41120
rect 152680 41120 152840 41280
rect 152680 41280 152840 41440
rect 152680 41440 152840 41600
rect 152680 41600 152840 41760
rect 152680 41760 152840 41920
rect 152680 41920 152840 42080
rect 152680 42080 152840 42240
rect 152680 42240 152840 42400
rect 152680 42400 152840 42560
rect 152680 42560 152840 42720
rect 152680 42720 152840 42880
rect 152680 42880 152840 43040
rect 152680 43040 152840 43200
rect 152680 43200 152840 43360
rect 152680 43360 152840 43520
rect 152680 43520 152840 43680
rect 152680 43680 152840 43840
rect 152680 43840 152840 44000
rect 152680 44000 152840 44160
rect 152680 44160 152840 44320
rect 152680 44320 152840 44480
rect 152680 44480 152840 44640
rect 152680 44640 152840 44800
rect 152680 44800 152840 44960
rect 152680 44960 152840 45120
rect 152680 45120 152840 45280
rect 152680 45280 152840 45440
rect 152680 45440 152840 45600
rect 152680 45600 152840 45760
rect 152680 45760 152840 45920
rect 152680 45920 152840 46080
rect 152680 46080 152840 46240
rect 152680 46240 152840 46400
rect 152680 46400 152840 46560
rect 152680 46560 152840 46720
rect 152680 46720 152840 46880
rect 152680 46880 152840 47040
rect 152680 47040 152840 47200
rect 152680 47200 152840 47360
rect 152680 47360 152840 47520
rect 152680 47520 152840 47680
rect 152680 47680 152840 47840
rect 152680 47840 152840 48000
rect 152680 48000 152840 48160
rect 152680 48160 152840 48320
rect 152680 48320 152840 48480
rect 152680 48480 152840 48640
rect 152680 48640 152840 48800
rect 152680 48800 152840 48960
rect 152680 48960 152840 49120
rect 152680 49120 152840 49280
rect 152680 49280 152840 49440
rect 152680 49440 152840 49600
rect 152680 49600 152840 49760
rect 152680 49760 152840 49920
rect 152680 49920 152840 50080
rect 152680 50080 152840 50240
rect 152680 50240 152840 50400
rect 152680 50400 152840 50560
rect 152680 50560 152840 50720
rect 152680 50720 152840 50880
rect 152680 50880 152840 51040
rect 152680 51040 152840 51200
rect 152680 51200 152840 51360
rect 152680 51360 152840 51520
rect 152680 51520 152840 51680
rect 152680 51680 152840 51840
rect 152680 51840 152840 52000
rect 152680 52000 152840 52160
rect 152680 52160 152840 52320
rect 152680 52320 152840 52480
rect 152680 52480 152840 52640
rect 152680 52640 152840 52800
rect 152840 35680 153000 35840
rect 152840 35840 153000 36000
rect 152840 36000 153000 36160
rect 152840 36160 153000 36320
rect 152840 36320 153000 36480
rect 152840 36480 153000 36640
rect 152840 36640 153000 36800
rect 152840 36800 153000 36960
rect 152840 36960 153000 37120
rect 152840 37120 153000 37280
rect 152840 37280 153000 37440
rect 152840 37440 153000 37600
rect 152840 37600 153000 37760
rect 152840 37760 153000 37920
rect 152840 37920 153000 38080
rect 152840 38080 153000 38240
rect 152840 38240 153000 38400
rect 152840 40960 153000 41120
rect 152840 41120 153000 41280
rect 152840 41280 153000 41440
rect 152840 41440 153000 41600
rect 152840 41600 153000 41760
rect 152840 41760 153000 41920
rect 152840 41920 153000 42080
rect 152840 42080 153000 42240
rect 152840 42240 153000 42400
rect 152840 42400 153000 42560
rect 152840 42560 153000 42720
rect 152840 42720 153000 42880
rect 152840 42880 153000 43040
rect 152840 43040 153000 43200
rect 152840 43200 153000 43360
rect 152840 43360 153000 43520
rect 152840 45920 153000 46080
rect 152840 46240 153000 46400
rect 152840 46400 153000 46560
rect 152840 46560 153000 46720
rect 152840 46720 153000 46880
rect 152840 46880 153000 47040
rect 152840 47040 153000 47200
rect 152840 47200 153000 47360
rect 152840 47360 153000 47520
rect 152840 47520 153000 47680
rect 152840 47680 153000 47840
rect 152840 47840 153000 48000
rect 152840 48000 153000 48160
rect 152840 48160 153000 48320
rect 152840 48320 153000 48480
rect 152840 48480 153000 48640
rect 152840 48640 153000 48800
rect 152840 48800 153000 48960
rect 152840 48960 153000 49120
rect 152840 49120 153000 49280
rect 152840 49280 153000 49440
rect 152840 49440 153000 49600
rect 152840 49600 153000 49760
rect 152840 49760 153000 49920
rect 152840 49920 153000 50080
rect 152840 50080 153000 50240
rect 152840 50240 153000 50400
rect 152840 50400 153000 50560
rect 152840 50560 153000 50720
rect 152840 50720 153000 50880
rect 152840 50880 153000 51040
rect 152840 51040 153000 51200
rect 152840 51200 153000 51360
rect 152840 51360 153000 51520
rect 152840 51520 153000 51680
rect 152840 51680 153000 51840
rect 152840 51840 153000 52000
rect 152840 52000 153000 52160
rect 152840 52160 153000 52320
rect 152840 52320 153000 52480
rect 153000 35680 153160 35840
rect 153000 35840 153160 36000
rect 153000 36000 153160 36160
rect 153000 36160 153160 36320
rect 153000 36320 153160 36480
rect 153000 36480 153160 36640
rect 153000 36640 153160 36800
rect 153000 36800 153160 36960
rect 153000 36960 153160 37120
rect 153000 37120 153160 37280
rect 153000 37280 153160 37440
rect 153000 37440 153160 37600
rect 153000 37600 153160 37760
rect 153000 37760 153160 37920
rect 153000 37920 153160 38080
rect 153000 38080 153160 38240
rect 153000 38240 153160 38400
rect 153000 38400 153160 38560
rect 153000 40960 153160 41120
rect 153000 41120 153160 41280
rect 153000 41280 153160 41440
rect 153000 41440 153160 41600
rect 153000 41600 153160 41760
rect 153000 41760 153160 41920
rect 153000 41920 153160 42080
rect 153000 42080 153160 42240
rect 153000 42240 153160 42400
rect 153000 42400 153160 42560
rect 153000 42560 153160 42720
rect 153000 42720 153160 42880
rect 153000 42880 153160 43040
rect 153000 43040 153160 43200
rect 153000 43200 153160 43360
rect 153000 43360 153160 43520
rect 153000 49120 153160 49280
rect 153000 49440 153160 49600
rect 153000 49600 153160 49760
rect 153000 49760 153160 49920
rect 153000 49920 153160 50080
rect 153000 50080 153160 50240
rect 153000 50240 153160 50400
rect 153000 50400 153160 50560
rect 153000 50560 153160 50720
rect 153000 50720 153160 50880
rect 153000 50880 153160 51040
rect 153000 51040 153160 51200
rect 153000 51200 153160 51360
rect 153000 51360 153160 51520
rect 153000 51520 153160 51680
rect 153000 51680 153160 51840
rect 153000 51840 153160 52000
rect 153000 52000 153160 52160
rect 153160 35680 153320 35840
rect 153160 35840 153320 36000
rect 153160 36000 153320 36160
rect 153160 36160 153320 36320
rect 153160 36320 153320 36480
rect 153160 36480 153320 36640
rect 153160 36640 153320 36800
rect 153160 36800 153320 36960
rect 153160 36960 153320 37120
rect 153160 37120 153320 37280
rect 153160 37280 153320 37440
rect 153160 37440 153320 37600
rect 153160 37600 153320 37760
rect 153160 37760 153320 37920
rect 153160 37920 153320 38080
rect 153160 38080 153320 38240
rect 153160 38240 153320 38400
rect 153160 38400 153320 38560
rect 153160 40800 153320 40960
rect 153160 40960 153320 41120
rect 153160 41120 153320 41280
rect 153160 41280 153320 41440
rect 153160 41440 153320 41600
rect 153160 41600 153320 41760
rect 153160 41760 153320 41920
rect 153160 41920 153320 42080
rect 153160 42080 153320 42240
rect 153160 42240 153320 42400
rect 153160 42400 153320 42560
rect 153160 42560 153320 42720
rect 153160 42720 153320 42880
rect 153160 42880 153320 43040
rect 153160 43040 153320 43200
rect 153160 43200 153320 43360
rect 153320 35680 153480 35840
rect 153320 35840 153480 36000
rect 153320 36000 153480 36160
rect 153320 36160 153480 36320
rect 153320 36320 153480 36480
rect 153320 36480 153480 36640
rect 153320 36640 153480 36800
rect 153320 36800 153480 36960
rect 153320 36960 153480 37120
rect 153320 37120 153480 37280
rect 153320 37280 153480 37440
rect 153320 37440 153480 37600
rect 153320 37600 153480 37760
rect 153320 37760 153480 37920
rect 153320 37920 153480 38080
rect 153320 38080 153480 38240
rect 153320 38240 153480 38400
rect 153320 38400 153480 38560
rect 153320 38560 153480 38720
rect 153320 40800 153480 40960
rect 153320 40960 153480 41120
rect 153320 41120 153480 41280
rect 153320 41280 153480 41440
rect 153320 41440 153480 41600
rect 153320 41600 153480 41760
rect 153320 41760 153480 41920
rect 153320 41920 153480 42080
rect 153320 42080 153480 42240
rect 153320 42240 153480 42400
rect 153320 42400 153480 42560
rect 153320 42560 153480 42720
rect 153320 42720 153480 42880
rect 153320 42880 153480 43040
rect 153320 43040 153480 43200
rect 153320 43200 153480 43360
rect 153480 35680 153640 35840
rect 153480 35840 153640 36000
rect 153480 36000 153640 36160
rect 153480 36160 153640 36320
rect 153480 36320 153640 36480
rect 153480 36480 153640 36640
rect 153480 36640 153640 36800
rect 153480 36800 153640 36960
rect 153480 36960 153640 37120
rect 153480 37120 153640 37280
rect 153480 37280 153640 37440
rect 153480 37440 153640 37600
rect 153480 37600 153640 37760
rect 153480 37760 153640 37920
rect 153480 37920 153640 38080
rect 153480 38080 153640 38240
rect 153480 38240 153640 38400
rect 153480 38400 153640 38560
rect 153480 38560 153640 38720
rect 153480 38720 153640 38880
rect 153480 40640 153640 40800
rect 153480 40800 153640 40960
rect 153480 40960 153640 41120
rect 153480 41120 153640 41280
rect 153480 41280 153640 41440
rect 153480 41440 153640 41600
rect 153480 41600 153640 41760
rect 153480 41760 153640 41920
rect 153480 41920 153640 42080
rect 153480 42080 153640 42240
rect 153480 42240 153640 42400
rect 153480 42400 153640 42560
rect 153480 42560 153640 42720
rect 153480 42720 153640 42880
rect 153480 42880 153640 43040
rect 153480 43040 153640 43200
rect 153480 43200 153640 43360
rect 153640 35520 153800 35680
rect 153640 35680 153800 35840
rect 153640 35840 153800 36000
rect 153640 36000 153800 36160
rect 153640 36160 153800 36320
rect 153640 36320 153800 36480
rect 153640 36480 153800 36640
rect 153640 36640 153800 36800
rect 153640 36800 153800 36960
rect 153640 36960 153800 37120
rect 153640 37120 153800 37280
rect 153640 37280 153800 37440
rect 153640 37440 153800 37600
rect 153640 37600 153800 37760
rect 153640 37760 153800 37920
rect 153640 37920 153800 38080
rect 153640 38080 153800 38240
rect 153640 38240 153800 38400
rect 153640 38400 153800 38560
rect 153640 38560 153800 38720
rect 153640 38720 153800 38880
rect 153640 38880 153800 39040
rect 153640 40480 153800 40640
rect 153640 40640 153800 40800
rect 153640 40800 153800 40960
rect 153640 40960 153800 41120
rect 153640 41120 153800 41280
rect 153640 41280 153800 41440
rect 153640 41440 153800 41600
rect 153640 41600 153800 41760
rect 153640 41760 153800 41920
rect 153640 41920 153800 42080
rect 153640 42080 153800 42240
rect 153640 42240 153800 42400
rect 153640 42400 153800 42560
rect 153640 42560 153800 42720
rect 153640 42720 153800 42880
rect 153640 42880 153800 43040
rect 153640 43040 153800 43200
rect 153800 35360 153960 35520
rect 153800 35520 153960 35680
rect 153800 35680 153960 35840
rect 153800 35840 153960 36000
rect 153800 36000 153960 36160
rect 153800 36160 153960 36320
rect 153800 36320 153960 36480
rect 153800 36480 153960 36640
rect 153800 36640 153960 36800
rect 153800 36800 153960 36960
rect 153800 36960 153960 37120
rect 153800 37120 153960 37280
rect 153800 37280 153960 37440
rect 153800 37440 153960 37600
rect 153800 37600 153960 37760
rect 153800 37760 153960 37920
rect 153800 37920 153960 38080
rect 153800 38080 153960 38240
rect 153800 38240 153960 38400
rect 153800 38400 153960 38560
rect 153800 38560 153960 38720
rect 153800 38720 153960 38880
rect 153800 38880 153960 39040
rect 153800 39040 153960 39200
rect 153800 40320 153960 40480
rect 153800 40480 153960 40640
rect 153800 40640 153960 40800
rect 153800 40800 153960 40960
rect 153800 40960 153960 41120
rect 153800 41120 153960 41280
rect 153800 41280 153960 41440
rect 153800 41440 153960 41600
rect 153800 41600 153960 41760
rect 153800 41760 153960 41920
rect 153800 41920 153960 42080
rect 153800 42080 153960 42240
rect 153800 42240 153960 42400
rect 153800 42400 153960 42560
rect 153800 42560 153960 42720
rect 153800 42720 153960 42880
rect 153800 42880 153960 43040
rect 153800 43040 153960 43200
rect 153960 35200 154120 35360
rect 153960 35360 154120 35520
rect 153960 35520 154120 35680
rect 153960 35680 154120 35840
rect 153960 35840 154120 36000
rect 153960 36000 154120 36160
rect 153960 36160 154120 36320
rect 153960 36320 154120 36480
rect 153960 36480 154120 36640
rect 153960 36640 154120 36800
rect 153960 36800 154120 36960
rect 153960 36960 154120 37120
rect 153960 37120 154120 37280
rect 153960 37280 154120 37440
rect 153960 37440 154120 37600
rect 153960 37600 154120 37760
rect 153960 37760 154120 37920
rect 153960 37920 154120 38080
rect 153960 38080 154120 38240
rect 153960 38240 154120 38400
rect 153960 38400 154120 38560
rect 153960 38560 154120 38720
rect 153960 38720 154120 38880
rect 153960 38880 154120 39040
rect 153960 39040 154120 39200
rect 153960 39200 154120 39360
rect 153960 39360 154120 39520
rect 153960 39520 154120 39680
rect 153960 39680 154120 39840
rect 153960 39840 154120 40000
rect 153960 40000 154120 40160
rect 153960 40160 154120 40320
rect 153960 40320 154120 40480
rect 153960 40480 154120 40640
rect 153960 40640 154120 40800
rect 153960 40800 154120 40960
rect 153960 40960 154120 41120
rect 153960 41120 154120 41280
rect 153960 41280 154120 41440
rect 153960 41440 154120 41600
rect 153960 41600 154120 41760
rect 153960 41760 154120 41920
rect 153960 41920 154120 42080
rect 153960 42080 154120 42240
rect 153960 42240 154120 42400
rect 153960 42400 154120 42560
rect 153960 42560 154120 42720
rect 153960 42720 154120 42880
rect 153960 42880 154120 43040
rect 153960 43040 154120 43200
rect 154120 35040 154280 35200
rect 154120 35200 154280 35360
rect 154120 35360 154280 35520
rect 154120 35520 154280 35680
rect 154120 35680 154280 35840
rect 154120 35840 154280 36000
rect 154120 36000 154280 36160
rect 154120 36160 154280 36320
rect 154120 36320 154280 36480
rect 154120 36480 154280 36640
rect 154120 36640 154280 36800
rect 154120 36800 154280 36960
rect 154120 36960 154280 37120
rect 154120 37120 154280 37280
rect 154120 37280 154280 37440
rect 154120 37440 154280 37600
rect 154120 37600 154280 37760
rect 154120 37760 154280 37920
rect 154120 37920 154280 38080
rect 154120 38080 154280 38240
rect 154120 38240 154280 38400
rect 154120 38400 154280 38560
rect 154120 38560 154280 38720
rect 154120 38720 154280 38880
rect 154120 38880 154280 39040
rect 154120 39040 154280 39200
rect 154120 39200 154280 39360
rect 154120 39360 154280 39520
rect 154120 39520 154280 39680
rect 154120 39680 154280 39840
rect 154120 39840 154280 40000
rect 154120 40000 154280 40160
rect 154120 40160 154280 40320
rect 154120 40320 154280 40480
rect 154120 40480 154280 40640
rect 154120 40640 154280 40800
rect 154120 40800 154280 40960
rect 154120 40960 154280 41120
rect 154120 41120 154280 41280
rect 154120 41280 154280 41440
rect 154120 41440 154280 41600
rect 154120 41600 154280 41760
rect 154120 41760 154280 41920
rect 154120 41920 154280 42080
rect 154120 42080 154280 42240
rect 154120 42240 154280 42400
rect 154120 42400 154280 42560
rect 154120 42560 154280 42720
rect 154120 42720 154280 42880
rect 154120 42880 154280 43040
rect 154280 34880 154440 35040
rect 154280 35040 154440 35200
rect 154280 35200 154440 35360
rect 154280 35360 154440 35520
rect 154280 35520 154440 35680
rect 154280 35680 154440 35840
rect 154280 35840 154440 36000
rect 154280 36000 154440 36160
rect 154280 36160 154440 36320
rect 154280 36320 154440 36480
rect 154280 36480 154440 36640
rect 154280 36640 154440 36800
rect 154280 36800 154440 36960
rect 154280 36960 154440 37120
rect 154280 37120 154440 37280
rect 154280 37280 154440 37440
rect 154280 37440 154440 37600
rect 154280 37600 154440 37760
rect 154280 37760 154440 37920
rect 154280 37920 154440 38080
rect 154280 38080 154440 38240
rect 154280 38240 154440 38400
rect 154280 38400 154440 38560
rect 154280 38560 154440 38720
rect 154280 38720 154440 38880
rect 154280 38880 154440 39040
rect 154280 39040 154440 39200
rect 154280 39200 154440 39360
rect 154280 39360 154440 39520
rect 154280 39520 154440 39680
rect 154280 39680 154440 39840
rect 154280 39840 154440 40000
rect 154280 40000 154440 40160
rect 154280 40160 154440 40320
rect 154280 40320 154440 40480
rect 154280 40480 154440 40640
rect 154280 40640 154440 40800
rect 154280 40800 154440 40960
rect 154280 40960 154440 41120
rect 154280 41120 154440 41280
rect 154280 41280 154440 41440
rect 154280 41440 154440 41600
rect 154280 41600 154440 41760
rect 154280 41760 154440 41920
rect 154280 41920 154440 42080
rect 154280 42080 154440 42240
rect 154280 42240 154440 42400
rect 154280 42400 154440 42560
rect 154280 42560 154440 42720
rect 154280 42720 154440 42880
rect 154280 42880 154440 43040
rect 154440 34720 154600 34880
rect 154440 34880 154600 35040
rect 154440 35040 154600 35200
rect 154440 35200 154600 35360
rect 154440 35360 154600 35520
rect 154440 35520 154600 35680
rect 154440 35680 154600 35840
rect 154440 35840 154600 36000
rect 154440 36000 154600 36160
rect 154440 36160 154600 36320
rect 154440 36320 154600 36480
rect 154440 36480 154600 36640
rect 154440 36640 154600 36800
rect 154440 36800 154600 36960
rect 154440 36960 154600 37120
rect 154440 37120 154600 37280
rect 154440 37280 154600 37440
rect 154440 37440 154600 37600
rect 154440 37600 154600 37760
rect 154440 37760 154600 37920
rect 154440 37920 154600 38080
rect 154440 38080 154600 38240
rect 154440 38240 154600 38400
rect 154440 38400 154600 38560
rect 154440 38560 154600 38720
rect 154440 38720 154600 38880
rect 154440 38880 154600 39040
rect 154440 39040 154600 39200
rect 154440 39200 154600 39360
rect 154440 39360 154600 39520
rect 154440 39520 154600 39680
rect 154440 39680 154600 39840
rect 154440 39840 154600 40000
rect 154440 40000 154600 40160
rect 154440 40160 154600 40320
rect 154440 40320 154600 40480
rect 154440 40480 154600 40640
rect 154440 40640 154600 40800
rect 154440 40800 154600 40960
rect 154440 40960 154600 41120
rect 154440 41120 154600 41280
rect 154440 41280 154600 41440
rect 154440 41440 154600 41600
rect 154440 41600 154600 41760
rect 154440 41760 154600 41920
rect 154440 41920 154600 42080
rect 154440 42080 154600 42240
rect 154440 42240 154600 42400
rect 154440 42400 154600 42560
rect 154440 42560 154600 42720
rect 154440 42720 154600 42880
rect 154440 42880 154600 43040
rect 154440 43040 154600 43200
rect 154600 34560 154760 34720
rect 154600 34720 154760 34880
rect 154600 34880 154760 35040
rect 154600 35040 154760 35200
rect 154600 35200 154760 35360
rect 154600 35360 154760 35520
rect 154600 35520 154760 35680
rect 154600 35680 154760 35840
rect 154600 35840 154760 36000
rect 154600 36000 154760 36160
rect 154600 36160 154760 36320
rect 154600 36320 154760 36480
rect 154600 36480 154760 36640
rect 154600 36640 154760 36800
rect 154600 36800 154760 36960
rect 154600 36960 154760 37120
rect 154600 37120 154760 37280
rect 154600 37280 154760 37440
rect 154600 37440 154760 37600
rect 154600 37600 154760 37760
rect 154600 37760 154760 37920
rect 154600 37920 154760 38080
rect 154600 38080 154760 38240
rect 154600 38240 154760 38400
rect 154600 38400 154760 38560
rect 154600 38560 154760 38720
rect 154600 38720 154760 38880
rect 154600 38880 154760 39040
rect 154600 39040 154760 39200
rect 154600 39200 154760 39360
rect 154600 39360 154760 39520
rect 154600 39520 154760 39680
rect 154600 39680 154760 39840
rect 154600 39840 154760 40000
rect 154600 40000 154760 40160
rect 154600 40160 154760 40320
rect 154600 40320 154760 40480
rect 154600 40480 154760 40640
rect 154600 40640 154760 40800
rect 154600 40800 154760 40960
rect 154600 40960 154760 41120
rect 154600 41120 154760 41280
rect 154600 41280 154760 41440
rect 154600 41440 154760 41600
rect 154600 41600 154760 41760
rect 154600 41760 154760 41920
rect 154600 41920 154760 42080
rect 154600 42080 154760 42240
rect 154600 42240 154760 42400
rect 154600 42400 154760 42560
rect 154600 42560 154760 42720
rect 154600 42720 154760 42880
rect 154600 42880 154760 43040
rect 154600 43040 154760 43200
rect 154600 43200 154760 43360
rect 154760 34400 154920 34560
rect 154760 34560 154920 34720
rect 154760 34720 154920 34880
rect 154760 34880 154920 35040
rect 154760 35040 154920 35200
rect 154760 35200 154920 35360
rect 154760 35360 154920 35520
rect 154760 35520 154920 35680
rect 154760 35680 154920 35840
rect 154760 35840 154920 36000
rect 154760 36000 154920 36160
rect 154760 36160 154920 36320
rect 154760 36320 154920 36480
rect 154760 36480 154920 36640
rect 154760 36640 154920 36800
rect 154760 36800 154920 36960
rect 154760 36960 154920 37120
rect 154760 37120 154920 37280
rect 154760 37280 154920 37440
rect 154760 37440 154920 37600
rect 154760 37600 154920 37760
rect 154760 37760 154920 37920
rect 154760 37920 154920 38080
rect 154760 38080 154920 38240
rect 154760 38240 154920 38400
rect 154760 38400 154920 38560
rect 154760 38560 154920 38720
rect 154760 38720 154920 38880
rect 154760 38880 154920 39040
rect 154760 39040 154920 39200
rect 154760 39200 154920 39360
rect 154760 39360 154920 39520
rect 154760 39520 154920 39680
rect 154760 39680 154920 39840
rect 154760 39840 154920 40000
rect 154760 40000 154920 40160
rect 154760 40160 154920 40320
rect 154760 40320 154920 40480
rect 154760 40480 154920 40640
rect 154760 40640 154920 40800
rect 154760 40800 154920 40960
rect 154760 40960 154920 41120
rect 154760 41120 154920 41280
rect 154760 41280 154920 41440
rect 154760 41440 154920 41600
rect 154760 41600 154920 41760
rect 154760 41760 154920 41920
rect 154760 41920 154920 42080
rect 154760 42080 154920 42240
rect 154760 42240 154920 42400
rect 154760 42400 154920 42560
rect 154760 42560 154920 42720
rect 154760 42720 154920 42880
rect 154760 42880 154920 43040
rect 154760 43040 154920 43200
rect 154760 43200 154920 43360
rect 154760 43360 154920 43520
rect 154920 34240 155080 34400
rect 154920 34400 155080 34560
rect 154920 34560 155080 34720
rect 154920 34720 155080 34880
rect 154920 34880 155080 35040
rect 154920 35040 155080 35200
rect 154920 35200 155080 35360
rect 154920 35360 155080 35520
rect 154920 35520 155080 35680
rect 154920 35680 155080 35840
rect 154920 35840 155080 36000
rect 154920 36000 155080 36160
rect 154920 36160 155080 36320
rect 154920 36320 155080 36480
rect 154920 36480 155080 36640
rect 154920 36640 155080 36800
rect 154920 36800 155080 36960
rect 154920 36960 155080 37120
rect 154920 37120 155080 37280
rect 154920 37280 155080 37440
rect 154920 37440 155080 37600
rect 154920 37600 155080 37760
rect 154920 37760 155080 37920
rect 154920 37920 155080 38080
rect 154920 38080 155080 38240
rect 154920 38240 155080 38400
rect 154920 38400 155080 38560
rect 154920 38560 155080 38720
rect 154920 38720 155080 38880
rect 154920 38880 155080 39040
rect 154920 39040 155080 39200
rect 154920 39200 155080 39360
rect 154920 39360 155080 39520
rect 154920 39520 155080 39680
rect 154920 39680 155080 39840
rect 154920 39840 155080 40000
rect 154920 40000 155080 40160
rect 154920 40160 155080 40320
rect 154920 40320 155080 40480
rect 154920 40480 155080 40640
rect 154920 40640 155080 40800
rect 154920 40800 155080 40960
rect 154920 40960 155080 41120
rect 154920 41120 155080 41280
rect 154920 41280 155080 41440
rect 154920 41440 155080 41600
rect 154920 41600 155080 41760
rect 154920 41760 155080 41920
rect 154920 41920 155080 42080
rect 154920 42080 155080 42240
rect 154920 42240 155080 42400
rect 154920 42400 155080 42560
rect 154920 42560 155080 42720
rect 154920 42720 155080 42880
rect 154920 42880 155080 43040
rect 154920 43040 155080 43200
rect 154920 43200 155080 43360
rect 154920 43360 155080 43520
rect 154920 43520 155080 43680
rect 154920 43680 155080 43840
rect 155080 34080 155240 34240
rect 155080 34240 155240 34400
rect 155080 34400 155240 34560
rect 155080 34560 155240 34720
rect 155080 34720 155240 34880
rect 155080 34880 155240 35040
rect 155080 35040 155240 35200
rect 155080 35200 155240 35360
rect 155080 35360 155240 35520
rect 155080 35520 155240 35680
rect 155080 35680 155240 35840
rect 155080 35840 155240 36000
rect 155080 36000 155240 36160
rect 155080 36160 155240 36320
rect 155080 36320 155240 36480
rect 155080 36480 155240 36640
rect 155080 36640 155240 36800
rect 155080 36800 155240 36960
rect 155080 36960 155240 37120
rect 155080 37120 155240 37280
rect 155080 37280 155240 37440
rect 155080 37440 155240 37600
rect 155080 37600 155240 37760
rect 155080 37760 155240 37920
rect 155080 37920 155240 38080
rect 155080 38080 155240 38240
rect 155080 38240 155240 38400
rect 155080 38400 155240 38560
rect 155080 38560 155240 38720
rect 155080 38720 155240 38880
rect 155080 38880 155240 39040
rect 155080 39040 155240 39200
rect 155080 39200 155240 39360
rect 155080 39360 155240 39520
rect 155080 39520 155240 39680
rect 155080 39680 155240 39840
rect 155080 39840 155240 40000
rect 155080 40000 155240 40160
rect 155080 40160 155240 40320
rect 155080 40320 155240 40480
rect 155080 40480 155240 40640
rect 155080 40640 155240 40800
rect 155080 40800 155240 40960
rect 155080 40960 155240 41120
rect 155080 41120 155240 41280
rect 155080 41280 155240 41440
rect 155080 41440 155240 41600
rect 155080 41600 155240 41760
rect 155080 41760 155240 41920
rect 155080 41920 155240 42080
rect 155080 42080 155240 42240
rect 155080 42240 155240 42400
rect 155080 42400 155240 42560
rect 155080 42560 155240 42720
rect 155080 42720 155240 42880
rect 155080 42880 155240 43040
rect 155080 43040 155240 43200
rect 155080 43200 155240 43360
rect 155080 43360 155240 43520
rect 155080 43520 155240 43680
rect 155080 43680 155240 43840
rect 155240 33920 155400 34080
rect 155240 34080 155400 34240
rect 155240 34240 155400 34400
rect 155240 34400 155400 34560
rect 155240 34560 155400 34720
rect 155240 34720 155400 34880
rect 155240 34880 155400 35040
rect 155240 35040 155400 35200
rect 155240 35200 155400 35360
rect 155240 35360 155400 35520
rect 155240 35520 155400 35680
rect 155240 35680 155400 35840
rect 155240 35840 155400 36000
rect 155240 36000 155400 36160
rect 155240 36160 155400 36320
rect 155240 36320 155400 36480
rect 155240 36480 155400 36640
rect 155240 36640 155400 36800
rect 155240 36800 155400 36960
rect 155240 36960 155400 37120
rect 155240 37120 155400 37280
rect 155240 37280 155400 37440
rect 155240 37440 155400 37600
rect 155240 37600 155400 37760
rect 155240 37760 155400 37920
rect 155240 37920 155400 38080
rect 155240 38080 155400 38240
rect 155240 38240 155400 38400
rect 155240 38400 155400 38560
rect 155240 38560 155400 38720
rect 155240 38720 155400 38880
rect 155240 38880 155400 39040
rect 155240 39040 155400 39200
rect 155240 39200 155400 39360
rect 155240 39360 155400 39520
rect 155240 39520 155400 39680
rect 155240 39680 155400 39840
rect 155240 39840 155400 40000
rect 155240 40000 155400 40160
rect 155240 40160 155400 40320
rect 155240 40320 155400 40480
rect 155240 40480 155400 40640
rect 155240 40640 155400 40800
rect 155240 40800 155400 40960
rect 155240 40960 155400 41120
rect 155240 41120 155400 41280
rect 155240 41280 155400 41440
rect 155240 41440 155400 41600
rect 155240 41600 155400 41760
rect 155240 41760 155400 41920
rect 155240 41920 155400 42080
rect 155240 42080 155400 42240
rect 155240 42240 155400 42400
rect 155240 42400 155400 42560
rect 155240 42560 155400 42720
rect 155240 42720 155400 42880
rect 155240 42880 155400 43040
rect 155240 43040 155400 43200
rect 155240 43200 155400 43360
rect 155240 43360 155400 43520
rect 155240 43520 155400 43680
rect 155240 43680 155400 43840
rect 155240 43840 155400 44000
rect 155240 44000 155400 44160
rect 155400 33760 155560 33920
rect 155400 33920 155560 34080
rect 155400 34080 155560 34240
rect 155400 34240 155560 34400
rect 155400 34400 155560 34560
rect 155400 34560 155560 34720
rect 155400 34720 155560 34880
rect 155400 34880 155560 35040
rect 155400 35040 155560 35200
rect 155400 35200 155560 35360
rect 155400 35360 155560 35520
rect 155400 35520 155560 35680
rect 155400 35680 155560 35840
rect 155400 35840 155560 36000
rect 155400 36000 155560 36160
rect 155400 36160 155560 36320
rect 155400 36320 155560 36480
rect 155400 36480 155560 36640
rect 155400 36640 155560 36800
rect 155400 36800 155560 36960
rect 155400 36960 155560 37120
rect 155400 37120 155560 37280
rect 155400 37280 155560 37440
rect 155400 37440 155560 37600
rect 155400 37600 155560 37760
rect 155400 37760 155560 37920
rect 155400 37920 155560 38080
rect 155400 38080 155560 38240
rect 155400 38240 155560 38400
rect 155400 38400 155560 38560
rect 155400 38560 155560 38720
rect 155400 38720 155560 38880
rect 155400 38880 155560 39040
rect 155400 39040 155560 39200
rect 155400 39200 155560 39360
rect 155400 39360 155560 39520
rect 155400 39520 155560 39680
rect 155400 39680 155560 39840
rect 155400 39840 155560 40000
rect 155400 40000 155560 40160
rect 155400 40160 155560 40320
rect 155400 40320 155560 40480
rect 155400 40480 155560 40640
rect 155400 40640 155560 40800
rect 155400 40800 155560 40960
rect 155400 40960 155560 41120
rect 155400 41120 155560 41280
rect 155400 41280 155560 41440
rect 155400 41440 155560 41600
rect 155400 41600 155560 41760
rect 155400 41760 155560 41920
rect 155400 41920 155560 42080
rect 155400 42080 155560 42240
rect 155400 42240 155560 42400
rect 155400 42400 155560 42560
rect 155400 42560 155560 42720
rect 155400 42720 155560 42880
rect 155400 42880 155560 43040
rect 155400 43040 155560 43200
rect 155400 43200 155560 43360
rect 155400 43360 155560 43520
rect 155400 43520 155560 43680
rect 155400 43680 155560 43840
rect 155400 43840 155560 44000
rect 155400 44000 155560 44160
rect 155400 44160 155560 44320
rect 155560 33600 155720 33760
rect 155560 33760 155720 33920
rect 155560 33920 155720 34080
rect 155560 34080 155720 34240
rect 155560 34240 155720 34400
rect 155560 34400 155720 34560
rect 155560 34560 155720 34720
rect 155560 34720 155720 34880
rect 155560 34880 155720 35040
rect 155560 35040 155720 35200
rect 155560 35200 155720 35360
rect 155560 35360 155720 35520
rect 155560 35520 155720 35680
rect 155560 35680 155720 35840
rect 155560 35840 155720 36000
rect 155560 36000 155720 36160
rect 155560 36160 155720 36320
rect 155560 36320 155720 36480
rect 155560 36480 155720 36640
rect 155560 36640 155720 36800
rect 155560 36800 155720 36960
rect 155560 36960 155720 37120
rect 155560 37120 155720 37280
rect 155560 37280 155720 37440
rect 155560 37440 155720 37600
rect 155560 37600 155720 37760
rect 155560 37760 155720 37920
rect 155560 37920 155720 38080
rect 155560 38080 155720 38240
rect 155560 38240 155720 38400
rect 155560 38400 155720 38560
rect 155560 38560 155720 38720
rect 155560 38720 155720 38880
rect 155560 38880 155720 39040
rect 155560 39040 155720 39200
rect 155560 39200 155720 39360
rect 155560 39360 155720 39520
rect 155560 39520 155720 39680
rect 155560 39680 155720 39840
rect 155560 39840 155720 40000
rect 155560 40000 155720 40160
rect 155560 40160 155720 40320
rect 155560 40320 155720 40480
rect 155560 40480 155720 40640
rect 155560 40640 155720 40800
rect 155560 40800 155720 40960
rect 155560 40960 155720 41120
rect 155560 41120 155720 41280
rect 155560 41280 155720 41440
rect 155560 41440 155720 41600
rect 155560 41600 155720 41760
rect 155560 41760 155720 41920
rect 155560 41920 155720 42080
rect 155560 42080 155720 42240
rect 155560 42240 155720 42400
rect 155560 42400 155720 42560
rect 155560 42560 155720 42720
rect 155560 42720 155720 42880
rect 155560 42880 155720 43040
rect 155560 43040 155720 43200
rect 155560 43200 155720 43360
rect 155560 43360 155720 43520
rect 155560 43520 155720 43680
rect 155560 43680 155720 43840
rect 155560 43840 155720 44000
rect 155560 44000 155720 44160
rect 155560 44160 155720 44320
rect 155560 44320 155720 44480
rect 155720 33440 155880 33600
rect 155720 33600 155880 33760
rect 155720 33760 155880 33920
rect 155720 33920 155880 34080
rect 155720 34080 155880 34240
rect 155720 34240 155880 34400
rect 155720 34400 155880 34560
rect 155720 34560 155880 34720
rect 155720 34720 155880 34880
rect 155720 34880 155880 35040
rect 155720 35040 155880 35200
rect 155720 35200 155880 35360
rect 155720 35360 155880 35520
rect 155720 35520 155880 35680
rect 155720 35680 155880 35840
rect 155720 35840 155880 36000
rect 155720 36000 155880 36160
rect 155720 36160 155880 36320
rect 155720 36320 155880 36480
rect 155720 36480 155880 36640
rect 155720 36640 155880 36800
rect 155720 36800 155880 36960
rect 155720 36960 155880 37120
rect 155720 37120 155880 37280
rect 155720 37280 155880 37440
rect 155720 37440 155880 37600
rect 155720 37600 155880 37760
rect 155720 37760 155880 37920
rect 155720 37920 155880 38080
rect 155720 38080 155880 38240
rect 155720 38240 155880 38400
rect 155720 38400 155880 38560
rect 155720 38560 155880 38720
rect 155720 38720 155880 38880
rect 155720 38880 155880 39040
rect 155720 39040 155880 39200
rect 155720 39200 155880 39360
rect 155720 39360 155880 39520
rect 155720 39520 155880 39680
rect 155720 39680 155880 39840
rect 155720 39840 155880 40000
rect 155720 40000 155880 40160
rect 155720 40160 155880 40320
rect 155720 40320 155880 40480
rect 155720 40480 155880 40640
rect 155720 40640 155880 40800
rect 155720 40800 155880 40960
rect 155720 40960 155880 41120
rect 155720 41120 155880 41280
rect 155720 41280 155880 41440
rect 155720 41440 155880 41600
rect 155720 41600 155880 41760
rect 155720 41760 155880 41920
rect 155720 41920 155880 42080
rect 155720 42080 155880 42240
rect 155720 42240 155880 42400
rect 155720 42400 155880 42560
rect 155720 42560 155880 42720
rect 155720 42720 155880 42880
rect 155720 42880 155880 43040
rect 155720 43040 155880 43200
rect 155720 43200 155880 43360
rect 155720 43360 155880 43520
rect 155720 43520 155880 43680
rect 155720 43680 155880 43840
rect 155720 43840 155880 44000
rect 155720 44000 155880 44160
rect 155720 44160 155880 44320
rect 155720 44320 155880 44480
rect 155720 44480 155880 44640
rect 155880 33280 156040 33440
rect 155880 33440 156040 33600
rect 155880 33600 156040 33760
rect 155880 33760 156040 33920
rect 155880 33920 156040 34080
rect 155880 34080 156040 34240
rect 155880 34240 156040 34400
rect 155880 34400 156040 34560
rect 155880 34560 156040 34720
rect 155880 34720 156040 34880
rect 155880 34880 156040 35040
rect 155880 35040 156040 35200
rect 155880 35200 156040 35360
rect 155880 35360 156040 35520
rect 155880 35520 156040 35680
rect 155880 35680 156040 35840
rect 155880 35840 156040 36000
rect 155880 36000 156040 36160
rect 155880 36160 156040 36320
rect 155880 36320 156040 36480
rect 155880 36480 156040 36640
rect 155880 36640 156040 36800
rect 155880 36800 156040 36960
rect 155880 36960 156040 37120
rect 155880 37120 156040 37280
rect 155880 37280 156040 37440
rect 155880 37440 156040 37600
rect 155880 37600 156040 37760
rect 155880 37760 156040 37920
rect 155880 37920 156040 38080
rect 155880 38080 156040 38240
rect 155880 38240 156040 38400
rect 155880 38400 156040 38560
rect 155880 38560 156040 38720
rect 155880 38720 156040 38880
rect 155880 38880 156040 39040
rect 155880 39040 156040 39200
rect 155880 39200 156040 39360
rect 155880 39360 156040 39520
rect 155880 39520 156040 39680
rect 155880 39680 156040 39840
rect 155880 39840 156040 40000
rect 155880 40000 156040 40160
rect 155880 40160 156040 40320
rect 155880 40320 156040 40480
rect 155880 40480 156040 40640
rect 155880 40640 156040 40800
rect 155880 40800 156040 40960
rect 155880 40960 156040 41120
rect 155880 41120 156040 41280
rect 155880 41280 156040 41440
rect 155880 41440 156040 41600
rect 155880 41600 156040 41760
rect 155880 41760 156040 41920
rect 155880 41920 156040 42080
rect 155880 42080 156040 42240
rect 155880 42240 156040 42400
rect 155880 42400 156040 42560
rect 155880 42560 156040 42720
rect 155880 42720 156040 42880
rect 155880 42880 156040 43040
rect 155880 43040 156040 43200
rect 155880 43200 156040 43360
rect 155880 43360 156040 43520
rect 155880 43520 156040 43680
rect 155880 43680 156040 43840
rect 155880 43840 156040 44000
rect 155880 44000 156040 44160
rect 155880 44160 156040 44320
rect 155880 44320 156040 44480
rect 155880 44480 156040 44640
rect 155880 44640 156040 44800
rect 156040 33120 156200 33280
rect 156040 33280 156200 33440
rect 156040 33440 156200 33600
rect 156040 33600 156200 33760
rect 156040 33760 156200 33920
rect 156040 33920 156200 34080
rect 156040 34080 156200 34240
rect 156040 34240 156200 34400
rect 156040 34400 156200 34560
rect 156040 34560 156200 34720
rect 156040 34720 156200 34880
rect 156040 34880 156200 35040
rect 156040 35040 156200 35200
rect 156040 35200 156200 35360
rect 156040 35360 156200 35520
rect 156040 35520 156200 35680
rect 156040 35680 156200 35840
rect 156040 35840 156200 36000
rect 156040 36000 156200 36160
rect 156040 36160 156200 36320
rect 156040 36320 156200 36480
rect 156040 36480 156200 36640
rect 156040 36640 156200 36800
rect 156040 36800 156200 36960
rect 156040 36960 156200 37120
rect 156040 37120 156200 37280
rect 156040 37280 156200 37440
rect 156040 37440 156200 37600
rect 156040 37600 156200 37760
rect 156040 37760 156200 37920
rect 156040 37920 156200 38080
rect 156040 38080 156200 38240
rect 156040 38240 156200 38400
rect 156040 38400 156200 38560
rect 156040 38560 156200 38720
rect 156040 38720 156200 38880
rect 156040 38880 156200 39040
rect 156040 39040 156200 39200
rect 156040 39200 156200 39360
rect 156040 39360 156200 39520
rect 156040 39520 156200 39680
rect 156040 39680 156200 39840
rect 156040 39840 156200 40000
rect 156040 40000 156200 40160
rect 156040 40160 156200 40320
rect 156040 40320 156200 40480
rect 156040 40480 156200 40640
rect 156040 40640 156200 40800
rect 156040 40800 156200 40960
rect 156040 40960 156200 41120
rect 156040 41120 156200 41280
rect 156040 41280 156200 41440
rect 156040 41440 156200 41600
rect 156040 41600 156200 41760
rect 156040 41760 156200 41920
rect 156040 41920 156200 42080
rect 156040 42080 156200 42240
rect 156040 42240 156200 42400
rect 156040 42400 156200 42560
rect 156040 42560 156200 42720
rect 156040 42720 156200 42880
rect 156040 42880 156200 43040
rect 156040 43040 156200 43200
rect 156040 43200 156200 43360
rect 156040 43360 156200 43520
rect 156040 43520 156200 43680
rect 156040 43680 156200 43840
rect 156040 43840 156200 44000
rect 156040 44000 156200 44160
rect 156040 44160 156200 44320
rect 156040 44320 156200 44480
rect 156040 44480 156200 44640
rect 156040 44640 156200 44800
rect 156040 44800 156200 44960
rect 156200 32960 156360 33120
rect 156200 33120 156360 33280
rect 156200 33280 156360 33440
rect 156200 33440 156360 33600
rect 156200 33600 156360 33760
rect 156200 33760 156360 33920
rect 156200 33920 156360 34080
rect 156200 34080 156360 34240
rect 156200 34240 156360 34400
rect 156200 34400 156360 34560
rect 156200 34560 156360 34720
rect 156200 34720 156360 34880
rect 156200 34880 156360 35040
rect 156200 35040 156360 35200
rect 156200 35200 156360 35360
rect 156200 35360 156360 35520
rect 156200 35520 156360 35680
rect 156200 35680 156360 35840
rect 156200 35840 156360 36000
rect 156200 36000 156360 36160
rect 156200 36160 156360 36320
rect 156200 36320 156360 36480
rect 156200 36480 156360 36640
rect 156200 36640 156360 36800
rect 156200 36800 156360 36960
rect 156200 36960 156360 37120
rect 156200 37120 156360 37280
rect 156200 37280 156360 37440
rect 156200 37440 156360 37600
rect 156200 37600 156360 37760
rect 156200 37760 156360 37920
rect 156200 38080 156360 38240
rect 156200 38240 156360 38400
rect 156200 38400 156360 38560
rect 156200 38560 156360 38720
rect 156200 38720 156360 38880
rect 156200 38880 156360 39040
rect 156200 39040 156360 39200
rect 156200 39200 156360 39360
rect 156200 39360 156360 39520
rect 156200 39520 156360 39680
rect 156200 39680 156360 39840
rect 156200 39840 156360 40000
rect 156200 40000 156360 40160
rect 156200 40320 156360 40480
rect 156200 40480 156360 40640
rect 156200 40640 156360 40800
rect 156200 40800 156360 40960
rect 156200 40960 156360 41120
rect 156200 41120 156360 41280
rect 156200 41280 156360 41440
rect 156200 41440 156360 41600
rect 156200 41600 156360 41760
rect 156200 41760 156360 41920
rect 156200 41920 156360 42080
rect 156200 42080 156360 42240
rect 156200 42240 156360 42400
rect 156200 42400 156360 42560
rect 156200 42560 156360 42720
rect 156200 42720 156360 42880
rect 156200 42880 156360 43040
rect 156200 43040 156360 43200
rect 156200 43200 156360 43360
rect 156200 43360 156360 43520
rect 156200 43520 156360 43680
rect 156200 43680 156360 43840
rect 156200 43840 156360 44000
rect 156200 44000 156360 44160
rect 156200 44160 156360 44320
rect 156200 44320 156360 44480
rect 156200 44480 156360 44640
rect 156200 44640 156360 44800
rect 156200 44800 156360 44960
rect 156200 44960 156360 45120
rect 156360 32800 156520 32960
rect 156360 32960 156520 33120
rect 156360 33120 156520 33280
rect 156360 33280 156520 33440
rect 156360 33440 156520 33600
rect 156360 33600 156520 33760
rect 156360 33760 156520 33920
rect 156360 33920 156520 34080
rect 156360 34080 156520 34240
rect 156360 34240 156520 34400
rect 156360 34400 156520 34560
rect 156360 34560 156520 34720
rect 156360 34720 156520 34880
rect 156360 34880 156520 35040
rect 156360 35040 156520 35200
rect 156360 35200 156520 35360
rect 156360 35360 156520 35520
rect 156360 35520 156520 35680
rect 156360 35680 156520 35840
rect 156360 35840 156520 36000
rect 156360 36000 156520 36160
rect 156360 36160 156520 36320
rect 156360 36320 156520 36480
rect 156360 36480 156520 36640
rect 156360 36640 156520 36800
rect 156360 36800 156520 36960
rect 156360 36960 156520 37120
rect 156360 37120 156520 37280
rect 156360 37280 156520 37440
rect 156360 37440 156520 37600
rect 156360 37600 156520 37760
rect 156360 40480 156520 40640
rect 156360 40640 156520 40800
rect 156360 40800 156520 40960
rect 156360 40960 156520 41120
rect 156360 41120 156520 41280
rect 156360 41280 156520 41440
rect 156360 41440 156520 41600
rect 156360 41600 156520 41760
rect 156360 41760 156520 41920
rect 156360 41920 156520 42080
rect 156360 42080 156520 42240
rect 156360 42240 156520 42400
rect 156360 42400 156520 42560
rect 156360 42560 156520 42720
rect 156360 42720 156520 42880
rect 156360 42880 156520 43040
rect 156360 43040 156520 43200
rect 156360 43200 156520 43360
rect 156360 43360 156520 43520
rect 156360 43520 156520 43680
rect 156360 43680 156520 43840
rect 156360 43840 156520 44000
rect 156360 44000 156520 44160
rect 156360 44160 156520 44320
rect 156360 44320 156520 44480
rect 156360 44480 156520 44640
rect 156360 44640 156520 44800
rect 156360 44800 156520 44960
rect 156360 44960 156520 45120
rect 156360 45120 156520 45280
rect 156520 32640 156680 32800
rect 156520 32800 156680 32960
rect 156520 32960 156680 33120
rect 156520 33120 156680 33280
rect 156520 33280 156680 33440
rect 156520 33440 156680 33600
rect 156520 33600 156680 33760
rect 156520 33760 156680 33920
rect 156520 33920 156680 34080
rect 156520 34080 156680 34240
rect 156520 34240 156680 34400
rect 156520 34400 156680 34560
rect 156520 34560 156680 34720
rect 156520 34720 156680 34880
rect 156520 34880 156680 35040
rect 156520 35040 156680 35200
rect 156520 35200 156680 35360
rect 156520 35360 156680 35520
rect 156520 35520 156680 35680
rect 156520 35680 156680 35840
rect 156520 35840 156680 36000
rect 156520 36000 156680 36160
rect 156520 36160 156680 36320
rect 156520 36320 156680 36480
rect 156520 36480 156680 36640
rect 156520 36640 156680 36800
rect 156520 36800 156680 36960
rect 156520 36960 156680 37120
rect 156520 37120 156680 37280
rect 156520 37280 156680 37440
rect 156520 37440 156680 37600
rect 156520 40640 156680 40800
rect 156520 40800 156680 40960
rect 156520 40960 156680 41120
rect 156520 41120 156680 41280
rect 156520 41280 156680 41440
rect 156520 41440 156680 41600
rect 156520 41600 156680 41760
rect 156520 41760 156680 41920
rect 156520 41920 156680 42080
rect 156520 42080 156680 42240
rect 156520 42240 156680 42400
rect 156520 42400 156680 42560
rect 156520 42560 156680 42720
rect 156520 42720 156680 42880
rect 156520 42880 156680 43040
rect 156520 43040 156680 43200
rect 156520 43200 156680 43360
rect 156520 43360 156680 43520
rect 156520 43520 156680 43680
rect 156520 43680 156680 43840
rect 156520 43840 156680 44000
rect 156520 44000 156680 44160
rect 156520 44160 156680 44320
rect 156520 44320 156680 44480
rect 156520 44480 156680 44640
rect 156520 44640 156680 44800
rect 156520 44800 156680 44960
rect 156520 44960 156680 45120
rect 156520 45120 156680 45280
rect 156520 45280 156680 45440
rect 156680 32480 156840 32640
rect 156680 32640 156840 32800
rect 156680 32800 156840 32960
rect 156680 32960 156840 33120
rect 156680 33120 156840 33280
rect 156680 33280 156840 33440
rect 156680 33440 156840 33600
rect 156680 33600 156840 33760
rect 156680 33760 156840 33920
rect 156680 33920 156840 34080
rect 156680 34080 156840 34240
rect 156680 34240 156840 34400
rect 156680 34400 156840 34560
rect 156680 34560 156840 34720
rect 156680 34720 156840 34880
rect 156680 34880 156840 35040
rect 156680 35040 156840 35200
rect 156680 35200 156840 35360
rect 156680 35360 156840 35520
rect 156680 35520 156840 35680
rect 156680 35680 156840 35840
rect 156680 35840 156840 36000
rect 156680 36000 156840 36160
rect 156680 36160 156840 36320
rect 156680 36320 156840 36480
rect 156680 36480 156840 36640
rect 156680 36640 156840 36800
rect 156680 36800 156840 36960
rect 156680 36960 156840 37120
rect 156680 37120 156840 37280
rect 156680 37280 156840 37440
rect 156680 40800 156840 40960
rect 156680 40960 156840 41120
rect 156680 41120 156840 41280
rect 156680 41280 156840 41440
rect 156680 41440 156840 41600
rect 156680 41600 156840 41760
rect 156680 41760 156840 41920
rect 156680 41920 156840 42080
rect 156680 42080 156840 42240
rect 156680 42240 156840 42400
rect 156680 42400 156840 42560
rect 156680 42560 156840 42720
rect 156680 42720 156840 42880
rect 156680 42880 156840 43040
rect 156680 43040 156840 43200
rect 156680 43200 156840 43360
rect 156680 43360 156840 43520
rect 156680 43520 156840 43680
rect 156680 43680 156840 43840
rect 156680 43840 156840 44000
rect 156680 44000 156840 44160
rect 156680 44160 156840 44320
rect 156680 44320 156840 44480
rect 156680 44480 156840 44640
rect 156680 44640 156840 44800
rect 156680 44800 156840 44960
rect 156680 44960 156840 45120
rect 156680 45120 156840 45280
rect 156680 45280 156840 45440
rect 156680 45440 156840 45600
rect 156840 32320 157000 32480
rect 156840 32480 157000 32640
rect 156840 32640 157000 32800
rect 156840 32800 157000 32960
rect 156840 32960 157000 33120
rect 156840 33120 157000 33280
rect 156840 33280 157000 33440
rect 156840 33440 157000 33600
rect 156840 33600 157000 33760
rect 156840 33760 157000 33920
rect 156840 33920 157000 34080
rect 156840 34080 157000 34240
rect 156840 34240 157000 34400
rect 156840 34400 157000 34560
rect 156840 34560 157000 34720
rect 156840 34720 157000 34880
rect 156840 34880 157000 35040
rect 156840 35040 157000 35200
rect 156840 35200 157000 35360
rect 156840 35360 157000 35520
rect 156840 35520 157000 35680
rect 156840 35680 157000 35840
rect 156840 35840 157000 36000
rect 156840 36000 157000 36160
rect 156840 36160 157000 36320
rect 156840 36320 157000 36480
rect 156840 36480 157000 36640
rect 156840 36640 157000 36800
rect 156840 36800 157000 36960
rect 156840 36960 157000 37120
rect 156840 37120 157000 37280
rect 156840 40960 157000 41120
rect 156840 41120 157000 41280
rect 156840 41280 157000 41440
rect 156840 41440 157000 41600
rect 156840 41600 157000 41760
rect 156840 41760 157000 41920
rect 156840 41920 157000 42080
rect 156840 42080 157000 42240
rect 156840 42240 157000 42400
rect 156840 42400 157000 42560
rect 156840 42560 157000 42720
rect 156840 42720 157000 42880
rect 156840 42880 157000 43040
rect 156840 43040 157000 43200
rect 156840 43200 157000 43360
rect 156840 43360 157000 43520
rect 156840 43520 157000 43680
rect 156840 43680 157000 43840
rect 156840 43840 157000 44000
rect 156840 44000 157000 44160
rect 156840 44160 157000 44320
rect 156840 44320 157000 44480
rect 156840 44480 157000 44640
rect 156840 44640 157000 44800
rect 156840 44800 157000 44960
rect 156840 44960 157000 45120
rect 156840 45120 157000 45280
rect 156840 45280 157000 45440
rect 156840 45440 157000 45600
rect 156840 45600 157000 45760
rect 157000 32160 157160 32320
rect 157000 32320 157160 32480
rect 157000 32480 157160 32640
rect 157000 32640 157160 32800
rect 157000 32800 157160 32960
rect 157000 32960 157160 33120
rect 157000 33120 157160 33280
rect 157000 33280 157160 33440
rect 157000 33440 157160 33600
rect 157000 33600 157160 33760
rect 157000 33760 157160 33920
rect 157000 33920 157160 34080
rect 157000 34080 157160 34240
rect 157000 34240 157160 34400
rect 157000 34400 157160 34560
rect 157000 34560 157160 34720
rect 157000 34720 157160 34880
rect 157000 34880 157160 35040
rect 157000 35040 157160 35200
rect 157000 35200 157160 35360
rect 157000 35360 157160 35520
rect 157000 35520 157160 35680
rect 157000 35680 157160 35840
rect 157000 35840 157160 36000
rect 157000 36000 157160 36160
rect 157000 36160 157160 36320
rect 157000 36320 157160 36480
rect 157000 36480 157160 36640
rect 157000 36640 157160 36800
rect 157000 36800 157160 36960
rect 157000 36960 157160 37120
rect 157000 41120 157160 41280
rect 157000 41280 157160 41440
rect 157000 41440 157160 41600
rect 157000 41600 157160 41760
rect 157000 41760 157160 41920
rect 157000 41920 157160 42080
rect 157000 42080 157160 42240
rect 157000 42240 157160 42400
rect 157000 42400 157160 42560
rect 157000 42560 157160 42720
rect 157000 42720 157160 42880
rect 157000 42880 157160 43040
rect 157000 43040 157160 43200
rect 157000 43200 157160 43360
rect 157000 43360 157160 43520
rect 157000 43520 157160 43680
rect 157000 43680 157160 43840
rect 157000 43840 157160 44000
rect 157000 44000 157160 44160
rect 157000 44160 157160 44320
rect 157000 44320 157160 44480
rect 157000 44480 157160 44640
rect 157000 44640 157160 44800
rect 157000 44800 157160 44960
rect 157000 44960 157160 45120
rect 157000 45120 157160 45280
rect 157000 45280 157160 45440
rect 157000 45440 157160 45600
rect 157000 45600 157160 45760
rect 157000 45760 157160 45920
rect 157000 45920 157160 46080
rect 157160 32000 157320 32160
rect 157160 32160 157320 32320
rect 157160 32320 157320 32480
rect 157160 32480 157320 32640
rect 157160 32640 157320 32800
rect 157160 32800 157320 32960
rect 157160 32960 157320 33120
rect 157160 33120 157320 33280
rect 157160 33280 157320 33440
rect 157160 33440 157320 33600
rect 157160 33600 157320 33760
rect 157160 33760 157320 33920
rect 157160 33920 157320 34080
rect 157160 34080 157320 34240
rect 157160 34240 157320 34400
rect 157160 34400 157320 34560
rect 157160 34560 157320 34720
rect 157160 34720 157320 34880
rect 157160 34880 157320 35040
rect 157160 35040 157320 35200
rect 157160 35200 157320 35360
rect 157160 35360 157320 35520
rect 157160 35520 157320 35680
rect 157160 35680 157320 35840
rect 157160 35840 157320 36000
rect 157160 36000 157320 36160
rect 157160 36160 157320 36320
rect 157160 36320 157320 36480
rect 157160 36480 157320 36640
rect 157160 36640 157320 36800
rect 157160 36800 157320 36960
rect 157160 41280 157320 41440
rect 157160 41440 157320 41600
rect 157160 41600 157320 41760
rect 157160 41760 157320 41920
rect 157160 41920 157320 42080
rect 157160 42080 157320 42240
rect 157160 42240 157320 42400
rect 157160 42400 157320 42560
rect 157160 42560 157320 42720
rect 157160 42720 157320 42880
rect 157160 42880 157320 43040
rect 157160 43040 157320 43200
rect 157160 43200 157320 43360
rect 157160 43360 157320 43520
rect 157160 43520 157320 43680
rect 157160 43680 157320 43840
rect 157160 43840 157320 44000
rect 157160 44000 157320 44160
rect 157160 44160 157320 44320
rect 157160 44320 157320 44480
rect 157160 44480 157320 44640
rect 157160 44640 157320 44800
rect 157160 44800 157320 44960
rect 157160 44960 157320 45120
rect 157160 45120 157320 45280
rect 157160 45280 157320 45440
rect 157160 45440 157320 45600
rect 157160 45600 157320 45760
rect 157160 45760 157320 45920
rect 157160 45920 157320 46080
rect 157160 46080 157320 46240
rect 157320 31840 157480 32000
rect 157320 32000 157480 32160
rect 157320 32160 157480 32320
rect 157320 32320 157480 32480
rect 157320 32480 157480 32640
rect 157320 32640 157480 32800
rect 157320 32800 157480 32960
rect 157320 32960 157480 33120
rect 157320 33120 157480 33280
rect 157320 33280 157480 33440
rect 157320 33440 157480 33600
rect 157320 33600 157480 33760
rect 157320 33760 157480 33920
rect 157320 33920 157480 34080
rect 157320 34080 157480 34240
rect 157320 34240 157480 34400
rect 157320 34400 157480 34560
rect 157320 34560 157480 34720
rect 157320 34720 157480 34880
rect 157320 34880 157480 35040
rect 157320 35040 157480 35200
rect 157320 35200 157480 35360
rect 157320 35360 157480 35520
rect 157320 35520 157480 35680
rect 157320 35680 157480 35840
rect 157320 35840 157480 36000
rect 157320 36000 157480 36160
rect 157320 36160 157480 36320
rect 157320 36320 157480 36480
rect 157320 36480 157480 36640
rect 157320 36640 157480 36800
rect 157320 41440 157480 41600
rect 157320 41600 157480 41760
rect 157320 41760 157480 41920
rect 157320 41920 157480 42080
rect 157320 42080 157480 42240
rect 157320 42240 157480 42400
rect 157320 42400 157480 42560
rect 157320 42560 157480 42720
rect 157320 42720 157480 42880
rect 157320 42880 157480 43040
rect 157320 43040 157480 43200
rect 157320 43200 157480 43360
rect 157320 43360 157480 43520
rect 157320 43520 157480 43680
rect 157320 43680 157480 43840
rect 157320 43840 157480 44000
rect 157320 44000 157480 44160
rect 157320 44160 157480 44320
rect 157320 44320 157480 44480
rect 157320 44480 157480 44640
rect 157320 44640 157480 44800
rect 157320 44800 157480 44960
rect 157320 44960 157480 45120
rect 157320 45120 157480 45280
rect 157320 45280 157480 45440
rect 157320 45440 157480 45600
rect 157320 45600 157480 45760
rect 157320 45760 157480 45920
rect 157320 45920 157480 46080
rect 157320 46080 157480 46240
rect 157320 46240 157480 46400
rect 157480 31680 157640 31840
rect 157480 31840 157640 32000
rect 157480 32000 157640 32160
rect 157480 32160 157640 32320
rect 157480 32320 157640 32480
rect 157480 32480 157640 32640
rect 157480 32640 157640 32800
rect 157480 32800 157640 32960
rect 157480 32960 157640 33120
rect 157480 33120 157640 33280
rect 157480 33280 157640 33440
rect 157480 33440 157640 33600
rect 157480 33600 157640 33760
rect 157480 33760 157640 33920
rect 157480 33920 157640 34080
rect 157480 34080 157640 34240
rect 157480 34240 157640 34400
rect 157480 34400 157640 34560
rect 157480 34560 157640 34720
rect 157480 34720 157640 34880
rect 157480 34880 157640 35040
rect 157480 35040 157640 35200
rect 157480 35200 157640 35360
rect 157480 35360 157640 35520
rect 157480 35520 157640 35680
rect 157480 35680 157640 35840
rect 157480 35840 157640 36000
rect 157480 36000 157640 36160
rect 157480 36160 157640 36320
rect 157480 36320 157640 36480
rect 157480 36480 157640 36640
rect 157480 41600 157640 41760
rect 157480 41760 157640 41920
rect 157480 41920 157640 42080
rect 157480 42080 157640 42240
rect 157480 42240 157640 42400
rect 157480 42400 157640 42560
rect 157480 42560 157640 42720
rect 157480 42720 157640 42880
rect 157480 42880 157640 43040
rect 157480 43040 157640 43200
rect 157480 43200 157640 43360
rect 157480 43360 157640 43520
rect 157480 43520 157640 43680
rect 157480 43680 157640 43840
rect 157480 43840 157640 44000
rect 157480 44000 157640 44160
rect 157480 44160 157640 44320
rect 157480 44320 157640 44480
rect 157480 44480 157640 44640
rect 157480 44640 157640 44800
rect 157480 44800 157640 44960
rect 157480 44960 157640 45120
rect 157480 45120 157640 45280
rect 157480 45280 157640 45440
rect 157480 45440 157640 45600
rect 157480 45600 157640 45760
rect 157480 45760 157640 45920
rect 157480 45920 157640 46080
rect 157480 46080 157640 46240
rect 157480 46240 157640 46400
rect 157480 46400 157640 46560
rect 157640 31520 157800 31680
rect 157640 31680 157800 31840
rect 157640 31840 157800 32000
rect 157640 32000 157800 32160
rect 157640 32160 157800 32320
rect 157640 32320 157800 32480
rect 157640 32480 157800 32640
rect 157640 32640 157800 32800
rect 157640 32800 157800 32960
rect 157640 32960 157800 33120
rect 157640 33120 157800 33280
rect 157640 33280 157800 33440
rect 157640 33440 157800 33600
rect 157640 33600 157800 33760
rect 157640 33760 157800 33920
rect 157640 33920 157800 34080
rect 157640 34080 157800 34240
rect 157640 34240 157800 34400
rect 157640 34400 157800 34560
rect 157640 34560 157800 34720
rect 157640 34720 157800 34880
rect 157640 34880 157800 35040
rect 157640 35040 157800 35200
rect 157640 35200 157800 35360
rect 157640 35360 157800 35520
rect 157640 35520 157800 35680
rect 157640 35680 157800 35840
rect 157640 35840 157800 36000
rect 157640 36000 157800 36160
rect 157640 36160 157800 36320
rect 157640 36320 157800 36480
rect 157640 41760 157800 41920
rect 157640 41920 157800 42080
rect 157640 42080 157800 42240
rect 157640 42240 157800 42400
rect 157640 42400 157800 42560
rect 157640 42560 157800 42720
rect 157640 42720 157800 42880
rect 157640 42880 157800 43040
rect 157640 43040 157800 43200
rect 157640 43200 157800 43360
rect 157640 43360 157800 43520
rect 157640 43520 157800 43680
rect 157640 43680 157800 43840
rect 157640 43840 157800 44000
rect 157640 44000 157800 44160
rect 157640 44160 157800 44320
rect 157640 44320 157800 44480
rect 157640 44480 157800 44640
rect 157640 44640 157800 44800
rect 157640 44800 157800 44960
rect 157640 44960 157800 45120
rect 157640 45120 157800 45280
rect 157640 45280 157800 45440
rect 157640 45440 157800 45600
rect 157640 45600 157800 45760
rect 157640 45760 157800 45920
rect 157640 45920 157800 46080
rect 157640 46080 157800 46240
rect 157640 46240 157800 46400
rect 157640 46400 157800 46560
rect 157640 46560 157800 46720
rect 157800 31360 157960 31520
rect 157800 31520 157960 31680
rect 157800 31680 157960 31840
rect 157800 31840 157960 32000
rect 157800 32000 157960 32160
rect 157800 32160 157960 32320
rect 157800 32320 157960 32480
rect 157800 32480 157960 32640
rect 157800 32640 157960 32800
rect 157800 32800 157960 32960
rect 157800 32960 157960 33120
rect 157800 33120 157960 33280
rect 157800 33280 157960 33440
rect 157800 33440 157960 33600
rect 157800 33600 157960 33760
rect 157800 33760 157960 33920
rect 157800 33920 157960 34080
rect 157800 34080 157960 34240
rect 157800 34240 157960 34400
rect 157800 34400 157960 34560
rect 157800 34560 157960 34720
rect 157800 34720 157960 34880
rect 157800 34880 157960 35040
rect 157800 35040 157960 35200
rect 157800 35200 157960 35360
rect 157800 35360 157960 35520
rect 157800 35520 157960 35680
rect 157800 35680 157960 35840
rect 157800 35840 157960 36000
rect 157800 36000 157960 36160
rect 157800 36160 157960 36320
rect 157800 41920 157960 42080
rect 157800 42080 157960 42240
rect 157800 42240 157960 42400
rect 157800 42400 157960 42560
rect 157800 42560 157960 42720
rect 157800 42720 157960 42880
rect 157800 42880 157960 43040
rect 157800 43040 157960 43200
rect 157800 43200 157960 43360
rect 157800 43360 157960 43520
rect 157800 43520 157960 43680
rect 157800 43680 157960 43840
rect 157800 43840 157960 44000
rect 157800 44000 157960 44160
rect 157800 44160 157960 44320
rect 157800 44320 157960 44480
rect 157800 44480 157960 44640
rect 157800 44640 157960 44800
rect 157800 44800 157960 44960
rect 157800 44960 157960 45120
rect 157800 45120 157960 45280
rect 157800 45280 157960 45440
rect 157800 45440 157960 45600
rect 157800 45600 157960 45760
rect 157800 45760 157960 45920
rect 157800 45920 157960 46080
rect 157800 46080 157960 46240
rect 157800 46240 157960 46400
rect 157800 46400 157960 46560
rect 157800 46560 157960 46720
rect 157800 46720 157960 46880
rect 157960 31200 158120 31360
rect 157960 31360 158120 31520
rect 157960 31520 158120 31680
rect 157960 31680 158120 31840
rect 157960 31840 158120 32000
rect 157960 32000 158120 32160
rect 157960 32160 158120 32320
rect 157960 32320 158120 32480
rect 157960 32480 158120 32640
rect 157960 32640 158120 32800
rect 157960 32800 158120 32960
rect 157960 32960 158120 33120
rect 157960 33120 158120 33280
rect 157960 33280 158120 33440
rect 157960 33440 158120 33600
rect 157960 33600 158120 33760
rect 157960 33760 158120 33920
rect 157960 33920 158120 34080
rect 157960 34080 158120 34240
rect 157960 34240 158120 34400
rect 157960 34400 158120 34560
rect 157960 34560 158120 34720
rect 157960 34720 158120 34880
rect 157960 34880 158120 35040
rect 157960 35040 158120 35200
rect 157960 35200 158120 35360
rect 157960 35360 158120 35520
rect 157960 35520 158120 35680
rect 157960 35680 158120 35840
rect 157960 35840 158120 36000
rect 157960 36000 158120 36160
rect 157960 42080 158120 42240
rect 157960 42240 158120 42400
rect 157960 42400 158120 42560
rect 157960 42560 158120 42720
rect 157960 42720 158120 42880
rect 157960 42880 158120 43040
rect 157960 43040 158120 43200
rect 157960 43200 158120 43360
rect 157960 43360 158120 43520
rect 157960 43520 158120 43680
rect 157960 43680 158120 43840
rect 157960 43840 158120 44000
rect 157960 44000 158120 44160
rect 157960 44160 158120 44320
rect 157960 44320 158120 44480
rect 157960 44480 158120 44640
rect 157960 44640 158120 44800
rect 157960 44800 158120 44960
rect 157960 44960 158120 45120
rect 157960 45120 158120 45280
rect 157960 45280 158120 45440
rect 157960 45440 158120 45600
rect 157960 45600 158120 45760
rect 157960 45760 158120 45920
rect 157960 45920 158120 46080
rect 157960 46080 158120 46240
rect 157960 46240 158120 46400
rect 157960 46400 158120 46560
rect 157960 46560 158120 46720
rect 157960 46720 158120 46880
rect 157960 46880 158120 47040
rect 158120 31040 158280 31200
rect 158120 31200 158280 31360
rect 158120 31360 158280 31520
rect 158120 31520 158280 31680
rect 158120 31680 158280 31840
rect 158120 31840 158280 32000
rect 158120 32000 158280 32160
rect 158120 32160 158280 32320
rect 158120 32320 158280 32480
rect 158120 32480 158280 32640
rect 158120 32640 158280 32800
rect 158120 32800 158280 32960
rect 158120 32960 158280 33120
rect 158120 33120 158280 33280
rect 158120 33280 158280 33440
rect 158120 33440 158280 33600
rect 158120 33600 158280 33760
rect 158120 33760 158280 33920
rect 158120 33920 158280 34080
rect 158120 34080 158280 34240
rect 158120 34240 158280 34400
rect 158120 34400 158280 34560
rect 158120 34560 158280 34720
rect 158120 34720 158280 34880
rect 158120 34880 158280 35040
rect 158120 35040 158280 35200
rect 158120 35200 158280 35360
rect 158120 35360 158280 35520
rect 158120 35520 158280 35680
rect 158120 35680 158280 35840
rect 158120 35840 158280 36000
rect 158120 42240 158280 42400
rect 158120 42400 158280 42560
rect 158120 42560 158280 42720
rect 158120 42720 158280 42880
rect 158120 42880 158280 43040
rect 158120 43040 158280 43200
rect 158120 43200 158280 43360
rect 158120 43360 158280 43520
rect 158120 43520 158280 43680
rect 158120 43680 158280 43840
rect 158120 43840 158280 44000
rect 158120 44000 158280 44160
rect 158120 44160 158280 44320
rect 158120 44320 158280 44480
rect 158120 44480 158280 44640
rect 158120 44640 158280 44800
rect 158120 44800 158280 44960
rect 158120 44960 158280 45120
rect 158120 45120 158280 45280
rect 158120 45280 158280 45440
rect 158120 45440 158280 45600
rect 158120 45600 158280 45760
rect 158120 45760 158280 45920
rect 158120 45920 158280 46080
rect 158120 46080 158280 46240
rect 158120 46240 158280 46400
rect 158120 46400 158280 46560
rect 158120 46560 158280 46720
rect 158120 46720 158280 46880
rect 158120 46880 158280 47040
rect 158120 47040 158280 47200
rect 158280 30880 158440 31040
rect 158280 31040 158440 31200
rect 158280 31200 158440 31360
rect 158280 31360 158440 31520
rect 158280 31520 158440 31680
rect 158280 31680 158440 31840
rect 158280 31840 158440 32000
rect 158280 32000 158440 32160
rect 158280 32160 158440 32320
rect 158280 32320 158440 32480
rect 158280 32480 158440 32640
rect 158280 32640 158440 32800
rect 158280 32800 158440 32960
rect 158280 32960 158440 33120
rect 158280 33120 158440 33280
rect 158280 33280 158440 33440
rect 158280 33440 158440 33600
rect 158280 33600 158440 33760
rect 158280 33760 158440 33920
rect 158280 33920 158440 34080
rect 158280 34080 158440 34240
rect 158280 34240 158440 34400
rect 158280 34400 158440 34560
rect 158280 34560 158440 34720
rect 158280 34720 158440 34880
rect 158280 34880 158440 35040
rect 158280 35040 158440 35200
rect 158280 35200 158440 35360
rect 158280 35360 158440 35520
rect 158280 35520 158440 35680
rect 158280 35680 158440 35840
rect 158280 42400 158440 42560
rect 158280 42560 158440 42720
rect 158280 42720 158440 42880
rect 158280 42880 158440 43040
rect 158280 43040 158440 43200
rect 158280 43200 158440 43360
rect 158280 43360 158440 43520
rect 158280 43520 158440 43680
rect 158280 43680 158440 43840
rect 158280 43840 158440 44000
rect 158280 44000 158440 44160
rect 158280 44160 158440 44320
rect 158280 44320 158440 44480
rect 158280 44480 158440 44640
rect 158280 44640 158440 44800
rect 158280 44800 158440 44960
rect 158280 44960 158440 45120
rect 158280 45120 158440 45280
rect 158280 45280 158440 45440
rect 158280 45440 158440 45600
rect 158280 45600 158440 45760
rect 158280 45760 158440 45920
rect 158280 45920 158440 46080
rect 158280 46080 158440 46240
rect 158280 46240 158440 46400
rect 158280 46400 158440 46560
rect 158280 46560 158440 46720
rect 158280 46720 158440 46880
rect 158280 46880 158440 47040
rect 158280 47040 158440 47200
rect 158280 47200 158440 47360
rect 158280 47360 158440 47520
rect 158440 30880 158600 31040
rect 158440 31040 158600 31200
rect 158440 31200 158600 31360
rect 158440 31360 158600 31520
rect 158440 31520 158600 31680
rect 158440 31680 158600 31840
rect 158440 31840 158600 32000
rect 158440 32000 158600 32160
rect 158440 32160 158600 32320
rect 158440 32320 158600 32480
rect 158440 32480 158600 32640
rect 158440 32640 158600 32800
rect 158440 32800 158600 32960
rect 158440 32960 158600 33120
rect 158440 33120 158600 33280
rect 158440 33280 158600 33440
rect 158440 33440 158600 33600
rect 158440 33600 158600 33760
rect 158440 33760 158600 33920
rect 158440 33920 158600 34080
rect 158440 34080 158600 34240
rect 158440 34240 158600 34400
rect 158440 34400 158600 34560
rect 158440 34560 158600 34720
rect 158440 34720 158600 34880
rect 158440 34880 158600 35040
rect 158440 35040 158600 35200
rect 158440 35200 158600 35360
rect 158440 35360 158600 35520
rect 158440 35520 158600 35680
rect 158440 42560 158600 42720
rect 158440 42720 158600 42880
rect 158440 42880 158600 43040
rect 158440 43040 158600 43200
rect 158440 43200 158600 43360
rect 158440 43360 158600 43520
rect 158440 43520 158600 43680
rect 158440 43680 158600 43840
rect 158440 43840 158600 44000
rect 158440 44000 158600 44160
rect 158440 44160 158600 44320
rect 158440 44320 158600 44480
rect 158440 44480 158600 44640
rect 158440 44640 158600 44800
rect 158440 44800 158600 44960
rect 158440 44960 158600 45120
rect 158440 45120 158600 45280
rect 158440 45280 158600 45440
rect 158440 45440 158600 45600
rect 158440 45600 158600 45760
rect 158440 45760 158600 45920
rect 158440 45920 158600 46080
rect 158440 46080 158600 46240
rect 158440 46240 158600 46400
rect 158440 46400 158600 46560
rect 158440 46560 158600 46720
rect 158440 46720 158600 46880
rect 158440 46880 158600 47040
rect 158440 47040 158600 47200
rect 158440 47200 158600 47360
rect 158440 47360 158600 47520
rect 158440 47520 158600 47680
rect 158600 30720 158760 30880
rect 158600 30880 158760 31040
rect 158600 31040 158760 31200
rect 158600 31200 158760 31360
rect 158600 31360 158760 31520
rect 158600 31520 158760 31680
rect 158600 31680 158760 31840
rect 158600 31840 158760 32000
rect 158600 32000 158760 32160
rect 158600 32160 158760 32320
rect 158600 32320 158760 32480
rect 158600 32480 158760 32640
rect 158600 32640 158760 32800
rect 158600 32800 158760 32960
rect 158600 32960 158760 33120
rect 158600 33120 158760 33280
rect 158600 33280 158760 33440
rect 158600 33440 158760 33600
rect 158600 33600 158760 33760
rect 158600 33760 158760 33920
rect 158600 33920 158760 34080
rect 158600 34080 158760 34240
rect 158600 34240 158760 34400
rect 158600 34400 158760 34560
rect 158600 34560 158760 34720
rect 158600 34720 158760 34880
rect 158600 34880 158760 35040
rect 158600 35040 158760 35200
rect 158600 35200 158760 35360
rect 158600 35360 158760 35520
rect 158600 42720 158760 42880
rect 158600 42880 158760 43040
rect 158600 43040 158760 43200
rect 158600 43200 158760 43360
rect 158600 43360 158760 43520
rect 158600 43520 158760 43680
rect 158600 43680 158760 43840
rect 158600 43840 158760 44000
rect 158600 44000 158760 44160
rect 158600 44160 158760 44320
rect 158600 44320 158760 44480
rect 158600 44480 158760 44640
rect 158600 44640 158760 44800
rect 158600 44800 158760 44960
rect 158600 44960 158760 45120
rect 158600 45120 158760 45280
rect 158600 45280 158760 45440
rect 158600 45440 158760 45600
rect 158600 45600 158760 45760
rect 158600 45760 158760 45920
rect 158600 45920 158760 46080
rect 158600 46080 158760 46240
rect 158600 46240 158760 46400
rect 158600 46400 158760 46560
rect 158600 46560 158760 46720
rect 158600 46720 158760 46880
rect 158600 46880 158760 47040
rect 158600 47040 158760 47200
rect 158600 47200 158760 47360
rect 158600 47360 158760 47520
rect 158600 47520 158760 47680
rect 158600 47680 158760 47840
rect 158760 30560 158920 30720
rect 158760 30720 158920 30880
rect 158760 30880 158920 31040
rect 158760 31040 158920 31200
rect 158760 31200 158920 31360
rect 158760 31360 158920 31520
rect 158760 31520 158920 31680
rect 158760 31680 158920 31840
rect 158760 31840 158920 32000
rect 158760 32000 158920 32160
rect 158760 32160 158920 32320
rect 158760 32320 158920 32480
rect 158760 32480 158920 32640
rect 158760 32640 158920 32800
rect 158760 32800 158920 32960
rect 158760 32960 158920 33120
rect 158760 33120 158920 33280
rect 158760 33280 158920 33440
rect 158760 33440 158920 33600
rect 158760 33600 158920 33760
rect 158760 33760 158920 33920
rect 158760 33920 158920 34080
rect 158760 34080 158920 34240
rect 158760 34240 158920 34400
rect 158760 34400 158920 34560
rect 158760 34560 158920 34720
rect 158760 34720 158920 34880
rect 158760 34880 158920 35040
rect 158760 35040 158920 35200
rect 158760 35200 158920 35360
rect 158760 42880 158920 43040
rect 158760 43040 158920 43200
rect 158760 43200 158920 43360
rect 158760 43360 158920 43520
rect 158760 43520 158920 43680
rect 158760 43680 158920 43840
rect 158760 43840 158920 44000
rect 158760 44000 158920 44160
rect 158760 44160 158920 44320
rect 158760 44320 158920 44480
rect 158760 44480 158920 44640
rect 158760 44640 158920 44800
rect 158760 44800 158920 44960
rect 158760 44960 158920 45120
rect 158760 45120 158920 45280
rect 158760 45280 158920 45440
rect 158760 45440 158920 45600
rect 158760 45600 158920 45760
rect 158760 45760 158920 45920
rect 158760 45920 158920 46080
rect 158760 46080 158920 46240
rect 158760 46240 158920 46400
rect 158760 46400 158920 46560
rect 158760 46560 158920 46720
rect 158760 46720 158920 46880
rect 158760 46880 158920 47040
rect 158760 47040 158920 47200
rect 158760 47200 158920 47360
rect 158760 47360 158920 47520
rect 158760 47520 158920 47680
rect 158760 47680 158920 47840
rect 158760 47840 158920 48000
rect 158920 30400 159080 30560
rect 158920 30560 159080 30720
rect 158920 30720 159080 30880
rect 158920 30880 159080 31040
rect 158920 31040 159080 31200
rect 158920 31200 159080 31360
rect 158920 31360 159080 31520
rect 158920 31520 159080 31680
rect 158920 31680 159080 31840
rect 158920 31840 159080 32000
rect 158920 32000 159080 32160
rect 158920 32160 159080 32320
rect 158920 32320 159080 32480
rect 158920 32480 159080 32640
rect 158920 32640 159080 32800
rect 158920 32800 159080 32960
rect 158920 32960 159080 33120
rect 158920 33120 159080 33280
rect 158920 33280 159080 33440
rect 158920 33440 159080 33600
rect 158920 33600 159080 33760
rect 158920 33760 159080 33920
rect 158920 33920 159080 34080
rect 158920 34080 159080 34240
rect 158920 34240 159080 34400
rect 158920 34400 159080 34560
rect 158920 34560 159080 34720
rect 158920 34720 159080 34880
rect 158920 34880 159080 35040
rect 158920 35040 159080 35200
rect 158920 43040 159080 43200
rect 158920 43200 159080 43360
rect 158920 43360 159080 43520
rect 158920 43520 159080 43680
rect 158920 43680 159080 43840
rect 158920 43840 159080 44000
rect 158920 44000 159080 44160
rect 158920 44160 159080 44320
rect 158920 44320 159080 44480
rect 158920 44480 159080 44640
rect 158920 44640 159080 44800
rect 158920 44800 159080 44960
rect 158920 44960 159080 45120
rect 158920 45120 159080 45280
rect 158920 45280 159080 45440
rect 158920 45440 159080 45600
rect 158920 45600 159080 45760
rect 158920 45760 159080 45920
rect 158920 45920 159080 46080
rect 158920 46080 159080 46240
rect 158920 46240 159080 46400
rect 158920 46400 159080 46560
rect 158920 46560 159080 46720
rect 158920 46720 159080 46880
rect 158920 46880 159080 47040
rect 158920 47040 159080 47200
rect 158920 47200 159080 47360
rect 158920 47360 159080 47520
rect 158920 47520 159080 47680
rect 158920 47680 159080 47840
rect 158920 47840 159080 48000
rect 158920 48000 159080 48160
rect 159080 30240 159240 30400
rect 159080 30400 159240 30560
rect 159080 30560 159240 30720
rect 159080 30720 159240 30880
rect 159080 30880 159240 31040
rect 159080 31040 159240 31200
rect 159080 31200 159240 31360
rect 159080 31360 159240 31520
rect 159080 31520 159240 31680
rect 159080 31680 159240 31840
rect 159080 31840 159240 32000
rect 159080 32000 159240 32160
rect 159080 32160 159240 32320
rect 159080 32320 159240 32480
rect 159080 32480 159240 32640
rect 159080 32640 159240 32800
rect 159080 32800 159240 32960
rect 159080 32960 159240 33120
rect 159080 33120 159240 33280
rect 159080 33280 159240 33440
rect 159080 33440 159240 33600
rect 159080 33600 159240 33760
rect 159080 33760 159240 33920
rect 159080 33920 159240 34080
rect 159080 34080 159240 34240
rect 159080 34240 159240 34400
rect 159080 34400 159240 34560
rect 159080 34560 159240 34720
rect 159080 34720 159240 34880
rect 159080 34880 159240 35040
rect 159080 43200 159240 43360
rect 159080 43360 159240 43520
rect 159080 43520 159240 43680
rect 159080 43680 159240 43840
rect 159080 43840 159240 44000
rect 159080 44000 159240 44160
rect 159080 44160 159240 44320
rect 159080 44320 159240 44480
rect 159080 44480 159240 44640
rect 159080 44640 159240 44800
rect 159080 44800 159240 44960
rect 159080 44960 159240 45120
rect 159080 45120 159240 45280
rect 159080 45280 159240 45440
rect 159080 45440 159240 45600
rect 159080 45600 159240 45760
rect 159080 45760 159240 45920
rect 159080 45920 159240 46080
rect 159080 46080 159240 46240
rect 159080 46240 159240 46400
rect 159080 46400 159240 46560
rect 159080 46560 159240 46720
rect 159080 46720 159240 46880
rect 159080 46880 159240 47040
rect 159080 47040 159240 47200
rect 159080 47200 159240 47360
rect 159080 47360 159240 47520
rect 159080 47520 159240 47680
rect 159080 47680 159240 47840
rect 159080 47840 159240 48000
rect 159080 48000 159240 48160
rect 159080 48160 159240 48320
rect 159240 30080 159400 30240
rect 159240 30240 159400 30400
rect 159240 30400 159400 30560
rect 159240 30560 159400 30720
rect 159240 30720 159400 30880
rect 159240 30880 159400 31040
rect 159240 31040 159400 31200
rect 159240 31200 159400 31360
rect 159240 31360 159400 31520
rect 159240 31520 159400 31680
rect 159240 31680 159400 31840
rect 159240 31840 159400 32000
rect 159240 32000 159400 32160
rect 159240 32160 159400 32320
rect 159240 32320 159400 32480
rect 159240 32480 159400 32640
rect 159240 32640 159400 32800
rect 159240 32800 159400 32960
rect 159240 32960 159400 33120
rect 159240 33120 159400 33280
rect 159240 33280 159400 33440
rect 159240 33440 159400 33600
rect 159240 33600 159400 33760
rect 159240 33760 159400 33920
rect 159240 33920 159400 34080
rect 159240 34080 159400 34240
rect 159240 34240 159400 34400
rect 159240 34400 159400 34560
rect 159240 34560 159400 34720
rect 159240 34720 159400 34880
rect 159240 43360 159400 43520
rect 159240 43520 159400 43680
rect 159240 43680 159400 43840
rect 159240 43840 159400 44000
rect 159240 44000 159400 44160
rect 159240 44160 159400 44320
rect 159240 44320 159400 44480
rect 159240 44480 159400 44640
rect 159240 44640 159400 44800
rect 159240 44800 159400 44960
rect 159240 44960 159400 45120
rect 159240 45120 159400 45280
rect 159240 45280 159400 45440
rect 159240 45440 159400 45600
rect 159240 45600 159400 45760
rect 159240 45760 159400 45920
rect 159240 45920 159400 46080
rect 159240 46080 159400 46240
rect 159240 46240 159400 46400
rect 159240 46400 159400 46560
rect 159240 46560 159400 46720
rect 159240 46720 159400 46880
rect 159240 46880 159400 47040
rect 159240 47040 159400 47200
rect 159240 47200 159400 47360
rect 159240 47360 159400 47520
rect 159240 47520 159400 47680
rect 159240 47680 159400 47840
rect 159240 47840 159400 48000
rect 159240 48000 159400 48160
rect 159240 48160 159400 48320
rect 159240 48320 159400 48480
rect 159240 48480 159400 48640
rect 159400 29920 159560 30080
rect 159400 30080 159560 30240
rect 159400 30240 159560 30400
rect 159400 30400 159560 30560
rect 159400 30560 159560 30720
rect 159400 30720 159560 30880
rect 159400 30880 159560 31040
rect 159400 31040 159560 31200
rect 159400 31200 159560 31360
rect 159400 31360 159560 31520
rect 159400 31520 159560 31680
rect 159400 31680 159560 31840
rect 159400 31840 159560 32000
rect 159400 32000 159560 32160
rect 159400 32160 159560 32320
rect 159400 32320 159560 32480
rect 159400 32480 159560 32640
rect 159400 32640 159560 32800
rect 159400 32800 159560 32960
rect 159400 32960 159560 33120
rect 159400 33120 159560 33280
rect 159400 33280 159560 33440
rect 159400 33440 159560 33600
rect 159400 33600 159560 33760
rect 159400 33760 159560 33920
rect 159400 33920 159560 34080
rect 159400 34080 159560 34240
rect 159400 34240 159560 34400
rect 159400 34400 159560 34560
rect 159400 34560 159560 34720
rect 159400 43520 159560 43680
rect 159400 43680 159560 43840
rect 159400 43840 159560 44000
rect 159400 44000 159560 44160
rect 159400 44160 159560 44320
rect 159400 44320 159560 44480
rect 159400 44480 159560 44640
rect 159400 44640 159560 44800
rect 159400 44800 159560 44960
rect 159400 44960 159560 45120
rect 159400 45120 159560 45280
rect 159400 45280 159560 45440
rect 159400 45440 159560 45600
rect 159400 45600 159560 45760
rect 159400 45760 159560 45920
rect 159400 45920 159560 46080
rect 159400 46080 159560 46240
rect 159400 46240 159560 46400
rect 159400 46400 159560 46560
rect 159400 46560 159560 46720
rect 159400 46720 159560 46880
rect 159400 46880 159560 47040
rect 159400 47040 159560 47200
rect 159400 47200 159560 47360
rect 159400 47360 159560 47520
rect 159400 47520 159560 47680
rect 159400 47680 159560 47840
rect 159400 47840 159560 48000
rect 159400 48000 159560 48160
rect 159400 48160 159560 48320
rect 159400 48320 159560 48480
rect 159400 48480 159560 48640
rect 159400 48640 159560 48800
rect 159560 29760 159720 29920
rect 159560 29920 159720 30080
rect 159560 30080 159720 30240
rect 159560 30240 159720 30400
rect 159560 30400 159720 30560
rect 159560 30560 159720 30720
rect 159560 30720 159720 30880
rect 159560 30880 159720 31040
rect 159560 31040 159720 31200
rect 159560 31200 159720 31360
rect 159560 31360 159720 31520
rect 159560 31520 159720 31680
rect 159560 31680 159720 31840
rect 159560 31840 159720 32000
rect 159560 32000 159720 32160
rect 159560 32160 159720 32320
rect 159560 32320 159720 32480
rect 159560 32480 159720 32640
rect 159560 32640 159720 32800
rect 159560 32800 159720 32960
rect 159560 32960 159720 33120
rect 159560 33120 159720 33280
rect 159560 33280 159720 33440
rect 159560 33440 159720 33600
rect 159560 33600 159720 33760
rect 159560 33760 159720 33920
rect 159560 33920 159720 34080
rect 159560 34080 159720 34240
rect 159560 34240 159720 34400
rect 159560 34400 159720 34560
rect 159560 34560 159720 34720
rect 159560 43680 159720 43840
rect 159560 43840 159720 44000
rect 159560 44000 159720 44160
rect 159560 44160 159720 44320
rect 159560 44320 159720 44480
rect 159560 44480 159720 44640
rect 159560 44640 159720 44800
rect 159560 44800 159720 44960
rect 159560 44960 159720 45120
rect 159560 45120 159720 45280
rect 159560 45280 159720 45440
rect 159560 45440 159720 45600
rect 159560 45600 159720 45760
rect 159560 45760 159720 45920
rect 159560 45920 159720 46080
rect 159560 46080 159720 46240
rect 159560 46240 159720 46400
rect 159560 46400 159720 46560
rect 159560 46560 159720 46720
rect 159560 46720 159720 46880
rect 159560 46880 159720 47040
rect 159560 47040 159720 47200
rect 159560 47200 159720 47360
rect 159560 47360 159720 47520
rect 159560 47520 159720 47680
rect 159560 47680 159720 47840
rect 159560 47840 159720 48000
rect 159560 48000 159720 48160
rect 159560 48160 159720 48320
rect 159560 48320 159720 48480
rect 159560 48480 159720 48640
rect 159560 48640 159720 48800
rect 159560 48800 159720 48960
rect 159720 29760 159880 29920
rect 159720 29920 159880 30080
rect 159720 30080 159880 30240
rect 159720 30240 159880 30400
rect 159720 30400 159880 30560
rect 159720 30560 159880 30720
rect 159720 30720 159880 30880
rect 159720 30880 159880 31040
rect 159720 31040 159880 31200
rect 159720 31200 159880 31360
rect 159720 31360 159880 31520
rect 159720 31520 159880 31680
rect 159720 31680 159880 31840
rect 159720 31840 159880 32000
rect 159720 32000 159880 32160
rect 159720 32160 159880 32320
rect 159720 32320 159880 32480
rect 159720 32480 159880 32640
rect 159720 32640 159880 32800
rect 159720 32800 159880 32960
rect 159720 32960 159880 33120
rect 159720 33120 159880 33280
rect 159720 33280 159880 33440
rect 159720 33440 159880 33600
rect 159720 33600 159880 33760
rect 159720 33760 159880 33920
rect 159720 33920 159880 34080
rect 159720 34080 159880 34240
rect 159720 34240 159880 34400
rect 159720 34400 159880 34560
rect 159720 43840 159880 44000
rect 159720 44000 159880 44160
rect 159720 44160 159880 44320
rect 159720 44320 159880 44480
rect 159720 44480 159880 44640
rect 159720 44640 159880 44800
rect 159720 44800 159880 44960
rect 159720 44960 159880 45120
rect 159720 45120 159880 45280
rect 159720 45280 159880 45440
rect 159720 45440 159880 45600
rect 159720 45600 159880 45760
rect 159720 45760 159880 45920
rect 159720 45920 159880 46080
rect 159720 46080 159880 46240
rect 159720 46240 159880 46400
rect 159720 46400 159880 46560
rect 159720 46560 159880 46720
rect 159720 46720 159880 46880
rect 159720 46880 159880 47040
rect 159720 47040 159880 47200
rect 159720 47200 159880 47360
rect 159720 47360 159880 47520
rect 159720 47520 159880 47680
rect 159720 47680 159880 47840
rect 159720 47840 159880 48000
rect 159720 48000 159880 48160
rect 159720 48160 159880 48320
rect 159720 48320 159880 48480
rect 159720 48480 159880 48640
rect 159720 48640 159880 48800
rect 159720 48800 159880 48960
rect 159720 48960 159880 49120
rect 159880 29600 160040 29760
rect 159880 29760 160040 29920
rect 159880 29920 160040 30080
rect 159880 30080 160040 30240
rect 159880 30240 160040 30400
rect 159880 30400 160040 30560
rect 159880 30560 160040 30720
rect 159880 30720 160040 30880
rect 159880 30880 160040 31040
rect 159880 31040 160040 31200
rect 159880 31200 160040 31360
rect 159880 31360 160040 31520
rect 159880 31520 160040 31680
rect 159880 31680 160040 31840
rect 159880 31840 160040 32000
rect 159880 32000 160040 32160
rect 159880 32160 160040 32320
rect 159880 32320 160040 32480
rect 159880 32480 160040 32640
rect 159880 32640 160040 32800
rect 159880 32800 160040 32960
rect 159880 32960 160040 33120
rect 159880 33120 160040 33280
rect 159880 33280 160040 33440
rect 159880 33440 160040 33600
rect 159880 33600 160040 33760
rect 159880 33760 160040 33920
rect 159880 33920 160040 34080
rect 159880 34080 160040 34240
rect 159880 34240 160040 34400
rect 159880 44000 160040 44160
rect 159880 44160 160040 44320
rect 159880 44320 160040 44480
rect 159880 44480 160040 44640
rect 159880 44640 160040 44800
rect 159880 44800 160040 44960
rect 159880 44960 160040 45120
rect 159880 45120 160040 45280
rect 159880 45280 160040 45440
rect 159880 45440 160040 45600
rect 159880 45600 160040 45760
rect 159880 45760 160040 45920
rect 159880 45920 160040 46080
rect 159880 46080 160040 46240
rect 159880 46240 160040 46400
rect 159880 46400 160040 46560
rect 159880 46560 160040 46720
rect 159880 46720 160040 46880
rect 159880 46880 160040 47040
rect 159880 47040 160040 47200
rect 159880 47200 160040 47360
rect 159880 47360 160040 47520
rect 159880 47520 160040 47680
rect 159880 47680 160040 47840
rect 159880 47840 160040 48000
rect 159880 48000 160040 48160
rect 159880 48160 160040 48320
rect 159880 48320 160040 48480
rect 159880 48480 160040 48640
rect 159880 48640 160040 48800
rect 159880 48800 160040 48960
rect 159880 48960 160040 49120
rect 159880 49120 160040 49280
rect 160040 29440 160200 29600
rect 160040 29600 160200 29760
rect 160040 29760 160200 29920
rect 160040 29920 160200 30080
rect 160040 30080 160200 30240
rect 160040 30240 160200 30400
rect 160040 30400 160200 30560
rect 160040 30560 160200 30720
rect 160040 30720 160200 30880
rect 160040 30880 160200 31040
rect 160040 31040 160200 31200
rect 160040 31200 160200 31360
rect 160040 31360 160200 31520
rect 160040 31520 160200 31680
rect 160040 31680 160200 31840
rect 160040 31840 160200 32000
rect 160040 32000 160200 32160
rect 160040 32160 160200 32320
rect 160040 32320 160200 32480
rect 160040 32480 160200 32640
rect 160040 32640 160200 32800
rect 160040 32800 160200 32960
rect 160040 32960 160200 33120
rect 160040 33120 160200 33280
rect 160040 33280 160200 33440
rect 160040 33440 160200 33600
rect 160040 33600 160200 33760
rect 160040 33760 160200 33920
rect 160040 33920 160200 34080
rect 160040 34080 160200 34240
rect 160040 44160 160200 44320
rect 160040 44320 160200 44480
rect 160040 44480 160200 44640
rect 160040 44640 160200 44800
rect 160040 44800 160200 44960
rect 160040 44960 160200 45120
rect 160040 45120 160200 45280
rect 160040 45280 160200 45440
rect 160040 45440 160200 45600
rect 160040 45600 160200 45760
rect 160040 45760 160200 45920
rect 160040 45920 160200 46080
rect 160040 46080 160200 46240
rect 160040 46240 160200 46400
rect 160040 46400 160200 46560
rect 160040 46560 160200 46720
rect 160040 46720 160200 46880
rect 160040 46880 160200 47040
rect 160040 47040 160200 47200
rect 160040 47200 160200 47360
rect 160040 47360 160200 47520
rect 160040 47520 160200 47680
rect 160040 47680 160200 47840
rect 160040 47840 160200 48000
rect 160040 48000 160200 48160
rect 160040 48160 160200 48320
rect 160040 48320 160200 48480
rect 160040 48480 160200 48640
rect 160040 48640 160200 48800
rect 160040 48800 160200 48960
rect 160040 48960 160200 49120
rect 160040 49120 160200 49280
rect 160040 49280 160200 49440
rect 160200 29280 160360 29440
rect 160200 29440 160360 29600
rect 160200 29600 160360 29760
rect 160200 29760 160360 29920
rect 160200 29920 160360 30080
rect 160200 30080 160360 30240
rect 160200 30240 160360 30400
rect 160200 30400 160360 30560
rect 160200 30560 160360 30720
rect 160200 30720 160360 30880
rect 160200 30880 160360 31040
rect 160200 31040 160360 31200
rect 160200 31200 160360 31360
rect 160200 31360 160360 31520
rect 160200 31520 160360 31680
rect 160200 31680 160360 31840
rect 160200 31840 160360 32000
rect 160200 32000 160360 32160
rect 160200 32160 160360 32320
rect 160200 32320 160360 32480
rect 160200 32480 160360 32640
rect 160200 32640 160360 32800
rect 160200 32800 160360 32960
rect 160200 32960 160360 33120
rect 160200 33120 160360 33280
rect 160200 33280 160360 33440
rect 160200 33440 160360 33600
rect 160200 33600 160360 33760
rect 160200 33760 160360 33920
rect 160200 33920 160360 34080
rect 160200 44320 160360 44480
rect 160200 44480 160360 44640
rect 160200 44640 160360 44800
rect 160200 44800 160360 44960
rect 160200 44960 160360 45120
rect 160200 45120 160360 45280
rect 160200 45280 160360 45440
rect 160200 45440 160360 45600
rect 160200 45600 160360 45760
rect 160200 45760 160360 45920
rect 160200 45920 160360 46080
rect 160200 46080 160360 46240
rect 160200 46240 160360 46400
rect 160200 46400 160360 46560
rect 160200 46560 160360 46720
rect 160200 46720 160360 46880
rect 160200 46880 160360 47040
rect 160200 47040 160360 47200
rect 160200 47200 160360 47360
rect 160200 47360 160360 47520
rect 160200 47520 160360 47680
rect 160200 47680 160360 47840
rect 160200 47840 160360 48000
rect 160200 48000 160360 48160
rect 160200 48160 160360 48320
rect 160200 48320 160360 48480
rect 160200 48480 160360 48640
rect 160200 48640 160360 48800
rect 160200 48800 160360 48960
rect 160200 48960 160360 49120
rect 160200 49120 160360 49280
rect 160200 49280 160360 49440
rect 160200 49440 160360 49600
rect 160360 29120 160520 29280
rect 160360 29280 160520 29440
rect 160360 29440 160520 29600
rect 160360 29600 160520 29760
rect 160360 29760 160520 29920
rect 160360 29920 160520 30080
rect 160360 30080 160520 30240
rect 160360 30240 160520 30400
rect 160360 30400 160520 30560
rect 160360 30560 160520 30720
rect 160360 30720 160520 30880
rect 160360 30880 160520 31040
rect 160360 31040 160520 31200
rect 160360 31200 160520 31360
rect 160360 31360 160520 31520
rect 160360 31520 160520 31680
rect 160360 31680 160520 31840
rect 160360 31840 160520 32000
rect 160360 32000 160520 32160
rect 160360 32160 160520 32320
rect 160360 32320 160520 32480
rect 160360 32480 160520 32640
rect 160360 32640 160520 32800
rect 160360 32800 160520 32960
rect 160360 32960 160520 33120
rect 160360 33120 160520 33280
rect 160360 33280 160520 33440
rect 160360 33440 160520 33600
rect 160360 33600 160520 33760
rect 160360 33760 160520 33920
rect 160360 44480 160520 44640
rect 160360 44640 160520 44800
rect 160360 44800 160520 44960
rect 160360 44960 160520 45120
rect 160360 45120 160520 45280
rect 160360 45280 160520 45440
rect 160360 45440 160520 45600
rect 160360 45600 160520 45760
rect 160360 45760 160520 45920
rect 160360 45920 160520 46080
rect 160360 46080 160520 46240
rect 160360 46240 160520 46400
rect 160360 46400 160520 46560
rect 160360 46560 160520 46720
rect 160360 46720 160520 46880
rect 160360 46880 160520 47040
rect 160360 47040 160520 47200
rect 160360 47200 160520 47360
rect 160360 47360 160520 47520
rect 160360 47520 160520 47680
rect 160360 47680 160520 47840
rect 160360 47840 160520 48000
rect 160360 48000 160520 48160
rect 160360 48160 160520 48320
rect 160360 48320 160520 48480
rect 160360 48480 160520 48640
rect 160360 48640 160520 48800
rect 160360 48800 160520 48960
rect 160360 48960 160520 49120
rect 160360 49120 160520 49280
rect 160360 49280 160520 49440
rect 160360 49440 160520 49600
rect 160360 49600 160520 49760
rect 160360 49760 160520 49920
rect 160520 29120 160680 29280
rect 160520 29280 160680 29440
rect 160520 29440 160680 29600
rect 160520 29600 160680 29760
rect 160520 29760 160680 29920
rect 160520 29920 160680 30080
rect 160520 30080 160680 30240
rect 160520 30240 160680 30400
rect 160520 30400 160680 30560
rect 160520 30560 160680 30720
rect 160520 30720 160680 30880
rect 160520 30880 160680 31040
rect 160520 31040 160680 31200
rect 160520 31200 160680 31360
rect 160520 31360 160680 31520
rect 160520 31520 160680 31680
rect 160520 31680 160680 31840
rect 160520 31840 160680 32000
rect 160520 32000 160680 32160
rect 160520 32160 160680 32320
rect 160520 32320 160680 32480
rect 160520 32480 160680 32640
rect 160520 32640 160680 32800
rect 160520 32800 160680 32960
rect 160520 32960 160680 33120
rect 160520 33120 160680 33280
rect 160520 33280 160680 33440
rect 160520 33440 160680 33600
rect 160520 33600 160680 33760
rect 160520 44640 160680 44800
rect 160520 44800 160680 44960
rect 160520 44960 160680 45120
rect 160520 45120 160680 45280
rect 160520 45280 160680 45440
rect 160520 45440 160680 45600
rect 160520 45600 160680 45760
rect 160520 45760 160680 45920
rect 160520 45920 160680 46080
rect 160520 46080 160680 46240
rect 160520 46240 160680 46400
rect 160520 46400 160680 46560
rect 160520 46560 160680 46720
rect 160520 46720 160680 46880
rect 160520 46880 160680 47040
rect 160520 47040 160680 47200
rect 160520 47200 160680 47360
rect 160520 47360 160680 47520
rect 160520 47520 160680 47680
rect 160520 47680 160680 47840
rect 160520 47840 160680 48000
rect 160520 48000 160680 48160
rect 160520 48160 160680 48320
rect 160520 48320 160680 48480
rect 160520 48480 160680 48640
rect 160520 48640 160680 48800
rect 160520 48800 160680 48960
rect 160520 48960 160680 49120
rect 160520 49120 160680 49280
rect 160520 49280 160680 49440
rect 160520 49440 160680 49600
rect 160520 49600 160680 49760
rect 160520 49760 160680 49920
rect 160520 49920 160680 50080
rect 160680 28960 160840 29120
rect 160680 29120 160840 29280
rect 160680 29280 160840 29440
rect 160680 29440 160840 29600
rect 160680 29600 160840 29760
rect 160680 29760 160840 29920
rect 160680 29920 160840 30080
rect 160680 30080 160840 30240
rect 160680 30240 160840 30400
rect 160680 30400 160840 30560
rect 160680 30560 160840 30720
rect 160680 30720 160840 30880
rect 160680 30880 160840 31040
rect 160680 31040 160840 31200
rect 160680 31200 160840 31360
rect 160680 31360 160840 31520
rect 160680 31520 160840 31680
rect 160680 31680 160840 31840
rect 160680 31840 160840 32000
rect 160680 32000 160840 32160
rect 160680 32160 160840 32320
rect 160680 32320 160840 32480
rect 160680 32480 160840 32640
rect 160680 32640 160840 32800
rect 160680 32800 160840 32960
rect 160680 32960 160840 33120
rect 160680 33120 160840 33280
rect 160680 33280 160840 33440
rect 160680 33440 160840 33600
rect 160680 44800 160840 44960
rect 160680 44960 160840 45120
rect 160680 45120 160840 45280
rect 160680 45280 160840 45440
rect 160680 45440 160840 45600
rect 160680 45600 160840 45760
rect 160680 45760 160840 45920
rect 160680 45920 160840 46080
rect 160680 46080 160840 46240
rect 160680 46240 160840 46400
rect 160680 46400 160840 46560
rect 160680 46560 160840 46720
rect 160680 46720 160840 46880
rect 160680 46880 160840 47040
rect 160680 47040 160840 47200
rect 160680 47200 160840 47360
rect 160680 47360 160840 47520
rect 160680 47520 160840 47680
rect 160680 47680 160840 47840
rect 160680 47840 160840 48000
rect 160680 48000 160840 48160
rect 160680 48160 160840 48320
rect 160680 48320 160840 48480
rect 160680 48480 160840 48640
rect 160680 48640 160840 48800
rect 160680 48800 160840 48960
rect 160680 48960 160840 49120
rect 160680 49120 160840 49280
rect 160680 49280 160840 49440
rect 160680 49440 160840 49600
rect 160680 49600 160840 49760
rect 160680 49760 160840 49920
rect 160680 49920 160840 50080
rect 160680 50080 160840 50240
rect 160840 28800 161000 28960
rect 160840 28960 161000 29120
rect 160840 29120 161000 29280
rect 160840 29280 161000 29440
rect 160840 29440 161000 29600
rect 160840 29600 161000 29760
rect 160840 29760 161000 29920
rect 160840 29920 161000 30080
rect 160840 30080 161000 30240
rect 160840 30240 161000 30400
rect 160840 30400 161000 30560
rect 160840 30560 161000 30720
rect 160840 30720 161000 30880
rect 160840 30880 161000 31040
rect 160840 31040 161000 31200
rect 160840 31200 161000 31360
rect 160840 31360 161000 31520
rect 160840 31520 161000 31680
rect 160840 31680 161000 31840
rect 160840 31840 161000 32000
rect 160840 32000 161000 32160
rect 160840 32160 161000 32320
rect 160840 32320 161000 32480
rect 160840 32480 161000 32640
rect 160840 32640 161000 32800
rect 160840 32800 161000 32960
rect 160840 32960 161000 33120
rect 160840 33120 161000 33280
rect 160840 33280 161000 33440
rect 160840 44960 161000 45120
rect 160840 45120 161000 45280
rect 160840 45280 161000 45440
rect 160840 45440 161000 45600
rect 160840 45600 161000 45760
rect 160840 45760 161000 45920
rect 160840 45920 161000 46080
rect 160840 46080 161000 46240
rect 160840 46240 161000 46400
rect 160840 46400 161000 46560
rect 160840 46560 161000 46720
rect 160840 46720 161000 46880
rect 160840 46880 161000 47040
rect 160840 47040 161000 47200
rect 160840 47200 161000 47360
rect 160840 47360 161000 47520
rect 160840 47520 161000 47680
rect 160840 47680 161000 47840
rect 160840 47840 161000 48000
rect 160840 48000 161000 48160
rect 160840 48160 161000 48320
rect 160840 48320 161000 48480
rect 160840 48480 161000 48640
rect 160840 48640 161000 48800
rect 160840 48800 161000 48960
rect 160840 48960 161000 49120
rect 160840 49120 161000 49280
rect 160840 49280 161000 49440
rect 160840 49440 161000 49600
rect 160840 49600 161000 49760
rect 160840 49760 161000 49920
rect 160840 49920 161000 50080
rect 160840 50080 161000 50240
rect 160840 50240 161000 50400
rect 161000 28640 161160 28800
rect 161000 28800 161160 28960
rect 161000 28960 161160 29120
rect 161000 29120 161160 29280
rect 161000 29280 161160 29440
rect 161000 29440 161160 29600
rect 161000 29600 161160 29760
rect 161000 29760 161160 29920
rect 161000 29920 161160 30080
rect 161000 30080 161160 30240
rect 161000 30240 161160 30400
rect 161000 30400 161160 30560
rect 161000 30560 161160 30720
rect 161000 30720 161160 30880
rect 161000 30880 161160 31040
rect 161000 31040 161160 31200
rect 161000 31200 161160 31360
rect 161000 31360 161160 31520
rect 161000 31520 161160 31680
rect 161000 31680 161160 31840
rect 161000 31840 161160 32000
rect 161000 32000 161160 32160
rect 161000 32160 161160 32320
rect 161000 32320 161160 32480
rect 161000 32480 161160 32640
rect 161000 32640 161160 32800
rect 161000 32800 161160 32960
rect 161000 32960 161160 33120
rect 161000 33120 161160 33280
rect 161000 45120 161160 45280
rect 161000 45280 161160 45440
rect 161000 45440 161160 45600
rect 161000 45600 161160 45760
rect 161000 45760 161160 45920
rect 161000 45920 161160 46080
rect 161000 46080 161160 46240
rect 161000 46240 161160 46400
rect 161000 46400 161160 46560
rect 161000 46560 161160 46720
rect 161000 46720 161160 46880
rect 161000 46880 161160 47040
rect 161000 47040 161160 47200
rect 161000 47200 161160 47360
rect 161000 47360 161160 47520
rect 161000 47520 161160 47680
rect 161000 47680 161160 47840
rect 161000 47840 161160 48000
rect 161000 48000 161160 48160
rect 161000 48160 161160 48320
rect 161000 48320 161160 48480
rect 161000 48480 161160 48640
rect 161000 48640 161160 48800
rect 161000 48800 161160 48960
rect 161000 48960 161160 49120
rect 161000 49120 161160 49280
rect 161000 49280 161160 49440
rect 161000 49440 161160 49600
rect 161000 49600 161160 49760
rect 161000 49760 161160 49920
rect 161000 49920 161160 50080
rect 161000 50080 161160 50240
rect 161000 50240 161160 50400
rect 161000 50400 161160 50560
rect 161160 28640 161320 28800
rect 161160 28800 161320 28960
rect 161160 28960 161320 29120
rect 161160 29120 161320 29280
rect 161160 29280 161320 29440
rect 161160 29440 161320 29600
rect 161160 29600 161320 29760
rect 161160 29760 161320 29920
rect 161160 29920 161320 30080
rect 161160 30080 161320 30240
rect 161160 30240 161320 30400
rect 161160 30400 161320 30560
rect 161160 30560 161320 30720
rect 161160 30720 161320 30880
rect 161160 30880 161320 31040
rect 161160 31040 161320 31200
rect 161160 31200 161320 31360
rect 161160 31360 161320 31520
rect 161160 31520 161320 31680
rect 161160 31680 161320 31840
rect 161160 31840 161320 32000
rect 161160 32000 161320 32160
rect 161160 32160 161320 32320
rect 161160 32320 161320 32480
rect 161160 32480 161320 32640
rect 161160 32640 161320 32800
rect 161160 32800 161320 32960
rect 161160 32960 161320 33120
rect 161160 45280 161320 45440
rect 161160 45440 161320 45600
rect 161160 45600 161320 45760
rect 161160 45760 161320 45920
rect 161160 45920 161320 46080
rect 161160 46080 161320 46240
rect 161160 46240 161320 46400
rect 161160 46400 161320 46560
rect 161160 46560 161320 46720
rect 161160 46720 161320 46880
rect 161160 46880 161320 47040
rect 161160 47040 161320 47200
rect 161160 47200 161320 47360
rect 161160 47360 161320 47520
rect 161160 47520 161320 47680
rect 161160 47680 161320 47840
rect 161160 47840 161320 48000
rect 161160 48000 161320 48160
rect 161160 48160 161320 48320
rect 161160 48320 161320 48480
rect 161160 48480 161320 48640
rect 161160 48640 161320 48800
rect 161160 48800 161320 48960
rect 161160 48960 161320 49120
rect 161160 49120 161320 49280
rect 161160 49280 161320 49440
rect 161160 49440 161320 49600
rect 161160 49600 161320 49760
rect 161160 49760 161320 49920
rect 161160 49920 161320 50080
rect 161160 50080 161320 50240
rect 161160 50240 161320 50400
rect 161160 50400 161320 50560
rect 161160 50560 161320 50720
rect 161320 28480 161480 28640
rect 161320 28640 161480 28800
rect 161320 28800 161480 28960
rect 161320 28960 161480 29120
rect 161320 29120 161480 29280
rect 161320 29280 161480 29440
rect 161320 29440 161480 29600
rect 161320 29600 161480 29760
rect 161320 29760 161480 29920
rect 161320 29920 161480 30080
rect 161320 30080 161480 30240
rect 161320 30240 161480 30400
rect 161320 30400 161480 30560
rect 161320 30560 161480 30720
rect 161320 30720 161480 30880
rect 161320 30880 161480 31040
rect 161320 31040 161480 31200
rect 161320 31200 161480 31360
rect 161320 31360 161480 31520
rect 161320 31520 161480 31680
rect 161320 31680 161480 31840
rect 161320 31840 161480 32000
rect 161320 32000 161480 32160
rect 161320 32160 161480 32320
rect 161320 32320 161480 32480
rect 161320 32480 161480 32640
rect 161320 32640 161480 32800
rect 161320 32800 161480 32960
rect 161320 45600 161480 45760
rect 161320 45760 161480 45920
rect 161320 45920 161480 46080
rect 161320 46080 161480 46240
rect 161320 46240 161480 46400
rect 161320 46400 161480 46560
rect 161320 46560 161480 46720
rect 161320 46720 161480 46880
rect 161320 46880 161480 47040
rect 161320 47040 161480 47200
rect 161320 47200 161480 47360
rect 161320 47360 161480 47520
rect 161320 47520 161480 47680
rect 161320 47680 161480 47840
rect 161320 47840 161480 48000
rect 161320 48000 161480 48160
rect 161320 48160 161480 48320
rect 161320 48320 161480 48480
rect 161320 48480 161480 48640
rect 161320 48640 161480 48800
rect 161320 48800 161480 48960
rect 161320 48960 161480 49120
rect 161320 49120 161480 49280
rect 161320 49280 161480 49440
rect 161320 49440 161480 49600
rect 161320 49600 161480 49760
rect 161320 49760 161480 49920
rect 161320 49920 161480 50080
rect 161320 50080 161480 50240
rect 161320 50240 161480 50400
rect 161320 50400 161480 50560
rect 161320 50560 161480 50720
rect 161320 50720 161480 50880
rect 161320 50880 161480 51040
rect 161480 28320 161640 28480
rect 161480 28480 161640 28640
rect 161480 28640 161640 28800
rect 161480 28800 161640 28960
rect 161480 28960 161640 29120
rect 161480 29120 161640 29280
rect 161480 29280 161640 29440
rect 161480 29440 161640 29600
rect 161480 29600 161640 29760
rect 161480 29760 161640 29920
rect 161480 29920 161640 30080
rect 161480 30080 161640 30240
rect 161480 30240 161640 30400
rect 161480 30400 161640 30560
rect 161480 30560 161640 30720
rect 161480 30720 161640 30880
rect 161480 30880 161640 31040
rect 161480 31040 161640 31200
rect 161480 31200 161640 31360
rect 161480 31360 161640 31520
rect 161480 31520 161640 31680
rect 161480 31680 161640 31840
rect 161480 31840 161640 32000
rect 161480 32000 161640 32160
rect 161480 32160 161640 32320
rect 161480 32320 161640 32480
rect 161480 32480 161640 32640
rect 161480 32640 161640 32800
rect 161480 45760 161640 45920
rect 161480 45920 161640 46080
rect 161480 46080 161640 46240
rect 161480 46240 161640 46400
rect 161480 46400 161640 46560
rect 161480 46560 161640 46720
rect 161480 46720 161640 46880
rect 161480 46880 161640 47040
rect 161480 47040 161640 47200
rect 161480 47200 161640 47360
rect 161480 47360 161640 47520
rect 161480 47520 161640 47680
rect 161480 47680 161640 47840
rect 161480 47840 161640 48000
rect 161480 48000 161640 48160
rect 161480 48160 161640 48320
rect 161480 48320 161640 48480
rect 161480 48480 161640 48640
rect 161480 48640 161640 48800
rect 161480 48800 161640 48960
rect 161480 48960 161640 49120
rect 161480 49120 161640 49280
rect 161480 49280 161640 49440
rect 161480 49440 161640 49600
rect 161480 49600 161640 49760
rect 161480 49760 161640 49920
rect 161480 49920 161640 50080
rect 161480 50080 161640 50240
rect 161480 50240 161640 50400
rect 161480 50400 161640 50560
rect 161480 50560 161640 50720
rect 161480 50720 161640 50880
rect 161480 50880 161640 51040
rect 161480 51040 161640 51200
rect 161640 28320 161800 28480
rect 161640 28480 161800 28640
rect 161640 28640 161800 28800
rect 161640 28800 161800 28960
rect 161640 28960 161800 29120
rect 161640 29120 161800 29280
rect 161640 29280 161800 29440
rect 161640 29440 161800 29600
rect 161640 29600 161800 29760
rect 161640 29760 161800 29920
rect 161640 29920 161800 30080
rect 161640 30080 161800 30240
rect 161640 30240 161800 30400
rect 161640 30400 161800 30560
rect 161640 30560 161800 30720
rect 161640 30720 161800 30880
rect 161640 30880 161800 31040
rect 161640 31040 161800 31200
rect 161640 31200 161800 31360
rect 161640 31360 161800 31520
rect 161640 31520 161800 31680
rect 161640 31680 161800 31840
rect 161640 31840 161800 32000
rect 161640 32000 161800 32160
rect 161640 32160 161800 32320
rect 161640 32320 161800 32480
rect 161640 32480 161800 32640
rect 161640 32640 161800 32800
rect 161640 45920 161800 46080
rect 161640 46080 161800 46240
rect 161640 46240 161800 46400
rect 161640 46400 161800 46560
rect 161640 46560 161800 46720
rect 161640 46720 161800 46880
rect 161640 46880 161800 47040
rect 161640 47040 161800 47200
rect 161640 47200 161800 47360
rect 161640 47360 161800 47520
rect 161640 47520 161800 47680
rect 161640 47680 161800 47840
rect 161640 47840 161800 48000
rect 161640 48000 161800 48160
rect 161640 48160 161800 48320
rect 161640 48320 161800 48480
rect 161640 48480 161800 48640
rect 161640 48640 161800 48800
rect 161640 48800 161800 48960
rect 161640 48960 161800 49120
rect 161640 49120 161800 49280
rect 161640 49280 161800 49440
rect 161640 49440 161800 49600
rect 161640 49600 161800 49760
rect 161640 49760 161800 49920
rect 161640 49920 161800 50080
rect 161640 50080 161800 50240
rect 161640 50240 161800 50400
rect 161640 50400 161800 50560
rect 161640 50560 161800 50720
rect 161640 50720 161800 50880
rect 161640 50880 161800 51040
rect 161640 51040 161800 51200
rect 161640 51200 161800 51360
rect 161800 28160 161960 28320
rect 161800 28320 161960 28480
rect 161800 28480 161960 28640
rect 161800 28640 161960 28800
rect 161800 28800 161960 28960
rect 161800 28960 161960 29120
rect 161800 29120 161960 29280
rect 161800 29280 161960 29440
rect 161800 29440 161960 29600
rect 161800 29600 161960 29760
rect 161800 29760 161960 29920
rect 161800 29920 161960 30080
rect 161800 30080 161960 30240
rect 161800 30240 161960 30400
rect 161800 30400 161960 30560
rect 161800 30560 161960 30720
rect 161800 30720 161960 30880
rect 161800 30880 161960 31040
rect 161800 31040 161960 31200
rect 161800 31200 161960 31360
rect 161800 31360 161960 31520
rect 161800 31520 161960 31680
rect 161800 31680 161960 31840
rect 161800 31840 161960 32000
rect 161800 32000 161960 32160
rect 161800 32160 161960 32320
rect 161800 32320 161960 32480
rect 161800 32480 161960 32640
rect 161800 46080 161960 46240
rect 161800 46240 161960 46400
rect 161800 46400 161960 46560
rect 161800 46560 161960 46720
rect 161800 46720 161960 46880
rect 161800 46880 161960 47040
rect 161800 47040 161960 47200
rect 161800 47200 161960 47360
rect 161800 47360 161960 47520
rect 161800 47520 161960 47680
rect 161800 47680 161960 47840
rect 161800 47840 161960 48000
rect 161800 48000 161960 48160
rect 161800 48160 161960 48320
rect 161800 48320 161960 48480
rect 161800 48480 161960 48640
rect 161800 48640 161960 48800
rect 161800 48800 161960 48960
rect 161800 48960 161960 49120
rect 161800 49120 161960 49280
rect 161800 49280 161960 49440
rect 161800 49440 161960 49600
rect 161800 49600 161960 49760
rect 161800 49760 161960 49920
rect 161800 49920 161960 50080
rect 161800 50080 161960 50240
rect 161800 50240 161960 50400
rect 161800 50400 161960 50560
rect 161800 50560 161960 50720
rect 161800 50720 161960 50880
rect 161800 50880 161960 51040
rect 161800 51040 161960 51200
rect 161800 51200 161960 51360
rect 161800 51360 161960 51520
rect 161960 28000 162120 28160
rect 161960 28160 162120 28320
rect 161960 28320 162120 28480
rect 161960 28480 162120 28640
rect 161960 28640 162120 28800
rect 161960 28800 162120 28960
rect 161960 28960 162120 29120
rect 161960 29120 162120 29280
rect 161960 29280 162120 29440
rect 161960 29440 162120 29600
rect 161960 29600 162120 29760
rect 161960 29760 162120 29920
rect 161960 29920 162120 30080
rect 161960 30080 162120 30240
rect 161960 30240 162120 30400
rect 161960 30400 162120 30560
rect 161960 30560 162120 30720
rect 161960 30720 162120 30880
rect 161960 30880 162120 31040
rect 161960 31040 162120 31200
rect 161960 31200 162120 31360
rect 161960 31360 162120 31520
rect 161960 31520 162120 31680
rect 161960 31680 162120 31840
rect 161960 31840 162120 32000
rect 161960 32000 162120 32160
rect 161960 32160 162120 32320
rect 161960 32320 162120 32480
rect 161960 46240 162120 46400
rect 161960 46400 162120 46560
rect 161960 46560 162120 46720
rect 161960 46720 162120 46880
rect 161960 46880 162120 47040
rect 161960 47040 162120 47200
rect 161960 47200 162120 47360
rect 161960 47360 162120 47520
rect 161960 47520 162120 47680
rect 161960 47680 162120 47840
rect 161960 47840 162120 48000
rect 161960 48000 162120 48160
rect 161960 48160 162120 48320
rect 161960 48320 162120 48480
rect 161960 48480 162120 48640
rect 161960 48640 162120 48800
rect 161960 48800 162120 48960
rect 161960 48960 162120 49120
rect 161960 49120 162120 49280
rect 161960 49280 162120 49440
rect 161960 49440 162120 49600
rect 161960 49600 162120 49760
rect 161960 49760 162120 49920
rect 161960 49920 162120 50080
rect 161960 50080 162120 50240
rect 161960 50240 162120 50400
rect 161960 50400 162120 50560
rect 161960 50560 162120 50720
rect 161960 50720 162120 50880
rect 161960 50880 162120 51040
rect 161960 51040 162120 51200
rect 161960 51200 162120 51360
rect 161960 51360 162120 51520
rect 161960 51520 162120 51680
rect 162120 28000 162280 28160
rect 162120 28160 162280 28320
rect 162120 28320 162280 28480
rect 162120 28480 162280 28640
rect 162120 28640 162280 28800
rect 162120 28800 162280 28960
rect 162120 28960 162280 29120
rect 162120 29120 162280 29280
rect 162120 29280 162280 29440
rect 162120 29440 162280 29600
rect 162120 29600 162280 29760
rect 162120 29760 162280 29920
rect 162120 29920 162280 30080
rect 162120 30080 162280 30240
rect 162120 30240 162280 30400
rect 162120 30400 162280 30560
rect 162120 30560 162280 30720
rect 162120 30720 162280 30880
rect 162120 30880 162280 31040
rect 162120 31040 162280 31200
rect 162120 31200 162280 31360
rect 162120 31360 162280 31520
rect 162120 31520 162280 31680
rect 162120 31680 162280 31840
rect 162120 31840 162280 32000
rect 162120 32000 162280 32160
rect 162120 32160 162280 32320
rect 162120 46400 162280 46560
rect 162120 46560 162280 46720
rect 162120 46720 162280 46880
rect 162120 46880 162280 47040
rect 162120 47040 162280 47200
rect 162120 47200 162280 47360
rect 162120 47360 162280 47520
rect 162120 47520 162280 47680
rect 162120 47680 162280 47840
rect 162120 47840 162280 48000
rect 162120 48000 162280 48160
rect 162120 48160 162280 48320
rect 162120 48320 162280 48480
rect 162120 48480 162280 48640
rect 162120 48640 162280 48800
rect 162120 48800 162280 48960
rect 162120 48960 162280 49120
rect 162120 49120 162280 49280
rect 162120 49280 162280 49440
rect 162120 49440 162280 49600
rect 162120 49600 162280 49760
rect 162120 49760 162280 49920
rect 162120 49920 162280 50080
rect 162120 50080 162280 50240
rect 162120 50240 162280 50400
rect 162120 50400 162280 50560
rect 162120 50560 162280 50720
rect 162120 50720 162280 50880
rect 162120 50880 162280 51040
rect 162120 51040 162280 51200
rect 162120 51200 162280 51360
rect 162120 51360 162280 51520
rect 162120 51520 162280 51680
rect 162120 51680 162280 51840
rect 162280 27840 162440 28000
rect 162280 28000 162440 28160
rect 162280 28160 162440 28320
rect 162280 28320 162440 28480
rect 162280 28480 162440 28640
rect 162280 28640 162440 28800
rect 162280 28800 162440 28960
rect 162280 28960 162440 29120
rect 162280 29120 162440 29280
rect 162280 29280 162440 29440
rect 162280 29440 162440 29600
rect 162280 29600 162440 29760
rect 162280 29760 162440 29920
rect 162280 29920 162440 30080
rect 162280 30080 162440 30240
rect 162280 30240 162440 30400
rect 162280 30400 162440 30560
rect 162280 30560 162440 30720
rect 162280 30720 162440 30880
rect 162280 30880 162440 31040
rect 162280 31040 162440 31200
rect 162280 31200 162440 31360
rect 162280 31360 162440 31520
rect 162280 31520 162440 31680
rect 162280 31680 162440 31840
rect 162280 31840 162440 32000
rect 162280 32000 162440 32160
rect 162280 46560 162440 46720
rect 162280 46720 162440 46880
rect 162280 46880 162440 47040
rect 162280 47040 162440 47200
rect 162280 47200 162440 47360
rect 162280 47360 162440 47520
rect 162280 47520 162440 47680
rect 162280 47680 162440 47840
rect 162280 47840 162440 48000
rect 162280 48000 162440 48160
rect 162280 48160 162440 48320
rect 162280 48320 162440 48480
rect 162280 48480 162440 48640
rect 162280 48640 162440 48800
rect 162280 48800 162440 48960
rect 162280 48960 162440 49120
rect 162280 49120 162440 49280
rect 162280 49280 162440 49440
rect 162280 49440 162440 49600
rect 162280 49600 162440 49760
rect 162280 49760 162440 49920
rect 162280 49920 162440 50080
rect 162280 50080 162440 50240
rect 162280 50240 162440 50400
rect 162280 50400 162440 50560
rect 162280 50560 162440 50720
rect 162280 50720 162440 50880
rect 162280 50880 162440 51040
rect 162280 51040 162440 51200
rect 162280 51200 162440 51360
rect 162280 51360 162440 51520
rect 162280 51520 162440 51680
rect 162280 51680 162440 51840
rect 162280 51840 162440 52000
rect 162280 52000 162440 52160
rect 162440 27840 162600 28000
rect 162440 28000 162600 28160
rect 162440 28160 162600 28320
rect 162440 28320 162600 28480
rect 162440 28480 162600 28640
rect 162440 28640 162600 28800
rect 162440 28800 162600 28960
rect 162440 28960 162600 29120
rect 162440 29120 162600 29280
rect 162440 29280 162600 29440
rect 162440 29440 162600 29600
rect 162440 29600 162600 29760
rect 162440 29760 162600 29920
rect 162440 29920 162600 30080
rect 162440 30080 162600 30240
rect 162440 30240 162600 30400
rect 162440 30400 162600 30560
rect 162440 30560 162600 30720
rect 162440 30720 162600 30880
rect 162440 30880 162600 31040
rect 162440 31040 162600 31200
rect 162440 31200 162600 31360
rect 162440 31360 162600 31520
rect 162440 31520 162600 31680
rect 162440 31680 162600 31840
rect 162440 31840 162600 32000
rect 162440 46880 162600 47040
rect 162440 47040 162600 47200
rect 162440 47200 162600 47360
rect 162440 47360 162600 47520
rect 162440 47520 162600 47680
rect 162440 47680 162600 47840
rect 162440 47840 162600 48000
rect 162440 48000 162600 48160
rect 162440 48160 162600 48320
rect 162440 48320 162600 48480
rect 162440 48480 162600 48640
rect 162440 48640 162600 48800
rect 162440 48800 162600 48960
rect 162440 48960 162600 49120
rect 162440 49120 162600 49280
rect 162440 49280 162600 49440
rect 162440 49440 162600 49600
rect 162440 49600 162600 49760
rect 162440 49760 162600 49920
rect 162440 49920 162600 50080
rect 162440 50080 162600 50240
rect 162440 50240 162600 50400
rect 162440 50400 162600 50560
rect 162440 50560 162600 50720
rect 162440 50720 162600 50880
rect 162440 50880 162600 51040
rect 162440 51040 162600 51200
rect 162440 51200 162600 51360
rect 162440 51360 162600 51520
rect 162440 51520 162600 51680
rect 162440 51680 162600 51840
rect 162440 51840 162600 52000
rect 162440 52000 162600 52160
rect 162440 52160 162600 52320
rect 162600 27680 162760 27840
rect 162600 27840 162760 28000
rect 162600 28000 162760 28160
rect 162600 28160 162760 28320
rect 162600 28320 162760 28480
rect 162600 28480 162760 28640
rect 162600 28640 162760 28800
rect 162600 28800 162760 28960
rect 162600 28960 162760 29120
rect 162600 29120 162760 29280
rect 162600 29280 162760 29440
rect 162600 29440 162760 29600
rect 162600 29600 162760 29760
rect 162600 29760 162760 29920
rect 162600 29920 162760 30080
rect 162600 30080 162760 30240
rect 162600 30240 162760 30400
rect 162600 30400 162760 30560
rect 162600 30560 162760 30720
rect 162600 30720 162760 30880
rect 162600 30880 162760 31040
rect 162600 31040 162760 31200
rect 162600 31200 162760 31360
rect 162600 31360 162760 31520
rect 162600 31520 162760 31680
rect 162600 31680 162760 31840
rect 162600 31840 162760 32000
rect 162600 47040 162760 47200
rect 162600 47200 162760 47360
rect 162600 47360 162760 47520
rect 162600 47520 162760 47680
rect 162600 47680 162760 47840
rect 162600 47840 162760 48000
rect 162600 48000 162760 48160
rect 162600 48160 162760 48320
rect 162600 48320 162760 48480
rect 162600 48480 162760 48640
rect 162600 48640 162760 48800
rect 162600 48800 162760 48960
rect 162600 48960 162760 49120
rect 162600 49120 162760 49280
rect 162600 49280 162760 49440
rect 162600 49440 162760 49600
rect 162600 49600 162760 49760
rect 162600 49760 162760 49920
rect 162600 49920 162760 50080
rect 162600 50080 162760 50240
rect 162600 50240 162760 50400
rect 162600 50400 162760 50560
rect 162600 50560 162760 50720
rect 162600 50720 162760 50880
rect 162600 50880 162760 51040
rect 162600 51040 162760 51200
rect 162600 51200 162760 51360
rect 162600 51360 162760 51520
rect 162600 51520 162760 51680
rect 162600 51680 162760 51840
rect 162600 51840 162760 52000
rect 162600 52000 162760 52160
rect 162600 52160 162760 52320
rect 162600 52320 162760 52480
rect 162760 27680 162920 27840
rect 162760 27840 162920 28000
rect 162760 28000 162920 28160
rect 162760 28160 162920 28320
rect 162760 28320 162920 28480
rect 162760 28480 162920 28640
rect 162760 28640 162920 28800
rect 162760 28800 162920 28960
rect 162760 28960 162920 29120
rect 162760 29120 162920 29280
rect 162760 29280 162920 29440
rect 162760 29440 162920 29600
rect 162760 29600 162920 29760
rect 162760 29760 162920 29920
rect 162760 29920 162920 30080
rect 162760 30080 162920 30240
rect 162760 30240 162920 30400
rect 162760 30400 162920 30560
rect 162760 30560 162920 30720
rect 162760 30720 162920 30880
rect 162760 30880 162920 31040
rect 162760 31040 162920 31200
rect 162760 31200 162920 31360
rect 162760 31360 162920 31520
rect 162760 31520 162920 31680
rect 162760 31680 162920 31840
rect 162760 47200 162920 47360
rect 162760 47360 162920 47520
rect 162760 47520 162920 47680
rect 162760 47680 162920 47840
rect 162760 47840 162920 48000
rect 162760 48000 162920 48160
rect 162760 48160 162920 48320
rect 162760 48320 162920 48480
rect 162760 48480 162920 48640
rect 162760 48640 162920 48800
rect 162760 48800 162920 48960
rect 162760 48960 162920 49120
rect 162760 49120 162920 49280
rect 162760 49280 162920 49440
rect 162760 49440 162920 49600
rect 162760 49600 162920 49760
rect 162760 49760 162920 49920
rect 162760 49920 162920 50080
rect 162760 50080 162920 50240
rect 162760 50240 162920 50400
rect 162760 50400 162920 50560
rect 162760 50560 162920 50720
rect 162760 50720 162920 50880
rect 162760 50880 162920 51040
rect 162760 51040 162920 51200
rect 162760 51200 162920 51360
rect 162760 51360 162920 51520
rect 162760 51520 162920 51680
rect 162760 51680 162920 51840
rect 162760 51840 162920 52000
rect 162760 52000 162920 52160
rect 162760 52160 162920 52320
rect 162760 52320 162920 52480
rect 162760 52480 162920 52640
rect 162920 27520 163080 27680
rect 162920 27680 163080 27840
rect 162920 27840 163080 28000
rect 162920 28000 163080 28160
rect 162920 28160 163080 28320
rect 162920 28320 163080 28480
rect 162920 28480 163080 28640
rect 162920 28640 163080 28800
rect 162920 28800 163080 28960
rect 162920 28960 163080 29120
rect 162920 29120 163080 29280
rect 162920 29280 163080 29440
rect 162920 29440 163080 29600
rect 162920 29600 163080 29760
rect 162920 29760 163080 29920
rect 162920 29920 163080 30080
rect 162920 30080 163080 30240
rect 162920 30240 163080 30400
rect 162920 30400 163080 30560
rect 162920 30560 163080 30720
rect 162920 30720 163080 30880
rect 162920 30880 163080 31040
rect 162920 31040 163080 31200
rect 162920 31200 163080 31360
rect 162920 31360 163080 31520
rect 162920 31520 163080 31680
rect 162920 47360 163080 47520
rect 162920 47520 163080 47680
rect 162920 47680 163080 47840
rect 162920 47840 163080 48000
rect 162920 48000 163080 48160
rect 162920 48160 163080 48320
rect 162920 48320 163080 48480
rect 162920 48480 163080 48640
rect 162920 48640 163080 48800
rect 162920 48800 163080 48960
rect 162920 48960 163080 49120
rect 162920 49120 163080 49280
rect 162920 49280 163080 49440
rect 162920 49440 163080 49600
rect 162920 49600 163080 49760
rect 162920 49760 163080 49920
rect 162920 49920 163080 50080
rect 162920 50080 163080 50240
rect 162920 50240 163080 50400
rect 162920 50400 163080 50560
rect 162920 50560 163080 50720
rect 162920 50720 163080 50880
rect 162920 50880 163080 51040
rect 162920 51040 163080 51200
rect 162920 51200 163080 51360
rect 162920 51360 163080 51520
rect 162920 51520 163080 51680
rect 162920 51680 163080 51840
rect 162920 51840 163080 52000
rect 162920 52000 163080 52160
rect 162920 52160 163080 52320
rect 162920 52320 163080 52480
rect 162920 52480 163080 52640
rect 162920 52640 163080 52800
rect 163080 27520 163240 27680
rect 163080 27680 163240 27840
rect 163080 27840 163240 28000
rect 163080 28000 163240 28160
rect 163080 28160 163240 28320
rect 163080 28320 163240 28480
rect 163080 28480 163240 28640
rect 163080 28640 163240 28800
rect 163080 28800 163240 28960
rect 163080 28960 163240 29120
rect 163080 29120 163240 29280
rect 163080 29280 163240 29440
rect 163080 29440 163240 29600
rect 163080 29600 163240 29760
rect 163080 29760 163240 29920
rect 163080 29920 163240 30080
rect 163080 30080 163240 30240
rect 163080 30240 163240 30400
rect 163080 30400 163240 30560
rect 163080 30560 163240 30720
rect 163080 30720 163240 30880
rect 163080 30880 163240 31040
rect 163080 31040 163240 31200
rect 163080 31200 163240 31360
rect 163080 31360 163240 31520
rect 163080 47520 163240 47680
rect 163080 47680 163240 47840
rect 163080 47840 163240 48000
rect 163080 48000 163240 48160
rect 163080 48160 163240 48320
rect 163080 48320 163240 48480
rect 163080 48480 163240 48640
rect 163080 48640 163240 48800
rect 163080 48800 163240 48960
rect 163080 48960 163240 49120
rect 163080 49120 163240 49280
rect 163080 49280 163240 49440
rect 163080 49440 163240 49600
rect 163080 49600 163240 49760
rect 163080 49760 163240 49920
rect 163080 49920 163240 50080
rect 163080 50080 163240 50240
rect 163080 50240 163240 50400
rect 163080 50400 163240 50560
rect 163080 50560 163240 50720
rect 163080 50720 163240 50880
rect 163080 50880 163240 51040
rect 163080 51040 163240 51200
rect 163080 51200 163240 51360
rect 163080 51360 163240 51520
rect 163080 51520 163240 51680
rect 163080 51680 163240 51840
rect 163080 51840 163240 52000
rect 163080 52000 163240 52160
rect 163080 52160 163240 52320
rect 163080 52320 163240 52480
rect 163080 52480 163240 52640
rect 163080 52640 163240 52800
rect 163240 27360 163400 27520
rect 163240 27520 163400 27680
rect 163240 27680 163400 27840
rect 163240 27840 163400 28000
rect 163240 28000 163400 28160
rect 163240 28160 163400 28320
rect 163240 28320 163400 28480
rect 163240 28480 163400 28640
rect 163240 28640 163400 28800
rect 163240 28800 163400 28960
rect 163240 28960 163400 29120
rect 163240 29120 163400 29280
rect 163240 29280 163400 29440
rect 163240 29440 163400 29600
rect 163240 29600 163400 29760
rect 163240 29760 163400 29920
rect 163240 29920 163400 30080
rect 163240 30080 163400 30240
rect 163240 30240 163400 30400
rect 163240 30400 163400 30560
rect 163240 30560 163400 30720
rect 163240 30720 163400 30880
rect 163240 30880 163400 31040
rect 163240 31040 163400 31200
rect 163240 31200 163400 31360
rect 163240 47680 163400 47840
rect 163240 47840 163400 48000
rect 163240 48000 163400 48160
rect 163240 48160 163400 48320
rect 163240 48320 163400 48480
rect 163240 48480 163400 48640
rect 163240 48640 163400 48800
rect 163240 48800 163400 48960
rect 163240 48960 163400 49120
rect 163240 49120 163400 49280
rect 163240 49280 163400 49440
rect 163240 49440 163400 49600
rect 163240 49600 163400 49760
rect 163240 49760 163400 49920
rect 163240 49920 163400 50080
rect 163240 50080 163400 50240
rect 163240 50240 163400 50400
rect 163240 50400 163400 50560
rect 163240 50560 163400 50720
rect 163240 50720 163400 50880
rect 163240 50880 163400 51040
rect 163240 51040 163400 51200
rect 163240 51200 163400 51360
rect 163240 51360 163400 51520
rect 163240 51520 163400 51680
rect 163240 51680 163400 51840
rect 163240 51840 163400 52000
rect 163240 52000 163400 52160
rect 163240 52160 163400 52320
rect 163240 52320 163400 52480
rect 163240 52480 163400 52640
rect 163240 52640 163400 52800
rect 163240 52800 163400 52960
rect 163400 27360 163560 27520
rect 163400 27520 163560 27680
rect 163400 27680 163560 27840
rect 163400 27840 163560 28000
rect 163400 28000 163560 28160
rect 163400 28160 163560 28320
rect 163400 28320 163560 28480
rect 163400 28480 163560 28640
rect 163400 28640 163560 28800
rect 163400 28800 163560 28960
rect 163400 28960 163560 29120
rect 163400 29120 163560 29280
rect 163400 29280 163560 29440
rect 163400 29440 163560 29600
rect 163400 29600 163560 29760
rect 163400 29760 163560 29920
rect 163400 29920 163560 30080
rect 163400 30080 163560 30240
rect 163400 30240 163560 30400
rect 163400 30400 163560 30560
rect 163400 30560 163560 30720
rect 163400 30720 163560 30880
rect 163400 30880 163560 31040
rect 163400 31040 163560 31200
rect 163400 31200 163560 31360
rect 163400 48000 163560 48160
rect 163400 48160 163560 48320
rect 163400 48320 163560 48480
rect 163400 48480 163560 48640
rect 163400 48640 163560 48800
rect 163400 48800 163560 48960
rect 163400 48960 163560 49120
rect 163400 49120 163560 49280
rect 163400 49280 163560 49440
rect 163400 49440 163560 49600
rect 163400 49600 163560 49760
rect 163400 49760 163560 49920
rect 163400 49920 163560 50080
rect 163400 50080 163560 50240
rect 163400 50240 163560 50400
rect 163400 50400 163560 50560
rect 163400 50560 163560 50720
rect 163400 50720 163560 50880
rect 163400 50880 163560 51040
rect 163400 51040 163560 51200
rect 163400 51200 163560 51360
rect 163400 51360 163560 51520
rect 163400 51520 163560 51680
rect 163400 51680 163560 51840
rect 163400 51840 163560 52000
rect 163400 52000 163560 52160
rect 163400 52160 163560 52320
rect 163400 52320 163560 52480
rect 163400 52480 163560 52640
rect 163400 52640 163560 52800
rect 163400 52800 163560 52960
rect 163560 27200 163720 27360
rect 163560 27360 163720 27520
rect 163560 27520 163720 27680
rect 163560 27680 163720 27840
rect 163560 27840 163720 28000
rect 163560 28000 163720 28160
rect 163560 28160 163720 28320
rect 163560 28320 163720 28480
rect 163560 28480 163720 28640
rect 163560 28640 163720 28800
rect 163560 28800 163720 28960
rect 163560 28960 163720 29120
rect 163560 29120 163720 29280
rect 163560 29280 163720 29440
rect 163560 29440 163720 29600
rect 163560 29600 163720 29760
rect 163560 29760 163720 29920
rect 163560 29920 163720 30080
rect 163560 30080 163720 30240
rect 163560 30240 163720 30400
rect 163560 30400 163720 30560
rect 163560 30560 163720 30720
rect 163560 30720 163720 30880
rect 163560 30880 163720 31040
rect 163560 31040 163720 31200
rect 163560 48160 163720 48320
rect 163560 48320 163720 48480
rect 163560 48480 163720 48640
rect 163560 48640 163720 48800
rect 163560 48800 163720 48960
rect 163560 48960 163720 49120
rect 163560 49120 163720 49280
rect 163560 49280 163720 49440
rect 163560 49440 163720 49600
rect 163560 49600 163720 49760
rect 163560 49760 163720 49920
rect 163560 49920 163720 50080
rect 163560 50080 163720 50240
rect 163560 50240 163720 50400
rect 163560 50400 163720 50560
rect 163560 50560 163720 50720
rect 163560 50720 163720 50880
rect 163560 50880 163720 51040
rect 163560 51040 163720 51200
rect 163560 51200 163720 51360
rect 163560 51360 163720 51520
rect 163560 51520 163720 51680
rect 163560 51680 163720 51840
rect 163560 51840 163720 52000
rect 163560 52000 163720 52160
rect 163560 52160 163720 52320
rect 163560 52320 163720 52480
rect 163560 52480 163720 52640
rect 163560 52640 163720 52800
rect 163560 52800 163720 52960
rect 163560 52960 163720 53120
rect 163720 27200 163880 27360
rect 163720 27360 163880 27520
rect 163720 27520 163880 27680
rect 163720 27680 163880 27840
rect 163720 27840 163880 28000
rect 163720 28000 163880 28160
rect 163720 28160 163880 28320
rect 163720 28320 163880 28480
rect 163720 28480 163880 28640
rect 163720 28640 163880 28800
rect 163720 28800 163880 28960
rect 163720 28960 163880 29120
rect 163720 29120 163880 29280
rect 163720 29280 163880 29440
rect 163720 29440 163880 29600
rect 163720 29600 163880 29760
rect 163720 29760 163880 29920
rect 163720 29920 163880 30080
rect 163720 30080 163880 30240
rect 163720 30240 163880 30400
rect 163720 30400 163880 30560
rect 163720 30560 163880 30720
rect 163720 30720 163880 30880
rect 163720 30880 163880 31040
rect 163720 48320 163880 48480
rect 163720 48480 163880 48640
rect 163720 48640 163880 48800
rect 163720 48800 163880 48960
rect 163720 48960 163880 49120
rect 163720 49120 163880 49280
rect 163720 49280 163880 49440
rect 163720 49440 163880 49600
rect 163720 49600 163880 49760
rect 163720 49760 163880 49920
rect 163720 49920 163880 50080
rect 163720 50080 163880 50240
rect 163720 50240 163880 50400
rect 163720 50400 163880 50560
rect 163720 50560 163880 50720
rect 163720 50720 163880 50880
rect 163720 50880 163880 51040
rect 163720 51040 163880 51200
rect 163720 51200 163880 51360
rect 163720 51360 163880 51520
rect 163720 51520 163880 51680
rect 163720 51680 163880 51840
rect 163720 51840 163880 52000
rect 163720 52000 163880 52160
rect 163720 52160 163880 52320
rect 163720 52320 163880 52480
rect 163720 52480 163880 52640
rect 163720 52640 163880 52800
rect 163720 52800 163880 52960
rect 163720 52960 163880 53120
rect 163880 27200 164040 27360
rect 163880 27360 164040 27520
rect 163880 27520 164040 27680
rect 163880 27680 164040 27840
rect 163880 27840 164040 28000
rect 163880 28000 164040 28160
rect 163880 28160 164040 28320
rect 163880 28320 164040 28480
rect 163880 28480 164040 28640
rect 163880 28640 164040 28800
rect 163880 28800 164040 28960
rect 163880 28960 164040 29120
rect 163880 29120 164040 29280
rect 163880 29280 164040 29440
rect 163880 29440 164040 29600
rect 163880 29600 164040 29760
rect 163880 29760 164040 29920
rect 163880 29920 164040 30080
rect 163880 30080 164040 30240
rect 163880 30240 164040 30400
rect 163880 30400 164040 30560
rect 163880 30560 164040 30720
rect 163880 30720 164040 30880
rect 163880 30880 164040 31040
rect 163880 48480 164040 48640
rect 163880 48640 164040 48800
rect 163880 48800 164040 48960
rect 163880 48960 164040 49120
rect 163880 49120 164040 49280
rect 163880 49280 164040 49440
rect 163880 49440 164040 49600
rect 163880 49600 164040 49760
rect 163880 49760 164040 49920
rect 163880 49920 164040 50080
rect 163880 50080 164040 50240
rect 163880 50240 164040 50400
rect 163880 50400 164040 50560
rect 163880 50560 164040 50720
rect 163880 50720 164040 50880
rect 163880 50880 164040 51040
rect 163880 51040 164040 51200
rect 163880 51200 164040 51360
rect 163880 51360 164040 51520
rect 163880 51520 164040 51680
rect 163880 51680 164040 51840
rect 163880 51840 164040 52000
rect 163880 52000 164040 52160
rect 163880 52160 164040 52320
rect 163880 52320 164040 52480
rect 163880 52480 164040 52640
rect 163880 52640 164040 52800
rect 163880 52800 164040 52960
rect 163880 52960 164040 53120
rect 164040 27040 164200 27200
rect 164040 27200 164200 27360
rect 164040 27360 164200 27520
rect 164040 27520 164200 27680
rect 164040 27680 164200 27840
rect 164040 27840 164200 28000
rect 164040 28000 164200 28160
rect 164040 28160 164200 28320
rect 164040 28320 164200 28480
rect 164040 28480 164200 28640
rect 164040 28640 164200 28800
rect 164040 28800 164200 28960
rect 164040 28960 164200 29120
rect 164040 29120 164200 29280
rect 164040 29280 164200 29440
rect 164040 29440 164200 29600
rect 164040 29600 164200 29760
rect 164040 29760 164200 29920
rect 164040 29920 164200 30080
rect 164040 30080 164200 30240
rect 164040 30240 164200 30400
rect 164040 30400 164200 30560
rect 164040 30560 164200 30720
rect 164040 30720 164200 30880
rect 164040 48800 164200 48960
rect 164040 48960 164200 49120
rect 164040 49120 164200 49280
rect 164040 49280 164200 49440
rect 164040 49440 164200 49600
rect 164040 49600 164200 49760
rect 164040 49760 164200 49920
rect 164040 49920 164200 50080
rect 164040 50080 164200 50240
rect 164040 50240 164200 50400
rect 164040 50400 164200 50560
rect 164040 50560 164200 50720
rect 164040 50720 164200 50880
rect 164040 50880 164200 51040
rect 164040 51040 164200 51200
rect 164040 51200 164200 51360
rect 164040 51360 164200 51520
rect 164040 51520 164200 51680
rect 164040 51680 164200 51840
rect 164040 51840 164200 52000
rect 164040 52000 164200 52160
rect 164040 52160 164200 52320
rect 164040 52320 164200 52480
rect 164040 52480 164200 52640
rect 164040 52640 164200 52800
rect 164040 52800 164200 52960
rect 164040 52960 164200 53120
rect 164200 27040 164360 27200
rect 164200 27200 164360 27360
rect 164200 27360 164360 27520
rect 164200 27520 164360 27680
rect 164200 27680 164360 27840
rect 164200 27840 164360 28000
rect 164200 28000 164360 28160
rect 164200 28160 164360 28320
rect 164200 28320 164360 28480
rect 164200 28480 164360 28640
rect 164200 28640 164360 28800
rect 164200 28800 164360 28960
rect 164200 28960 164360 29120
rect 164200 29120 164360 29280
rect 164200 29280 164360 29440
rect 164200 29440 164360 29600
rect 164200 29600 164360 29760
rect 164200 29760 164360 29920
rect 164200 29920 164360 30080
rect 164200 30080 164360 30240
rect 164200 30240 164360 30400
rect 164200 30400 164360 30560
rect 164200 30560 164360 30720
rect 164200 30720 164360 30880
rect 164200 48960 164360 49120
rect 164200 49120 164360 49280
rect 164200 49280 164360 49440
rect 164200 49440 164360 49600
rect 164200 49600 164360 49760
rect 164200 49760 164360 49920
rect 164200 49920 164360 50080
rect 164200 50080 164360 50240
rect 164200 50240 164360 50400
rect 164200 50400 164360 50560
rect 164200 50560 164360 50720
rect 164200 50720 164360 50880
rect 164200 50880 164360 51040
rect 164200 51040 164360 51200
rect 164200 51200 164360 51360
rect 164200 51360 164360 51520
rect 164200 51520 164360 51680
rect 164200 51680 164360 51840
rect 164200 51840 164360 52000
rect 164200 52000 164360 52160
rect 164200 52160 164360 52320
rect 164200 52320 164360 52480
rect 164200 52480 164360 52640
rect 164200 52640 164360 52800
rect 164200 52800 164360 52960
rect 164360 27040 164520 27200
rect 164360 27200 164520 27360
rect 164360 27360 164520 27520
rect 164360 27520 164520 27680
rect 164360 27680 164520 27840
rect 164360 27840 164520 28000
rect 164360 28000 164520 28160
rect 164360 28160 164520 28320
rect 164360 28320 164520 28480
rect 164360 28480 164520 28640
rect 164360 28640 164520 28800
rect 164360 28800 164520 28960
rect 164360 28960 164520 29120
rect 164360 29120 164520 29280
rect 164360 29280 164520 29440
rect 164360 29440 164520 29600
rect 164360 29600 164520 29760
rect 164360 29760 164520 29920
rect 164360 29920 164520 30080
rect 164360 30080 164520 30240
rect 164360 30240 164520 30400
rect 164360 30400 164520 30560
rect 164360 30560 164520 30720
rect 164360 49120 164520 49280
rect 164360 49280 164520 49440
rect 164360 49440 164520 49600
rect 164360 49600 164520 49760
rect 164360 49760 164520 49920
rect 164360 49920 164520 50080
rect 164360 50080 164520 50240
rect 164360 50240 164520 50400
rect 164360 50400 164520 50560
rect 164360 50560 164520 50720
rect 164360 50720 164520 50880
rect 164360 50880 164520 51040
rect 164360 51040 164520 51200
rect 164360 51200 164520 51360
rect 164360 51360 164520 51520
rect 164360 51520 164520 51680
rect 164360 51680 164520 51840
rect 164360 51840 164520 52000
rect 164360 52000 164520 52160
rect 164360 52160 164520 52320
rect 164360 52320 164520 52480
rect 164360 52480 164520 52640
rect 164360 52640 164520 52800
rect 164360 52800 164520 52960
rect 164520 27040 164680 27200
rect 164520 27200 164680 27360
rect 164520 27360 164680 27520
rect 164520 27520 164680 27680
rect 164520 27680 164680 27840
rect 164520 27840 164680 28000
rect 164520 28000 164680 28160
rect 164520 28160 164680 28320
rect 164520 28320 164680 28480
rect 164520 28480 164680 28640
rect 164520 28640 164680 28800
rect 164520 28800 164680 28960
rect 164520 28960 164680 29120
rect 164520 29120 164680 29280
rect 164520 29280 164680 29440
rect 164520 29440 164680 29600
rect 164520 29600 164680 29760
rect 164520 29760 164680 29920
rect 164520 29920 164680 30080
rect 164520 30080 164680 30240
rect 164520 30240 164680 30400
rect 164520 30400 164680 30560
rect 164520 30560 164680 30720
rect 164520 49440 164680 49600
rect 164520 49600 164680 49760
rect 164520 49760 164680 49920
rect 164520 49920 164680 50080
rect 164520 50080 164680 50240
rect 164520 50240 164680 50400
rect 164520 50400 164680 50560
rect 164520 50560 164680 50720
rect 164520 50720 164680 50880
rect 164520 50880 164680 51040
rect 164520 51040 164680 51200
rect 164520 51200 164680 51360
rect 164520 51360 164680 51520
rect 164520 51520 164680 51680
rect 164520 51680 164680 51840
rect 164520 51840 164680 52000
rect 164520 52000 164680 52160
rect 164520 52160 164680 52320
rect 164520 52320 164680 52480
rect 164520 52480 164680 52640
rect 164520 52640 164680 52800
rect 164520 52800 164680 52960
rect 164680 27040 164840 27200
rect 164680 27200 164840 27360
rect 164680 27360 164840 27520
rect 164680 27520 164840 27680
rect 164680 27680 164840 27840
rect 164680 27840 164840 28000
rect 164680 28000 164840 28160
rect 164680 28160 164840 28320
rect 164680 28320 164840 28480
rect 164680 28480 164840 28640
rect 164680 28640 164840 28800
rect 164680 28800 164840 28960
rect 164680 28960 164840 29120
rect 164680 29120 164840 29280
rect 164680 29280 164840 29440
rect 164680 29440 164840 29600
rect 164680 29600 164840 29760
rect 164680 29760 164840 29920
rect 164680 29920 164840 30080
rect 164680 30080 164840 30240
rect 164680 30240 164840 30400
rect 164680 30400 164840 30560
rect 164680 49600 164840 49760
rect 164680 49760 164840 49920
rect 164680 49920 164840 50080
rect 164680 50080 164840 50240
rect 164680 50240 164840 50400
rect 164680 50400 164840 50560
rect 164680 50560 164840 50720
rect 164680 50720 164840 50880
rect 164680 50880 164840 51040
rect 164680 51040 164840 51200
rect 164680 51200 164840 51360
rect 164680 51360 164840 51520
rect 164680 51520 164840 51680
rect 164680 51680 164840 51840
rect 164680 51840 164840 52000
rect 164680 52000 164840 52160
rect 164680 52160 164840 52320
rect 164680 52320 164840 52480
rect 164680 52480 164840 52640
rect 164680 52640 164840 52800
rect 164840 27040 165000 27200
rect 164840 27200 165000 27360
rect 164840 27360 165000 27520
rect 164840 27520 165000 27680
rect 164840 27680 165000 27840
rect 164840 27840 165000 28000
rect 164840 28000 165000 28160
rect 164840 28160 165000 28320
rect 164840 28320 165000 28480
rect 164840 28480 165000 28640
rect 164840 28640 165000 28800
rect 164840 28800 165000 28960
rect 164840 28960 165000 29120
rect 164840 29120 165000 29280
rect 164840 29280 165000 29440
rect 164840 29440 165000 29600
rect 164840 29600 165000 29760
rect 164840 29760 165000 29920
rect 164840 29920 165000 30080
rect 164840 30080 165000 30240
rect 164840 30240 165000 30400
rect 164840 30400 165000 30560
rect 164840 49760 165000 49920
rect 164840 49920 165000 50080
rect 164840 50080 165000 50240
rect 164840 50240 165000 50400
rect 164840 50400 165000 50560
rect 164840 50560 165000 50720
rect 164840 50720 165000 50880
rect 164840 50880 165000 51040
rect 164840 51040 165000 51200
rect 164840 51200 165000 51360
rect 164840 51360 165000 51520
rect 164840 51520 165000 51680
rect 164840 51680 165000 51840
rect 164840 51840 165000 52000
rect 164840 52000 165000 52160
rect 164840 52160 165000 52320
rect 164840 52320 165000 52480
rect 164840 52480 165000 52640
rect 164840 52640 165000 52800
rect 165000 27040 165160 27200
rect 165000 27200 165160 27360
rect 165000 27360 165160 27520
rect 165000 27520 165160 27680
rect 165000 27680 165160 27840
rect 165000 27840 165160 28000
rect 165000 28000 165160 28160
rect 165000 28160 165160 28320
rect 165000 28320 165160 28480
rect 165000 28480 165160 28640
rect 165000 28640 165160 28800
rect 165000 28800 165160 28960
rect 165000 28960 165160 29120
rect 165000 29120 165160 29280
rect 165000 29280 165160 29440
rect 165000 29440 165160 29600
rect 165000 29600 165160 29760
rect 165000 29760 165160 29920
rect 165000 29920 165160 30080
rect 165000 30080 165160 30240
rect 165000 30240 165160 30400
rect 165000 50080 165160 50240
rect 165000 50240 165160 50400
rect 165000 50400 165160 50560
rect 165000 50560 165160 50720
rect 165000 50720 165160 50880
rect 165000 50880 165160 51040
rect 165000 51040 165160 51200
rect 165000 51200 165160 51360
rect 165000 51360 165160 51520
rect 165000 51520 165160 51680
rect 165000 51680 165160 51840
rect 165000 51840 165160 52000
rect 165000 52000 165160 52160
rect 165000 52160 165160 52320
rect 165000 52320 165160 52480
rect 165000 52480 165160 52640
rect 165160 27040 165320 27200
rect 165160 27200 165320 27360
rect 165160 27360 165320 27520
rect 165160 27520 165320 27680
rect 165160 27680 165320 27840
rect 165160 27840 165320 28000
rect 165160 28000 165320 28160
rect 165160 28160 165320 28320
rect 165160 28320 165320 28480
rect 165160 28480 165320 28640
rect 165160 28640 165320 28800
rect 165160 28800 165320 28960
rect 165160 28960 165320 29120
rect 165160 29120 165320 29280
rect 165160 29280 165320 29440
rect 165160 29440 165320 29600
rect 165160 29600 165320 29760
rect 165160 29760 165320 29920
rect 165160 29920 165320 30080
rect 165160 30080 165320 30240
rect 165160 30240 165320 30400
rect 165160 50400 165320 50560
rect 165160 50560 165320 50720
rect 165160 50720 165320 50880
rect 165160 50880 165320 51040
rect 165160 51040 165320 51200
rect 165160 51200 165320 51360
rect 165160 51360 165320 51520
rect 165160 51520 165320 51680
rect 165160 51680 165320 51840
rect 165160 51840 165320 52000
rect 165160 52000 165320 52160
rect 165160 52160 165320 52320
rect 165160 52320 165320 52480
rect 165320 27040 165480 27200
rect 165320 27200 165480 27360
rect 165320 27360 165480 27520
rect 165320 27520 165480 27680
rect 165320 27680 165480 27840
rect 165320 27840 165480 28000
rect 165320 28000 165480 28160
rect 165320 28160 165480 28320
rect 165320 28320 165480 28480
rect 165320 28480 165480 28640
rect 165320 28640 165480 28800
rect 165320 28800 165480 28960
rect 165320 28960 165480 29120
rect 165320 29120 165480 29280
rect 165320 29280 165480 29440
rect 165320 29440 165480 29600
rect 165320 29600 165480 29760
rect 165320 29760 165480 29920
rect 165320 29920 165480 30080
rect 165320 30080 165480 30240
rect 165320 30240 165480 30400
rect 165320 50560 165480 50720
rect 165320 50720 165480 50880
rect 165320 50880 165480 51040
rect 165320 51040 165480 51200
rect 165320 51200 165480 51360
rect 165320 51360 165480 51520
rect 165320 51520 165480 51680
rect 165320 51680 165480 51840
rect 165320 51840 165480 52000
rect 165320 52000 165480 52160
rect 165480 27040 165640 27200
rect 165480 27200 165640 27360
rect 165480 27360 165640 27520
rect 165480 27520 165640 27680
rect 165480 27680 165640 27840
rect 165480 27840 165640 28000
rect 165480 28000 165640 28160
rect 165480 28160 165640 28320
rect 165480 28320 165640 28480
rect 165480 28480 165640 28640
rect 165480 28640 165640 28800
rect 165480 28800 165640 28960
rect 165480 28960 165640 29120
rect 165480 29120 165640 29280
rect 165480 29280 165640 29440
rect 165480 29440 165640 29600
rect 165480 29600 165640 29760
rect 165480 29760 165640 29920
rect 165480 29920 165640 30080
rect 165480 30080 165640 30240
rect 165480 51040 165640 51200
rect 165480 51200 165640 51360
rect 165480 51360 165640 51520
rect 165480 51520 165640 51680
rect 165480 51680 165640 51840
rect 165640 27200 165800 27360
rect 165640 27360 165800 27520
rect 165640 27520 165800 27680
rect 165640 27680 165800 27840
rect 165640 27840 165800 28000
rect 165640 28000 165800 28160
rect 165640 28160 165800 28320
rect 165640 28320 165800 28480
rect 165640 28480 165800 28640
rect 165640 28640 165800 28800
rect 165640 28800 165800 28960
rect 165640 28960 165800 29120
rect 165640 29120 165800 29280
rect 165640 29280 165800 29440
rect 165640 29440 165800 29600
rect 165640 29600 165800 29760
rect 165640 29760 165800 29920
rect 165640 29920 165800 30080
rect 165640 30080 165800 30240
rect 165800 27200 165960 27360
rect 165800 27360 165960 27520
rect 165800 27520 165960 27680
rect 165800 27680 165960 27840
rect 165800 27840 165960 28000
rect 165800 28000 165960 28160
rect 165800 28160 165960 28320
rect 165800 28320 165960 28480
rect 165800 28480 165960 28640
rect 165800 28640 165960 28800
rect 165800 28800 165960 28960
rect 165800 28960 165960 29120
rect 165800 29120 165960 29280
rect 165800 29280 165960 29440
rect 165800 29440 165960 29600
rect 165800 29600 165960 29760
rect 165800 29760 165960 29920
rect 165800 29920 165960 30080
rect 165960 27360 166120 27520
rect 165960 27520 166120 27680
rect 165960 27680 166120 27840
rect 165960 27840 166120 28000
rect 165960 28000 166120 28160
rect 165960 28160 166120 28320
rect 165960 28320 166120 28480
rect 165960 28480 166120 28640
rect 165960 28640 166120 28800
rect 165960 28800 166120 28960
rect 165960 28960 166120 29120
rect 165960 29120 166120 29280
rect 165960 29280 166120 29440
rect 165960 29440 166120 29600
rect 165960 29600 166120 29760
rect 165960 29760 166120 29920
rect 166120 27520 166280 27680
rect 166120 27680 166280 27840
rect 166120 27840 166280 28000
rect 166120 28000 166280 28160
rect 166120 28160 166280 28320
rect 166120 28320 166280 28480
rect 166120 28480 166280 28640
rect 166120 28640 166280 28800
rect 166120 28800 166280 28960
rect 166120 28960 166280 29120
rect 166120 29120 166280 29280
rect 166120 29280 166280 29440
rect 166120 29440 166280 29600
rect 166120 29600 166280 29760
rect 166280 27840 166440 28000
rect 166280 28000 166440 28160
rect 166280 28160 166440 28320
rect 166280 28320 166440 28480
rect 166280 28480 166440 28640
rect 166280 28640 166440 28800
rect 166280 28800 166440 28960
rect 166280 28960 166440 29120
rect 166280 29120 166440 29280
rect 166280 29280 166440 29440
rect 166280 29440 166440 29600
rect 166440 28160 166600 28320
rect 166440 28320 166600 28480
rect 166440 28480 166600 28640
rect 166440 28640 166600 28800
rect 166440 28800 166600 28960
rect 166440 28960 166600 29120
rect 166440 29120 166600 29280
rect 169000 51520 169160 51680
rect 169000 51840 169160 52000
rect 169160 50880 169320 51040
rect 169160 51040 169320 51200
rect 169160 51200 169320 51360
rect 169160 51360 169320 51520
rect 169160 51520 169320 51680
rect 169160 51680 169320 51840
rect 169160 51840 169320 52000
rect 169160 52000 169320 52160
rect 169160 52160 169320 52320
rect 169160 52320 169320 52480
rect 169320 50400 169480 50560
rect 169320 50560 169480 50720
rect 169320 50720 169480 50880
rect 169320 50880 169480 51040
rect 169320 51040 169480 51200
rect 169320 51200 169480 51360
rect 169320 51360 169480 51520
rect 169320 51520 169480 51680
rect 169320 51680 169480 51840
rect 169320 51840 169480 52000
rect 169320 52000 169480 52160
rect 169320 52160 169480 52320
rect 169320 52320 169480 52480
rect 169320 52480 169480 52640
rect 169320 52640 169480 52800
rect 169480 49920 169640 50080
rect 169480 50080 169640 50240
rect 169480 50240 169640 50400
rect 169480 50400 169640 50560
rect 169480 50560 169640 50720
rect 169480 50720 169640 50880
rect 169480 50880 169640 51040
rect 169480 51040 169640 51200
rect 169480 51200 169640 51360
rect 169480 51360 169640 51520
rect 169480 51520 169640 51680
rect 169480 51680 169640 51840
rect 169480 51840 169640 52000
rect 169480 52000 169640 52160
rect 169480 52160 169640 52320
rect 169480 52320 169640 52480
rect 169480 52480 169640 52640
rect 169480 52640 169640 52800
rect 169480 52800 169640 52960
rect 169640 49440 169800 49600
rect 169640 49600 169800 49760
rect 169640 49760 169800 49920
rect 169640 49920 169800 50080
rect 169640 50080 169800 50240
rect 169640 50240 169800 50400
rect 169640 50400 169800 50560
rect 169640 50560 169800 50720
rect 169640 50720 169800 50880
rect 169640 50880 169800 51040
rect 169640 51040 169800 51200
rect 169640 51200 169800 51360
rect 169640 51360 169800 51520
rect 169640 51520 169800 51680
rect 169640 51680 169800 51840
rect 169640 51840 169800 52000
rect 169640 52000 169800 52160
rect 169640 52160 169800 52320
rect 169640 52320 169800 52480
rect 169640 52480 169800 52640
rect 169640 52640 169800 52800
rect 169640 52800 169800 52960
rect 169800 48960 169960 49120
rect 169800 49120 169960 49280
rect 169800 49280 169960 49440
rect 169800 49440 169960 49600
rect 169800 49600 169960 49760
rect 169800 49760 169960 49920
rect 169800 49920 169960 50080
rect 169800 50080 169960 50240
rect 169800 50240 169960 50400
rect 169800 50400 169960 50560
rect 169800 50560 169960 50720
rect 169800 50720 169960 50880
rect 169800 50880 169960 51040
rect 169800 51040 169960 51200
rect 169800 51200 169960 51360
rect 169800 51360 169960 51520
rect 169800 51520 169960 51680
rect 169800 51680 169960 51840
rect 169800 51840 169960 52000
rect 169800 52000 169960 52160
rect 169800 52160 169960 52320
rect 169800 52320 169960 52480
rect 169800 52480 169960 52640
rect 169800 52640 169960 52800
rect 169800 52800 169960 52960
rect 169800 52960 169960 53120
rect 169960 48480 170120 48640
rect 169960 48640 170120 48800
rect 169960 48800 170120 48960
rect 169960 48960 170120 49120
rect 169960 49120 170120 49280
rect 169960 49280 170120 49440
rect 169960 49440 170120 49600
rect 169960 49600 170120 49760
rect 169960 49760 170120 49920
rect 169960 49920 170120 50080
rect 169960 50080 170120 50240
rect 169960 50240 170120 50400
rect 169960 50400 170120 50560
rect 169960 50560 170120 50720
rect 169960 50720 170120 50880
rect 169960 50880 170120 51040
rect 169960 51040 170120 51200
rect 169960 51200 170120 51360
rect 169960 51360 170120 51520
rect 169960 51520 170120 51680
rect 169960 51680 170120 51840
rect 169960 51840 170120 52000
rect 169960 52000 170120 52160
rect 169960 52160 170120 52320
rect 169960 52320 170120 52480
rect 169960 52480 170120 52640
rect 169960 52640 170120 52800
rect 169960 52800 170120 52960
rect 169960 52960 170120 53120
rect 170120 48000 170280 48160
rect 170120 48160 170280 48320
rect 170120 48320 170280 48480
rect 170120 48480 170280 48640
rect 170120 48640 170280 48800
rect 170120 48800 170280 48960
rect 170120 48960 170280 49120
rect 170120 49120 170280 49280
rect 170120 49280 170280 49440
rect 170120 49440 170280 49600
rect 170120 49600 170280 49760
rect 170120 49760 170280 49920
rect 170120 49920 170280 50080
rect 170120 50080 170280 50240
rect 170120 50240 170280 50400
rect 170120 50400 170280 50560
rect 170120 50560 170280 50720
rect 170120 50720 170280 50880
rect 170120 50880 170280 51040
rect 170120 51040 170280 51200
rect 170120 51200 170280 51360
rect 170120 51360 170280 51520
rect 170120 51520 170280 51680
rect 170120 51680 170280 51840
rect 170120 51840 170280 52000
rect 170120 52000 170280 52160
rect 170120 52160 170280 52320
rect 170120 52320 170280 52480
rect 170120 52480 170280 52640
rect 170120 52640 170280 52800
rect 170120 52800 170280 52960
rect 170120 52960 170280 53120
rect 170120 53120 170280 53280
rect 170280 47520 170440 47680
rect 170280 47680 170440 47840
rect 170280 47840 170440 48000
rect 170280 48000 170440 48160
rect 170280 48160 170440 48320
rect 170280 48320 170440 48480
rect 170280 48480 170440 48640
rect 170280 48640 170440 48800
rect 170280 48800 170440 48960
rect 170280 48960 170440 49120
rect 170280 49120 170440 49280
rect 170280 49280 170440 49440
rect 170280 49440 170440 49600
rect 170280 49600 170440 49760
rect 170280 49760 170440 49920
rect 170280 49920 170440 50080
rect 170280 50080 170440 50240
rect 170280 50240 170440 50400
rect 170280 50400 170440 50560
rect 170280 50560 170440 50720
rect 170280 50720 170440 50880
rect 170280 50880 170440 51040
rect 170280 51040 170440 51200
rect 170280 51200 170440 51360
rect 170280 51360 170440 51520
rect 170280 51520 170440 51680
rect 170280 51680 170440 51840
rect 170280 51840 170440 52000
rect 170280 52000 170440 52160
rect 170280 52160 170440 52320
rect 170280 52320 170440 52480
rect 170280 52480 170440 52640
rect 170280 52640 170440 52800
rect 170280 52800 170440 52960
rect 170280 52960 170440 53120
rect 170280 53120 170440 53280
rect 170440 47040 170600 47200
rect 170440 47200 170600 47360
rect 170440 47360 170600 47520
rect 170440 47520 170600 47680
rect 170440 47680 170600 47840
rect 170440 47840 170600 48000
rect 170440 48000 170600 48160
rect 170440 48160 170600 48320
rect 170440 48320 170600 48480
rect 170440 48480 170600 48640
rect 170440 48640 170600 48800
rect 170440 48800 170600 48960
rect 170440 48960 170600 49120
rect 170440 49120 170600 49280
rect 170440 49280 170600 49440
rect 170440 49440 170600 49600
rect 170440 49600 170600 49760
rect 170440 49760 170600 49920
rect 170440 49920 170600 50080
rect 170440 50080 170600 50240
rect 170440 50240 170600 50400
rect 170440 50400 170600 50560
rect 170440 50560 170600 50720
rect 170440 50720 170600 50880
rect 170440 50880 170600 51040
rect 170440 51040 170600 51200
rect 170440 51200 170600 51360
rect 170440 51360 170600 51520
rect 170440 51520 170600 51680
rect 170440 51680 170600 51840
rect 170440 51840 170600 52000
rect 170440 52000 170600 52160
rect 170440 52160 170600 52320
rect 170440 52320 170600 52480
rect 170440 52480 170600 52640
rect 170440 52640 170600 52800
rect 170440 52800 170600 52960
rect 170440 52960 170600 53120
rect 170440 53120 170600 53280
rect 170600 46560 170760 46720
rect 170600 46720 170760 46880
rect 170600 46880 170760 47040
rect 170600 47040 170760 47200
rect 170600 47200 170760 47360
rect 170600 47360 170760 47520
rect 170600 47520 170760 47680
rect 170600 47680 170760 47840
rect 170600 47840 170760 48000
rect 170600 48000 170760 48160
rect 170600 48160 170760 48320
rect 170600 48320 170760 48480
rect 170600 48480 170760 48640
rect 170600 48640 170760 48800
rect 170600 48800 170760 48960
rect 170600 48960 170760 49120
rect 170600 49120 170760 49280
rect 170600 49280 170760 49440
rect 170600 49440 170760 49600
rect 170600 49600 170760 49760
rect 170600 49760 170760 49920
rect 170600 49920 170760 50080
rect 170600 50080 170760 50240
rect 170600 50240 170760 50400
rect 170600 50400 170760 50560
rect 170600 50560 170760 50720
rect 170600 50720 170760 50880
rect 170600 50880 170760 51040
rect 170600 51040 170760 51200
rect 170600 51200 170760 51360
rect 170600 51360 170760 51520
rect 170600 51520 170760 51680
rect 170600 51680 170760 51840
rect 170600 51840 170760 52000
rect 170600 52000 170760 52160
rect 170600 52160 170760 52320
rect 170600 52320 170760 52480
rect 170600 52480 170760 52640
rect 170600 52640 170760 52800
rect 170600 52800 170760 52960
rect 170600 52960 170760 53120
rect 170600 53120 170760 53280
rect 170760 46080 170920 46240
rect 170760 46240 170920 46400
rect 170760 46400 170920 46560
rect 170760 46560 170920 46720
rect 170760 46720 170920 46880
rect 170760 46880 170920 47040
rect 170760 47040 170920 47200
rect 170760 47200 170920 47360
rect 170760 47360 170920 47520
rect 170760 47520 170920 47680
rect 170760 47680 170920 47840
rect 170760 47840 170920 48000
rect 170760 48000 170920 48160
rect 170760 48160 170920 48320
rect 170760 48320 170920 48480
rect 170760 48480 170920 48640
rect 170760 48640 170920 48800
rect 170760 48800 170920 48960
rect 170760 48960 170920 49120
rect 170760 49120 170920 49280
rect 170760 49280 170920 49440
rect 170760 49440 170920 49600
rect 170760 49600 170920 49760
rect 170760 49760 170920 49920
rect 170760 49920 170920 50080
rect 170760 50080 170920 50240
rect 170760 50240 170920 50400
rect 170760 50400 170920 50560
rect 170760 50560 170920 50720
rect 170760 50720 170920 50880
rect 170760 50880 170920 51040
rect 170760 51040 170920 51200
rect 170760 51200 170920 51360
rect 170760 51360 170920 51520
rect 170760 51520 170920 51680
rect 170760 51680 170920 51840
rect 170760 51840 170920 52000
rect 170760 52000 170920 52160
rect 170760 52160 170920 52320
rect 170760 52320 170920 52480
rect 170760 52480 170920 52640
rect 170760 52640 170920 52800
rect 170760 52800 170920 52960
rect 170760 52960 170920 53120
rect 170760 53120 170920 53280
rect 170920 45600 171080 45760
rect 170920 45760 171080 45920
rect 170920 45920 171080 46080
rect 170920 46080 171080 46240
rect 170920 46240 171080 46400
rect 170920 46400 171080 46560
rect 170920 46560 171080 46720
rect 170920 46720 171080 46880
rect 170920 46880 171080 47040
rect 170920 47040 171080 47200
rect 170920 47200 171080 47360
rect 170920 47360 171080 47520
rect 170920 47520 171080 47680
rect 170920 47680 171080 47840
rect 170920 47840 171080 48000
rect 170920 48000 171080 48160
rect 170920 48160 171080 48320
rect 170920 48320 171080 48480
rect 170920 48480 171080 48640
rect 170920 48640 171080 48800
rect 170920 48800 171080 48960
rect 170920 48960 171080 49120
rect 170920 49120 171080 49280
rect 170920 49280 171080 49440
rect 170920 49440 171080 49600
rect 170920 49600 171080 49760
rect 170920 49760 171080 49920
rect 170920 49920 171080 50080
rect 170920 50080 171080 50240
rect 170920 50240 171080 50400
rect 170920 50400 171080 50560
rect 170920 50560 171080 50720
rect 170920 50720 171080 50880
rect 170920 50880 171080 51040
rect 170920 51040 171080 51200
rect 170920 51200 171080 51360
rect 170920 51360 171080 51520
rect 170920 51520 171080 51680
rect 170920 51680 171080 51840
rect 170920 51840 171080 52000
rect 170920 52000 171080 52160
rect 170920 52160 171080 52320
rect 170920 52320 171080 52480
rect 170920 52480 171080 52640
rect 170920 52640 171080 52800
rect 170920 52800 171080 52960
rect 170920 52960 171080 53120
rect 170920 53120 171080 53280
rect 171080 44960 171240 45120
rect 171080 45120 171240 45280
rect 171080 45280 171240 45440
rect 171080 45440 171240 45600
rect 171080 45600 171240 45760
rect 171080 45760 171240 45920
rect 171080 45920 171240 46080
rect 171080 46080 171240 46240
rect 171080 46240 171240 46400
rect 171080 46400 171240 46560
rect 171080 46560 171240 46720
rect 171080 46720 171240 46880
rect 171080 46880 171240 47040
rect 171080 47040 171240 47200
rect 171080 47200 171240 47360
rect 171080 47360 171240 47520
rect 171080 47520 171240 47680
rect 171080 47680 171240 47840
rect 171080 47840 171240 48000
rect 171080 48000 171240 48160
rect 171080 48160 171240 48320
rect 171080 48320 171240 48480
rect 171080 48480 171240 48640
rect 171080 48640 171240 48800
rect 171080 48800 171240 48960
rect 171080 48960 171240 49120
rect 171080 49120 171240 49280
rect 171080 49280 171240 49440
rect 171080 49440 171240 49600
rect 171080 49600 171240 49760
rect 171080 49760 171240 49920
rect 171080 49920 171240 50080
rect 171080 50080 171240 50240
rect 171080 50240 171240 50400
rect 171080 50400 171240 50560
rect 171080 50560 171240 50720
rect 171080 50720 171240 50880
rect 171080 50880 171240 51040
rect 171080 51040 171240 51200
rect 171080 51200 171240 51360
rect 171080 51360 171240 51520
rect 171080 51520 171240 51680
rect 171080 51680 171240 51840
rect 171080 51840 171240 52000
rect 171080 52000 171240 52160
rect 171080 52160 171240 52320
rect 171080 52320 171240 52480
rect 171080 52480 171240 52640
rect 171080 52640 171240 52800
rect 171080 52800 171240 52960
rect 171080 52960 171240 53120
rect 171080 53120 171240 53280
rect 171240 44480 171400 44640
rect 171240 44640 171400 44800
rect 171240 44800 171400 44960
rect 171240 44960 171400 45120
rect 171240 45120 171400 45280
rect 171240 45280 171400 45440
rect 171240 45440 171400 45600
rect 171240 45600 171400 45760
rect 171240 45760 171400 45920
rect 171240 45920 171400 46080
rect 171240 46080 171400 46240
rect 171240 46240 171400 46400
rect 171240 46400 171400 46560
rect 171240 46560 171400 46720
rect 171240 46720 171400 46880
rect 171240 46880 171400 47040
rect 171240 47040 171400 47200
rect 171240 47200 171400 47360
rect 171240 47360 171400 47520
rect 171240 47520 171400 47680
rect 171240 47680 171400 47840
rect 171240 47840 171400 48000
rect 171240 48000 171400 48160
rect 171240 48160 171400 48320
rect 171240 48320 171400 48480
rect 171240 48480 171400 48640
rect 171240 48640 171400 48800
rect 171240 48800 171400 48960
rect 171240 48960 171400 49120
rect 171240 49120 171400 49280
rect 171240 49280 171400 49440
rect 171240 49440 171400 49600
rect 171240 49600 171400 49760
rect 171240 49760 171400 49920
rect 171240 49920 171400 50080
rect 171240 50080 171400 50240
rect 171240 50240 171400 50400
rect 171240 50400 171400 50560
rect 171240 50560 171400 50720
rect 171240 50720 171400 50880
rect 171240 50880 171400 51040
rect 171240 51040 171400 51200
rect 171240 51200 171400 51360
rect 171240 51360 171400 51520
rect 171240 51520 171400 51680
rect 171240 51680 171400 51840
rect 171240 51840 171400 52000
rect 171240 52000 171400 52160
rect 171240 52160 171400 52320
rect 171240 52320 171400 52480
rect 171240 52480 171400 52640
rect 171240 52640 171400 52800
rect 171240 52800 171400 52960
rect 171240 52960 171400 53120
rect 171240 53120 171400 53280
rect 171400 44000 171560 44160
rect 171400 44160 171560 44320
rect 171400 44320 171560 44480
rect 171400 44480 171560 44640
rect 171400 44640 171560 44800
rect 171400 44800 171560 44960
rect 171400 44960 171560 45120
rect 171400 45120 171560 45280
rect 171400 45280 171560 45440
rect 171400 45440 171560 45600
rect 171400 45600 171560 45760
rect 171400 45760 171560 45920
rect 171400 45920 171560 46080
rect 171400 46080 171560 46240
rect 171400 46240 171560 46400
rect 171400 46400 171560 46560
rect 171400 46560 171560 46720
rect 171400 46720 171560 46880
rect 171400 46880 171560 47040
rect 171400 47040 171560 47200
rect 171400 47200 171560 47360
rect 171400 47360 171560 47520
rect 171400 47520 171560 47680
rect 171400 47680 171560 47840
rect 171400 47840 171560 48000
rect 171400 48000 171560 48160
rect 171400 48160 171560 48320
rect 171400 48320 171560 48480
rect 171400 48480 171560 48640
rect 171400 48640 171560 48800
rect 171400 48800 171560 48960
rect 171400 48960 171560 49120
rect 171400 49120 171560 49280
rect 171400 49280 171560 49440
rect 171400 49440 171560 49600
rect 171400 49600 171560 49760
rect 171400 49760 171560 49920
rect 171400 49920 171560 50080
rect 171400 50080 171560 50240
rect 171400 50240 171560 50400
rect 171400 50400 171560 50560
rect 171400 50560 171560 50720
rect 171400 50720 171560 50880
rect 171400 50880 171560 51040
rect 171400 51040 171560 51200
rect 171400 51200 171560 51360
rect 171400 51360 171560 51520
rect 171400 51520 171560 51680
rect 171400 51680 171560 51840
rect 171400 51840 171560 52000
rect 171400 52000 171560 52160
rect 171400 52160 171560 52320
rect 171400 52320 171560 52480
rect 171400 52480 171560 52640
rect 171400 52640 171560 52800
rect 171400 52800 171560 52960
rect 171400 52960 171560 53120
rect 171560 43520 171720 43680
rect 171560 43680 171720 43840
rect 171560 43840 171720 44000
rect 171560 44000 171720 44160
rect 171560 44160 171720 44320
rect 171560 44320 171720 44480
rect 171560 44480 171720 44640
rect 171560 44640 171720 44800
rect 171560 44800 171720 44960
rect 171560 44960 171720 45120
rect 171560 45120 171720 45280
rect 171560 45280 171720 45440
rect 171560 45440 171720 45600
rect 171560 45600 171720 45760
rect 171560 45760 171720 45920
rect 171560 45920 171720 46080
rect 171560 46080 171720 46240
rect 171560 46240 171720 46400
rect 171560 46400 171720 46560
rect 171560 46560 171720 46720
rect 171560 46720 171720 46880
rect 171560 46880 171720 47040
rect 171560 47040 171720 47200
rect 171560 47200 171720 47360
rect 171560 47360 171720 47520
rect 171560 47520 171720 47680
rect 171560 47680 171720 47840
rect 171560 47840 171720 48000
rect 171560 48000 171720 48160
rect 171560 48160 171720 48320
rect 171560 48320 171720 48480
rect 171560 48480 171720 48640
rect 171560 48640 171720 48800
rect 171560 48800 171720 48960
rect 171560 48960 171720 49120
rect 171560 49120 171720 49280
rect 171560 49280 171720 49440
rect 171560 49440 171720 49600
rect 171560 49600 171720 49760
rect 171560 49760 171720 49920
rect 171560 49920 171720 50080
rect 171560 50080 171720 50240
rect 171560 50240 171720 50400
rect 171560 50400 171720 50560
rect 171560 50560 171720 50720
rect 171560 50720 171720 50880
rect 171560 50880 171720 51040
rect 171560 51040 171720 51200
rect 171560 51200 171720 51360
rect 171560 51360 171720 51520
rect 171560 51520 171720 51680
rect 171560 51680 171720 51840
rect 171560 51840 171720 52000
rect 171560 52000 171720 52160
rect 171560 52160 171720 52320
rect 171560 52320 171720 52480
rect 171560 52480 171720 52640
rect 171560 52640 171720 52800
rect 171560 52800 171720 52960
rect 171560 52960 171720 53120
rect 171720 43040 171880 43200
rect 171720 43200 171880 43360
rect 171720 43360 171880 43520
rect 171720 43520 171880 43680
rect 171720 43680 171880 43840
rect 171720 43840 171880 44000
rect 171720 44000 171880 44160
rect 171720 44160 171880 44320
rect 171720 44320 171880 44480
rect 171720 44480 171880 44640
rect 171720 44640 171880 44800
rect 171720 44800 171880 44960
rect 171720 44960 171880 45120
rect 171720 45120 171880 45280
rect 171720 45280 171880 45440
rect 171720 45440 171880 45600
rect 171720 45600 171880 45760
rect 171720 45760 171880 45920
rect 171720 45920 171880 46080
rect 171720 46080 171880 46240
rect 171720 46240 171880 46400
rect 171720 46400 171880 46560
rect 171720 46560 171880 46720
rect 171720 46720 171880 46880
rect 171720 46880 171880 47040
rect 171720 47040 171880 47200
rect 171720 47200 171880 47360
rect 171720 47360 171880 47520
rect 171720 47520 171880 47680
rect 171720 47680 171880 47840
rect 171720 47840 171880 48000
rect 171720 48000 171880 48160
rect 171720 48160 171880 48320
rect 171720 48320 171880 48480
rect 171720 48480 171880 48640
rect 171720 48640 171880 48800
rect 171720 48800 171880 48960
rect 171720 48960 171880 49120
rect 171720 49120 171880 49280
rect 171720 49280 171880 49440
rect 171720 49440 171880 49600
rect 171720 49600 171880 49760
rect 171720 49760 171880 49920
rect 171720 49920 171880 50080
rect 171720 50080 171880 50240
rect 171720 50240 171880 50400
rect 171720 50400 171880 50560
rect 171720 50560 171880 50720
rect 171720 50720 171880 50880
rect 171720 50880 171880 51040
rect 171720 51040 171880 51200
rect 171720 51200 171880 51360
rect 171720 51360 171880 51520
rect 171720 51520 171880 51680
rect 171720 51680 171880 51840
rect 171720 51840 171880 52000
rect 171720 52000 171880 52160
rect 171720 52160 171880 52320
rect 171720 52320 171880 52480
rect 171720 52480 171880 52640
rect 171720 52640 171880 52800
rect 171720 52800 171880 52960
rect 171880 42400 172040 42560
rect 171880 42560 172040 42720
rect 171880 42720 172040 42880
rect 171880 42880 172040 43040
rect 171880 43040 172040 43200
rect 171880 43200 172040 43360
rect 171880 43360 172040 43520
rect 171880 43520 172040 43680
rect 171880 43680 172040 43840
rect 171880 43840 172040 44000
rect 171880 44000 172040 44160
rect 171880 44160 172040 44320
rect 171880 44320 172040 44480
rect 171880 44480 172040 44640
rect 171880 44640 172040 44800
rect 171880 44800 172040 44960
rect 171880 44960 172040 45120
rect 171880 45120 172040 45280
rect 171880 45280 172040 45440
rect 171880 45440 172040 45600
rect 171880 45600 172040 45760
rect 171880 45760 172040 45920
rect 171880 45920 172040 46080
rect 171880 46080 172040 46240
rect 171880 46240 172040 46400
rect 171880 46400 172040 46560
rect 171880 46560 172040 46720
rect 171880 46720 172040 46880
rect 171880 46880 172040 47040
rect 171880 47040 172040 47200
rect 171880 47200 172040 47360
rect 171880 47360 172040 47520
rect 171880 47520 172040 47680
rect 171880 47680 172040 47840
rect 171880 47840 172040 48000
rect 171880 48000 172040 48160
rect 171880 48160 172040 48320
rect 171880 48320 172040 48480
rect 171880 48480 172040 48640
rect 171880 48640 172040 48800
rect 171880 48800 172040 48960
rect 171880 48960 172040 49120
rect 171880 49120 172040 49280
rect 171880 49280 172040 49440
rect 171880 49440 172040 49600
rect 171880 49600 172040 49760
rect 171880 49760 172040 49920
rect 171880 49920 172040 50080
rect 171880 50080 172040 50240
rect 171880 50240 172040 50400
rect 171880 50400 172040 50560
rect 171880 50560 172040 50720
rect 171880 50720 172040 50880
rect 171880 50880 172040 51040
rect 171880 51040 172040 51200
rect 171880 51200 172040 51360
rect 171880 51360 172040 51520
rect 171880 51520 172040 51680
rect 171880 51680 172040 51840
rect 171880 51840 172040 52000
rect 171880 52000 172040 52160
rect 171880 52160 172040 52320
rect 171880 52320 172040 52480
rect 171880 52480 172040 52640
rect 171880 52640 172040 52800
rect 172040 41920 172200 42080
rect 172040 42080 172200 42240
rect 172040 42240 172200 42400
rect 172040 42400 172200 42560
rect 172040 42560 172200 42720
rect 172040 42720 172200 42880
rect 172040 42880 172200 43040
rect 172040 43040 172200 43200
rect 172040 43200 172200 43360
rect 172040 43360 172200 43520
rect 172040 43520 172200 43680
rect 172040 43680 172200 43840
rect 172040 43840 172200 44000
rect 172040 44000 172200 44160
rect 172040 44160 172200 44320
rect 172040 44320 172200 44480
rect 172040 44480 172200 44640
rect 172040 44640 172200 44800
rect 172040 44800 172200 44960
rect 172040 44960 172200 45120
rect 172040 45120 172200 45280
rect 172040 45280 172200 45440
rect 172040 45440 172200 45600
rect 172040 45600 172200 45760
rect 172040 45760 172200 45920
rect 172040 45920 172200 46080
rect 172040 46080 172200 46240
rect 172040 46240 172200 46400
rect 172040 46400 172200 46560
rect 172040 46560 172200 46720
rect 172040 46720 172200 46880
rect 172040 46880 172200 47040
rect 172040 47040 172200 47200
rect 172040 47200 172200 47360
rect 172040 47360 172200 47520
rect 172040 47520 172200 47680
rect 172040 47680 172200 47840
rect 172040 47840 172200 48000
rect 172040 48000 172200 48160
rect 172040 48160 172200 48320
rect 172040 48320 172200 48480
rect 172040 48480 172200 48640
rect 172040 48640 172200 48800
rect 172040 48800 172200 48960
rect 172040 48960 172200 49120
rect 172040 49120 172200 49280
rect 172040 49280 172200 49440
rect 172040 49440 172200 49600
rect 172040 49600 172200 49760
rect 172040 49760 172200 49920
rect 172040 49920 172200 50080
rect 172040 50080 172200 50240
rect 172040 50240 172200 50400
rect 172040 50400 172200 50560
rect 172040 50560 172200 50720
rect 172040 50720 172200 50880
rect 172040 50880 172200 51040
rect 172040 51040 172200 51200
rect 172040 51200 172200 51360
rect 172040 51360 172200 51520
rect 172040 51520 172200 51680
rect 172040 51680 172200 51840
rect 172040 51840 172200 52000
rect 172040 52000 172200 52160
rect 172040 52160 172200 52320
rect 172040 52320 172200 52480
rect 172040 52480 172200 52640
rect 172200 41440 172360 41600
rect 172200 41600 172360 41760
rect 172200 41760 172360 41920
rect 172200 41920 172360 42080
rect 172200 42080 172360 42240
rect 172200 42240 172360 42400
rect 172200 42400 172360 42560
rect 172200 42560 172360 42720
rect 172200 42720 172360 42880
rect 172200 42880 172360 43040
rect 172200 43040 172360 43200
rect 172200 43200 172360 43360
rect 172200 43360 172360 43520
rect 172200 43520 172360 43680
rect 172200 43680 172360 43840
rect 172200 43840 172360 44000
rect 172200 44000 172360 44160
rect 172200 44160 172360 44320
rect 172200 44320 172360 44480
rect 172200 44480 172360 44640
rect 172200 44640 172360 44800
rect 172200 44800 172360 44960
rect 172200 44960 172360 45120
rect 172200 45120 172360 45280
rect 172200 45280 172360 45440
rect 172200 45440 172360 45600
rect 172200 45600 172360 45760
rect 172200 45760 172360 45920
rect 172200 45920 172360 46080
rect 172200 46080 172360 46240
rect 172200 46240 172360 46400
rect 172200 46400 172360 46560
rect 172200 46560 172360 46720
rect 172200 46720 172360 46880
rect 172200 46880 172360 47040
rect 172200 47040 172360 47200
rect 172200 47200 172360 47360
rect 172200 47360 172360 47520
rect 172200 47520 172360 47680
rect 172200 47680 172360 47840
rect 172200 47840 172360 48000
rect 172200 48000 172360 48160
rect 172200 48160 172360 48320
rect 172200 48320 172360 48480
rect 172200 48480 172360 48640
rect 172200 48640 172360 48800
rect 172200 48800 172360 48960
rect 172200 48960 172360 49120
rect 172200 49120 172360 49280
rect 172200 49280 172360 49440
rect 172200 49440 172360 49600
rect 172200 49600 172360 49760
rect 172200 49760 172360 49920
rect 172200 49920 172360 50080
rect 172200 50080 172360 50240
rect 172200 50240 172360 50400
rect 172200 50400 172360 50560
rect 172200 50560 172360 50720
rect 172200 50720 172360 50880
rect 172200 50880 172360 51040
rect 172200 51040 172360 51200
rect 172200 51200 172360 51360
rect 172200 51360 172360 51520
rect 172200 51520 172360 51680
rect 172200 51680 172360 51840
rect 172200 51840 172360 52000
rect 172200 52000 172360 52160
rect 172200 52160 172360 52320
rect 172200 52320 172360 52480
rect 172360 40800 172520 40960
rect 172360 40960 172520 41120
rect 172360 41120 172520 41280
rect 172360 41280 172520 41440
rect 172360 41440 172520 41600
rect 172360 41600 172520 41760
rect 172360 41760 172520 41920
rect 172360 41920 172520 42080
rect 172360 42080 172520 42240
rect 172360 42240 172520 42400
rect 172360 42400 172520 42560
rect 172360 42560 172520 42720
rect 172360 42720 172520 42880
rect 172360 42880 172520 43040
rect 172360 43040 172520 43200
rect 172360 43200 172520 43360
rect 172360 43360 172520 43520
rect 172360 43520 172520 43680
rect 172360 43680 172520 43840
rect 172360 43840 172520 44000
rect 172360 44000 172520 44160
rect 172360 44160 172520 44320
rect 172360 44320 172520 44480
rect 172360 44480 172520 44640
rect 172360 44640 172520 44800
rect 172360 44800 172520 44960
rect 172360 44960 172520 45120
rect 172360 45120 172520 45280
rect 172360 45280 172520 45440
rect 172360 45440 172520 45600
rect 172360 45600 172520 45760
rect 172360 45760 172520 45920
rect 172360 45920 172520 46080
rect 172360 46080 172520 46240
rect 172360 46240 172520 46400
rect 172360 46400 172520 46560
rect 172360 46560 172520 46720
rect 172360 46720 172520 46880
rect 172360 46880 172520 47040
rect 172360 47040 172520 47200
rect 172360 47200 172520 47360
rect 172360 47360 172520 47520
rect 172360 47520 172520 47680
rect 172360 47680 172520 47840
rect 172360 47840 172520 48000
rect 172360 48000 172520 48160
rect 172360 48160 172520 48320
rect 172360 48320 172520 48480
rect 172360 48480 172520 48640
rect 172360 48640 172520 48800
rect 172360 48800 172520 48960
rect 172360 48960 172520 49120
rect 172360 49120 172520 49280
rect 172360 49280 172520 49440
rect 172360 49440 172520 49600
rect 172360 49600 172520 49760
rect 172360 49760 172520 49920
rect 172360 49920 172520 50080
rect 172360 50080 172520 50240
rect 172360 50240 172520 50400
rect 172360 50400 172520 50560
rect 172360 50560 172520 50720
rect 172360 50720 172520 50880
rect 172360 50880 172520 51040
rect 172360 51040 172520 51200
rect 172360 51200 172520 51360
rect 172360 51360 172520 51520
rect 172360 51520 172520 51680
rect 172360 51680 172520 51840
rect 172360 51840 172520 52000
rect 172360 52000 172520 52160
rect 172360 52160 172520 52320
rect 172520 40160 172680 40320
rect 172520 40320 172680 40480
rect 172520 40480 172680 40640
rect 172520 40640 172680 40800
rect 172520 40800 172680 40960
rect 172520 40960 172680 41120
rect 172520 41120 172680 41280
rect 172520 41280 172680 41440
rect 172520 41440 172680 41600
rect 172520 41600 172680 41760
rect 172520 41760 172680 41920
rect 172520 41920 172680 42080
rect 172520 42080 172680 42240
rect 172520 42240 172680 42400
rect 172520 42400 172680 42560
rect 172520 42560 172680 42720
rect 172520 42720 172680 42880
rect 172520 42880 172680 43040
rect 172520 43040 172680 43200
rect 172520 43200 172680 43360
rect 172520 43360 172680 43520
rect 172520 43520 172680 43680
rect 172520 43680 172680 43840
rect 172520 43840 172680 44000
rect 172520 44000 172680 44160
rect 172520 44160 172680 44320
rect 172520 44320 172680 44480
rect 172520 44480 172680 44640
rect 172520 44640 172680 44800
rect 172520 44800 172680 44960
rect 172520 44960 172680 45120
rect 172520 45120 172680 45280
rect 172520 45280 172680 45440
rect 172520 45440 172680 45600
rect 172520 45600 172680 45760
rect 172520 45760 172680 45920
rect 172520 45920 172680 46080
rect 172520 46080 172680 46240
rect 172520 46240 172680 46400
rect 172520 46400 172680 46560
rect 172520 46560 172680 46720
rect 172520 46720 172680 46880
rect 172520 46880 172680 47040
rect 172520 47040 172680 47200
rect 172520 47200 172680 47360
rect 172520 47360 172680 47520
rect 172520 47520 172680 47680
rect 172520 47680 172680 47840
rect 172520 47840 172680 48000
rect 172520 48000 172680 48160
rect 172520 48160 172680 48320
rect 172520 48320 172680 48480
rect 172520 48480 172680 48640
rect 172520 48640 172680 48800
rect 172520 48800 172680 48960
rect 172520 48960 172680 49120
rect 172520 49120 172680 49280
rect 172520 49280 172680 49440
rect 172520 49440 172680 49600
rect 172520 49600 172680 49760
rect 172520 49760 172680 49920
rect 172520 49920 172680 50080
rect 172520 50080 172680 50240
rect 172520 50240 172680 50400
rect 172520 50400 172680 50560
rect 172520 50560 172680 50720
rect 172520 50720 172680 50880
rect 172520 50880 172680 51040
rect 172520 51040 172680 51200
rect 172520 51200 172680 51360
rect 172520 51360 172680 51520
rect 172520 51520 172680 51680
rect 172520 51680 172680 51840
rect 172680 39680 172840 39840
rect 172680 39840 172840 40000
rect 172680 40000 172840 40160
rect 172680 40160 172840 40320
rect 172680 40320 172840 40480
rect 172680 40480 172840 40640
rect 172680 40640 172840 40800
rect 172680 40800 172840 40960
rect 172680 40960 172840 41120
rect 172680 41120 172840 41280
rect 172680 41280 172840 41440
rect 172680 41440 172840 41600
rect 172680 41600 172840 41760
rect 172680 41760 172840 41920
rect 172680 41920 172840 42080
rect 172680 42080 172840 42240
rect 172680 42240 172840 42400
rect 172680 42400 172840 42560
rect 172680 42560 172840 42720
rect 172680 42720 172840 42880
rect 172680 42880 172840 43040
rect 172680 43040 172840 43200
rect 172680 43200 172840 43360
rect 172680 43360 172840 43520
rect 172680 43520 172840 43680
rect 172680 43680 172840 43840
rect 172680 43840 172840 44000
rect 172680 44000 172840 44160
rect 172680 44160 172840 44320
rect 172680 44320 172840 44480
rect 172680 44480 172840 44640
rect 172680 44640 172840 44800
rect 172680 44800 172840 44960
rect 172680 44960 172840 45120
rect 172680 45120 172840 45280
rect 172680 45280 172840 45440
rect 172680 45440 172840 45600
rect 172680 45600 172840 45760
rect 172680 45760 172840 45920
rect 172680 45920 172840 46080
rect 172680 46080 172840 46240
rect 172680 46240 172840 46400
rect 172680 46400 172840 46560
rect 172680 46560 172840 46720
rect 172680 46720 172840 46880
rect 172680 46880 172840 47040
rect 172680 47040 172840 47200
rect 172680 47200 172840 47360
rect 172680 47360 172840 47520
rect 172680 47520 172840 47680
rect 172680 47680 172840 47840
rect 172680 47840 172840 48000
rect 172680 48000 172840 48160
rect 172680 48160 172840 48320
rect 172680 48320 172840 48480
rect 172680 48480 172840 48640
rect 172680 48640 172840 48800
rect 172680 48800 172840 48960
rect 172680 48960 172840 49120
rect 172680 49120 172840 49280
rect 172680 49280 172840 49440
rect 172680 49440 172840 49600
rect 172680 49600 172840 49760
rect 172680 49760 172840 49920
rect 172680 49920 172840 50080
rect 172680 50080 172840 50240
rect 172680 50240 172840 50400
rect 172680 50400 172840 50560
rect 172680 50560 172840 50720
rect 172680 50720 172840 50880
rect 172680 50880 172840 51040
rect 172680 51040 172840 51200
rect 172680 51200 172840 51360
rect 172680 51360 172840 51520
rect 172840 39040 173000 39200
rect 172840 39200 173000 39360
rect 172840 39360 173000 39520
rect 172840 39520 173000 39680
rect 172840 39680 173000 39840
rect 172840 39840 173000 40000
rect 172840 40000 173000 40160
rect 172840 40160 173000 40320
rect 172840 40320 173000 40480
rect 172840 40480 173000 40640
rect 172840 40640 173000 40800
rect 172840 40800 173000 40960
rect 172840 40960 173000 41120
rect 172840 41120 173000 41280
rect 172840 41280 173000 41440
rect 172840 41440 173000 41600
rect 172840 41600 173000 41760
rect 172840 41760 173000 41920
rect 172840 41920 173000 42080
rect 172840 42080 173000 42240
rect 172840 42240 173000 42400
rect 172840 42400 173000 42560
rect 172840 42560 173000 42720
rect 172840 42720 173000 42880
rect 172840 42880 173000 43040
rect 172840 43040 173000 43200
rect 172840 43200 173000 43360
rect 172840 43360 173000 43520
rect 172840 43520 173000 43680
rect 172840 43680 173000 43840
rect 172840 43840 173000 44000
rect 172840 44000 173000 44160
rect 172840 44160 173000 44320
rect 172840 44320 173000 44480
rect 172840 44480 173000 44640
rect 172840 44640 173000 44800
rect 172840 44800 173000 44960
rect 172840 44960 173000 45120
rect 172840 45120 173000 45280
rect 172840 45280 173000 45440
rect 172840 45440 173000 45600
rect 172840 45600 173000 45760
rect 172840 45760 173000 45920
rect 172840 45920 173000 46080
rect 172840 46080 173000 46240
rect 172840 46240 173000 46400
rect 172840 46400 173000 46560
rect 172840 46560 173000 46720
rect 172840 46720 173000 46880
rect 172840 46880 173000 47040
rect 172840 47040 173000 47200
rect 172840 47200 173000 47360
rect 172840 47360 173000 47520
rect 172840 47520 173000 47680
rect 172840 47680 173000 47840
rect 172840 47840 173000 48000
rect 172840 48000 173000 48160
rect 172840 48160 173000 48320
rect 172840 48320 173000 48480
rect 172840 48480 173000 48640
rect 172840 48640 173000 48800
rect 172840 48800 173000 48960
rect 172840 48960 173000 49120
rect 172840 49120 173000 49280
rect 172840 49280 173000 49440
rect 172840 49440 173000 49600
rect 172840 49600 173000 49760
rect 172840 49760 173000 49920
rect 172840 49920 173000 50080
rect 172840 50080 173000 50240
rect 172840 50240 173000 50400
rect 172840 50400 173000 50560
rect 172840 50560 173000 50720
rect 172840 50720 173000 50880
rect 172840 50880 173000 51040
rect 173000 38400 173160 38560
rect 173000 38560 173160 38720
rect 173000 38720 173160 38880
rect 173000 38880 173160 39040
rect 173000 39040 173160 39200
rect 173000 39200 173160 39360
rect 173000 39360 173160 39520
rect 173000 39520 173160 39680
rect 173000 39680 173160 39840
rect 173000 39840 173160 40000
rect 173000 40000 173160 40160
rect 173000 40160 173160 40320
rect 173000 40320 173160 40480
rect 173000 40480 173160 40640
rect 173000 40640 173160 40800
rect 173000 40800 173160 40960
rect 173000 40960 173160 41120
rect 173000 41120 173160 41280
rect 173000 41280 173160 41440
rect 173000 41440 173160 41600
rect 173000 41600 173160 41760
rect 173000 41760 173160 41920
rect 173000 41920 173160 42080
rect 173000 42080 173160 42240
rect 173000 42240 173160 42400
rect 173000 42400 173160 42560
rect 173000 42560 173160 42720
rect 173000 42720 173160 42880
rect 173000 42880 173160 43040
rect 173000 43040 173160 43200
rect 173000 43200 173160 43360
rect 173000 43360 173160 43520
rect 173000 43520 173160 43680
rect 173000 43680 173160 43840
rect 173000 43840 173160 44000
rect 173000 44000 173160 44160
rect 173000 44160 173160 44320
rect 173000 44320 173160 44480
rect 173000 44480 173160 44640
rect 173000 44640 173160 44800
rect 173000 44800 173160 44960
rect 173000 44960 173160 45120
rect 173000 45120 173160 45280
rect 173000 45280 173160 45440
rect 173000 45440 173160 45600
rect 173000 45600 173160 45760
rect 173000 45760 173160 45920
rect 173000 45920 173160 46080
rect 173000 46080 173160 46240
rect 173000 46240 173160 46400
rect 173000 46400 173160 46560
rect 173000 46560 173160 46720
rect 173000 46720 173160 46880
rect 173000 46880 173160 47040
rect 173000 47040 173160 47200
rect 173000 47200 173160 47360
rect 173000 47360 173160 47520
rect 173000 47520 173160 47680
rect 173000 47680 173160 47840
rect 173000 47840 173160 48000
rect 173000 48000 173160 48160
rect 173000 48160 173160 48320
rect 173000 48320 173160 48480
rect 173000 48480 173160 48640
rect 173000 48640 173160 48800
rect 173000 48800 173160 48960
rect 173000 48960 173160 49120
rect 173000 49120 173160 49280
rect 173000 49280 173160 49440
rect 173000 49440 173160 49600
rect 173000 49600 173160 49760
rect 173000 49760 173160 49920
rect 173000 49920 173160 50080
rect 173000 50080 173160 50240
rect 173000 50240 173160 50400
rect 173000 50400 173160 50560
rect 173160 37600 173320 37760
rect 173160 37760 173320 37920
rect 173160 37920 173320 38080
rect 173160 38080 173320 38240
rect 173160 38240 173320 38400
rect 173160 38400 173320 38560
rect 173160 38560 173320 38720
rect 173160 38720 173320 38880
rect 173160 38880 173320 39040
rect 173160 39040 173320 39200
rect 173160 39200 173320 39360
rect 173160 39360 173320 39520
rect 173160 39520 173320 39680
rect 173160 39680 173320 39840
rect 173160 39840 173320 40000
rect 173160 40000 173320 40160
rect 173160 40160 173320 40320
rect 173160 40320 173320 40480
rect 173160 40480 173320 40640
rect 173160 40640 173320 40800
rect 173160 40800 173320 40960
rect 173160 40960 173320 41120
rect 173160 41120 173320 41280
rect 173160 41280 173320 41440
rect 173160 41440 173320 41600
rect 173160 41600 173320 41760
rect 173160 41760 173320 41920
rect 173160 41920 173320 42080
rect 173160 42080 173320 42240
rect 173160 42240 173320 42400
rect 173160 42400 173320 42560
rect 173160 42560 173320 42720
rect 173160 42720 173320 42880
rect 173160 42880 173320 43040
rect 173160 43040 173320 43200
rect 173160 43200 173320 43360
rect 173160 43360 173320 43520
rect 173160 43520 173320 43680
rect 173160 43680 173320 43840
rect 173160 43840 173320 44000
rect 173160 44000 173320 44160
rect 173160 44160 173320 44320
rect 173160 44320 173320 44480
rect 173160 44480 173320 44640
rect 173160 44640 173320 44800
rect 173160 44800 173320 44960
rect 173160 44960 173320 45120
rect 173160 45120 173320 45280
rect 173160 45280 173320 45440
rect 173160 45440 173320 45600
rect 173160 45600 173320 45760
rect 173160 45760 173320 45920
rect 173160 45920 173320 46080
rect 173160 46080 173320 46240
rect 173160 46240 173320 46400
rect 173160 46400 173320 46560
rect 173160 46560 173320 46720
rect 173160 46720 173320 46880
rect 173160 46880 173320 47040
rect 173160 47040 173320 47200
rect 173160 47200 173320 47360
rect 173160 47360 173320 47520
rect 173160 47520 173320 47680
rect 173160 47680 173320 47840
rect 173160 47840 173320 48000
rect 173160 48000 173320 48160
rect 173160 48160 173320 48320
rect 173160 48320 173320 48480
rect 173160 48480 173320 48640
rect 173160 48640 173320 48800
rect 173160 48800 173320 48960
rect 173160 48960 173320 49120
rect 173160 49120 173320 49280
rect 173160 49280 173320 49440
rect 173160 49440 173320 49600
rect 173160 49600 173320 49760
rect 173160 49760 173320 49920
rect 173160 49920 173320 50080
rect 173320 36960 173480 37120
rect 173320 37120 173480 37280
rect 173320 37280 173480 37440
rect 173320 37440 173480 37600
rect 173320 37600 173480 37760
rect 173320 37760 173480 37920
rect 173320 37920 173480 38080
rect 173320 38080 173480 38240
rect 173320 38240 173480 38400
rect 173320 38400 173480 38560
rect 173320 38560 173480 38720
rect 173320 38720 173480 38880
rect 173320 38880 173480 39040
rect 173320 39040 173480 39200
rect 173320 39200 173480 39360
rect 173320 39360 173480 39520
rect 173320 39520 173480 39680
rect 173320 39680 173480 39840
rect 173320 39840 173480 40000
rect 173320 40000 173480 40160
rect 173320 40160 173480 40320
rect 173320 40320 173480 40480
rect 173320 40480 173480 40640
rect 173320 40640 173480 40800
rect 173320 40800 173480 40960
rect 173320 40960 173480 41120
rect 173320 41120 173480 41280
rect 173320 41280 173480 41440
rect 173320 41440 173480 41600
rect 173320 41600 173480 41760
rect 173320 41760 173480 41920
rect 173320 41920 173480 42080
rect 173320 42080 173480 42240
rect 173320 42240 173480 42400
rect 173320 42400 173480 42560
rect 173320 42560 173480 42720
rect 173320 42720 173480 42880
rect 173320 42880 173480 43040
rect 173320 43040 173480 43200
rect 173320 43200 173480 43360
rect 173320 43360 173480 43520
rect 173320 43520 173480 43680
rect 173320 43680 173480 43840
rect 173320 43840 173480 44000
rect 173320 44000 173480 44160
rect 173320 44160 173480 44320
rect 173320 44320 173480 44480
rect 173320 44480 173480 44640
rect 173320 44640 173480 44800
rect 173320 44800 173480 44960
rect 173320 44960 173480 45120
rect 173320 45120 173480 45280
rect 173320 45280 173480 45440
rect 173320 45440 173480 45600
rect 173320 45600 173480 45760
rect 173320 45760 173480 45920
rect 173320 45920 173480 46080
rect 173320 46080 173480 46240
rect 173320 46240 173480 46400
rect 173320 46400 173480 46560
rect 173320 46560 173480 46720
rect 173320 46720 173480 46880
rect 173320 46880 173480 47040
rect 173320 47040 173480 47200
rect 173320 47200 173480 47360
rect 173320 47360 173480 47520
rect 173320 47520 173480 47680
rect 173320 47680 173480 47840
rect 173320 47840 173480 48000
rect 173320 48000 173480 48160
rect 173320 48160 173480 48320
rect 173320 48320 173480 48480
rect 173320 48480 173480 48640
rect 173320 48640 173480 48800
rect 173320 48800 173480 48960
rect 173320 48960 173480 49120
rect 173320 49120 173480 49280
rect 173320 49280 173480 49440
rect 173320 49440 173480 49600
rect 173480 36160 173640 36320
rect 173480 36320 173640 36480
rect 173480 36480 173640 36640
rect 173480 36640 173640 36800
rect 173480 36800 173640 36960
rect 173480 36960 173640 37120
rect 173480 37120 173640 37280
rect 173480 37280 173640 37440
rect 173480 37440 173640 37600
rect 173480 37600 173640 37760
rect 173480 37760 173640 37920
rect 173480 37920 173640 38080
rect 173480 38080 173640 38240
rect 173480 38240 173640 38400
rect 173480 38400 173640 38560
rect 173480 38560 173640 38720
rect 173480 38720 173640 38880
rect 173480 38880 173640 39040
rect 173480 39040 173640 39200
rect 173480 39200 173640 39360
rect 173480 39360 173640 39520
rect 173480 39520 173640 39680
rect 173480 39680 173640 39840
rect 173480 39840 173640 40000
rect 173480 40000 173640 40160
rect 173480 40160 173640 40320
rect 173480 40320 173640 40480
rect 173480 40480 173640 40640
rect 173480 40640 173640 40800
rect 173480 40800 173640 40960
rect 173480 40960 173640 41120
rect 173480 41120 173640 41280
rect 173480 41280 173640 41440
rect 173480 41440 173640 41600
rect 173480 41600 173640 41760
rect 173480 41760 173640 41920
rect 173480 41920 173640 42080
rect 173480 42080 173640 42240
rect 173480 42240 173640 42400
rect 173480 42400 173640 42560
rect 173480 42560 173640 42720
rect 173480 42720 173640 42880
rect 173480 42880 173640 43040
rect 173480 43040 173640 43200
rect 173480 43200 173640 43360
rect 173480 43360 173640 43520
rect 173480 43520 173640 43680
rect 173480 43680 173640 43840
rect 173480 43840 173640 44000
rect 173480 44000 173640 44160
rect 173480 44160 173640 44320
rect 173480 44320 173640 44480
rect 173480 44480 173640 44640
rect 173480 44640 173640 44800
rect 173480 44800 173640 44960
rect 173480 44960 173640 45120
rect 173480 45120 173640 45280
rect 173480 45280 173640 45440
rect 173480 45440 173640 45600
rect 173480 45600 173640 45760
rect 173480 45760 173640 45920
rect 173480 45920 173640 46080
rect 173480 46080 173640 46240
rect 173480 46240 173640 46400
rect 173480 46400 173640 46560
rect 173480 46560 173640 46720
rect 173480 46720 173640 46880
rect 173480 46880 173640 47040
rect 173480 47040 173640 47200
rect 173480 47200 173640 47360
rect 173480 47360 173640 47520
rect 173480 47520 173640 47680
rect 173480 47680 173640 47840
rect 173480 47840 173640 48000
rect 173480 48000 173640 48160
rect 173480 48160 173640 48320
rect 173480 48320 173640 48480
rect 173480 48480 173640 48640
rect 173480 48640 173640 48800
rect 173480 48800 173640 48960
rect 173480 48960 173640 49120
rect 173640 35520 173800 35680
rect 173640 35680 173800 35840
rect 173640 35840 173800 36000
rect 173640 36000 173800 36160
rect 173640 36160 173800 36320
rect 173640 36320 173800 36480
rect 173640 36480 173800 36640
rect 173640 36640 173800 36800
rect 173640 36800 173800 36960
rect 173640 36960 173800 37120
rect 173640 37120 173800 37280
rect 173640 37280 173800 37440
rect 173640 37440 173800 37600
rect 173640 37600 173800 37760
rect 173640 37760 173800 37920
rect 173640 37920 173800 38080
rect 173640 38080 173800 38240
rect 173640 38240 173800 38400
rect 173640 38400 173800 38560
rect 173640 38560 173800 38720
rect 173640 38720 173800 38880
rect 173640 38880 173800 39040
rect 173640 39040 173800 39200
rect 173640 39200 173800 39360
rect 173640 39360 173800 39520
rect 173640 39520 173800 39680
rect 173640 39680 173800 39840
rect 173640 39840 173800 40000
rect 173640 40000 173800 40160
rect 173640 40160 173800 40320
rect 173640 40320 173800 40480
rect 173640 40480 173800 40640
rect 173640 40640 173800 40800
rect 173640 40800 173800 40960
rect 173640 40960 173800 41120
rect 173640 41120 173800 41280
rect 173640 41280 173800 41440
rect 173640 41440 173800 41600
rect 173640 41600 173800 41760
rect 173640 41760 173800 41920
rect 173640 41920 173800 42080
rect 173640 42080 173800 42240
rect 173640 42240 173800 42400
rect 173640 42400 173800 42560
rect 173640 42560 173800 42720
rect 173640 42720 173800 42880
rect 173640 42880 173800 43040
rect 173640 43040 173800 43200
rect 173640 43200 173800 43360
rect 173640 43360 173800 43520
rect 173640 43520 173800 43680
rect 173640 43680 173800 43840
rect 173640 43840 173800 44000
rect 173640 44000 173800 44160
rect 173640 44160 173800 44320
rect 173640 44320 173800 44480
rect 173640 44480 173800 44640
rect 173640 44640 173800 44800
rect 173640 44800 173800 44960
rect 173640 44960 173800 45120
rect 173640 45120 173800 45280
rect 173640 45280 173800 45440
rect 173640 45440 173800 45600
rect 173640 45600 173800 45760
rect 173640 45760 173800 45920
rect 173640 45920 173800 46080
rect 173640 46080 173800 46240
rect 173640 46240 173800 46400
rect 173640 46400 173800 46560
rect 173640 46560 173800 46720
rect 173640 46720 173800 46880
rect 173640 46880 173800 47040
rect 173640 47040 173800 47200
rect 173640 47200 173800 47360
rect 173640 47360 173800 47520
rect 173640 47520 173800 47680
rect 173640 47680 173800 47840
rect 173640 47840 173800 48000
rect 173640 48000 173800 48160
rect 173640 48160 173800 48320
rect 173640 48320 173800 48480
rect 173640 48480 173800 48640
rect 173800 34720 173960 34880
rect 173800 34880 173960 35040
rect 173800 35040 173960 35200
rect 173800 35200 173960 35360
rect 173800 35360 173960 35520
rect 173800 35520 173960 35680
rect 173800 35680 173960 35840
rect 173800 35840 173960 36000
rect 173800 36000 173960 36160
rect 173800 36160 173960 36320
rect 173800 36320 173960 36480
rect 173800 36480 173960 36640
rect 173800 36640 173960 36800
rect 173800 36800 173960 36960
rect 173800 36960 173960 37120
rect 173800 37120 173960 37280
rect 173800 37280 173960 37440
rect 173800 37440 173960 37600
rect 173800 37600 173960 37760
rect 173800 37760 173960 37920
rect 173800 37920 173960 38080
rect 173800 38080 173960 38240
rect 173800 38240 173960 38400
rect 173800 38400 173960 38560
rect 173800 38560 173960 38720
rect 173800 38720 173960 38880
rect 173800 38880 173960 39040
rect 173800 39040 173960 39200
rect 173800 39200 173960 39360
rect 173800 39360 173960 39520
rect 173800 39520 173960 39680
rect 173800 39680 173960 39840
rect 173800 39840 173960 40000
rect 173800 40000 173960 40160
rect 173800 40160 173960 40320
rect 173800 40320 173960 40480
rect 173800 40480 173960 40640
rect 173800 40640 173960 40800
rect 173800 40800 173960 40960
rect 173800 40960 173960 41120
rect 173800 41120 173960 41280
rect 173800 41280 173960 41440
rect 173800 41440 173960 41600
rect 173800 41600 173960 41760
rect 173800 41760 173960 41920
rect 173800 41920 173960 42080
rect 173800 42080 173960 42240
rect 173800 42240 173960 42400
rect 173800 42400 173960 42560
rect 173800 42560 173960 42720
rect 173800 42720 173960 42880
rect 173800 42880 173960 43040
rect 173800 43040 173960 43200
rect 173800 43200 173960 43360
rect 173800 43360 173960 43520
rect 173800 43520 173960 43680
rect 173800 43680 173960 43840
rect 173800 43840 173960 44000
rect 173800 44000 173960 44160
rect 173800 44160 173960 44320
rect 173800 44320 173960 44480
rect 173800 44480 173960 44640
rect 173800 44640 173960 44800
rect 173800 44800 173960 44960
rect 173800 44960 173960 45120
rect 173800 45120 173960 45280
rect 173800 45280 173960 45440
rect 173800 45440 173960 45600
rect 173800 45600 173960 45760
rect 173800 45760 173960 45920
rect 173800 45920 173960 46080
rect 173800 46080 173960 46240
rect 173800 46240 173960 46400
rect 173800 46400 173960 46560
rect 173800 46560 173960 46720
rect 173800 46720 173960 46880
rect 173800 46880 173960 47040
rect 173800 47040 173960 47200
rect 173800 47200 173960 47360
rect 173800 47360 173960 47520
rect 173800 47520 173960 47680
rect 173800 47680 173960 47840
rect 173800 47840 173960 48000
rect 173800 48000 173960 48160
rect 173960 34080 174120 34240
rect 173960 34240 174120 34400
rect 173960 34400 174120 34560
rect 173960 34560 174120 34720
rect 173960 34720 174120 34880
rect 173960 34880 174120 35040
rect 173960 35040 174120 35200
rect 173960 35200 174120 35360
rect 173960 35360 174120 35520
rect 173960 35520 174120 35680
rect 173960 35680 174120 35840
rect 173960 35840 174120 36000
rect 173960 36000 174120 36160
rect 173960 36160 174120 36320
rect 173960 36320 174120 36480
rect 173960 36480 174120 36640
rect 173960 36640 174120 36800
rect 173960 36800 174120 36960
rect 173960 36960 174120 37120
rect 173960 37120 174120 37280
rect 173960 37280 174120 37440
rect 173960 37440 174120 37600
rect 173960 37600 174120 37760
rect 173960 37760 174120 37920
rect 173960 37920 174120 38080
rect 173960 38080 174120 38240
rect 173960 38240 174120 38400
rect 173960 38400 174120 38560
rect 173960 38560 174120 38720
rect 173960 38720 174120 38880
rect 173960 38880 174120 39040
rect 173960 39040 174120 39200
rect 173960 39200 174120 39360
rect 173960 39360 174120 39520
rect 173960 39520 174120 39680
rect 173960 39680 174120 39840
rect 173960 39840 174120 40000
rect 173960 40000 174120 40160
rect 173960 40160 174120 40320
rect 173960 40320 174120 40480
rect 173960 40480 174120 40640
rect 173960 40640 174120 40800
rect 173960 40800 174120 40960
rect 173960 40960 174120 41120
rect 173960 41120 174120 41280
rect 173960 41280 174120 41440
rect 173960 41440 174120 41600
rect 173960 41600 174120 41760
rect 173960 41760 174120 41920
rect 173960 41920 174120 42080
rect 173960 42080 174120 42240
rect 173960 42240 174120 42400
rect 173960 42400 174120 42560
rect 173960 42560 174120 42720
rect 173960 42720 174120 42880
rect 173960 42880 174120 43040
rect 173960 43040 174120 43200
rect 173960 43200 174120 43360
rect 173960 43360 174120 43520
rect 173960 43520 174120 43680
rect 173960 43680 174120 43840
rect 173960 43840 174120 44000
rect 173960 44000 174120 44160
rect 173960 44160 174120 44320
rect 173960 44320 174120 44480
rect 173960 44480 174120 44640
rect 173960 44640 174120 44800
rect 173960 44800 174120 44960
rect 173960 44960 174120 45120
rect 173960 45120 174120 45280
rect 173960 45280 174120 45440
rect 173960 45440 174120 45600
rect 173960 45600 174120 45760
rect 173960 45760 174120 45920
rect 173960 45920 174120 46080
rect 173960 46080 174120 46240
rect 173960 46240 174120 46400
rect 173960 46400 174120 46560
rect 173960 46560 174120 46720
rect 173960 46720 174120 46880
rect 173960 46880 174120 47040
rect 173960 47040 174120 47200
rect 173960 47200 174120 47360
rect 173960 47360 174120 47520
rect 173960 47520 174120 47680
rect 174120 33280 174280 33440
rect 174120 33440 174280 33600
rect 174120 33600 174280 33760
rect 174120 33760 174280 33920
rect 174120 33920 174280 34080
rect 174120 34080 174280 34240
rect 174120 34240 174280 34400
rect 174120 34400 174280 34560
rect 174120 34560 174280 34720
rect 174120 34720 174280 34880
rect 174120 34880 174280 35040
rect 174120 35040 174280 35200
rect 174120 35200 174280 35360
rect 174120 35360 174280 35520
rect 174120 35520 174280 35680
rect 174120 35680 174280 35840
rect 174120 35840 174280 36000
rect 174120 36000 174280 36160
rect 174120 36160 174280 36320
rect 174120 36320 174280 36480
rect 174120 36480 174280 36640
rect 174120 36640 174280 36800
rect 174120 36800 174280 36960
rect 174120 36960 174280 37120
rect 174120 37120 174280 37280
rect 174120 37280 174280 37440
rect 174120 37440 174280 37600
rect 174120 37600 174280 37760
rect 174120 37760 174280 37920
rect 174120 37920 174280 38080
rect 174120 38080 174280 38240
rect 174120 38240 174280 38400
rect 174120 38400 174280 38560
rect 174120 38560 174280 38720
rect 174120 38720 174280 38880
rect 174120 38880 174280 39040
rect 174120 39040 174280 39200
rect 174120 39200 174280 39360
rect 174120 39360 174280 39520
rect 174120 39520 174280 39680
rect 174120 39680 174280 39840
rect 174120 39840 174280 40000
rect 174120 40000 174280 40160
rect 174120 40160 174280 40320
rect 174120 40320 174280 40480
rect 174120 40480 174280 40640
rect 174120 40640 174280 40800
rect 174120 40800 174280 40960
rect 174120 40960 174280 41120
rect 174120 41120 174280 41280
rect 174120 41280 174280 41440
rect 174120 41440 174280 41600
rect 174120 41600 174280 41760
rect 174120 41760 174280 41920
rect 174120 41920 174280 42080
rect 174120 42080 174280 42240
rect 174120 42240 174280 42400
rect 174120 42400 174280 42560
rect 174120 42560 174280 42720
rect 174120 42720 174280 42880
rect 174120 42880 174280 43040
rect 174120 43040 174280 43200
rect 174120 43200 174280 43360
rect 174120 43360 174280 43520
rect 174120 43520 174280 43680
rect 174120 43680 174280 43840
rect 174120 43840 174280 44000
rect 174120 44000 174280 44160
rect 174120 44160 174280 44320
rect 174120 44320 174280 44480
rect 174120 44480 174280 44640
rect 174120 44640 174280 44800
rect 174120 44800 174280 44960
rect 174120 44960 174280 45120
rect 174120 45120 174280 45280
rect 174120 45280 174280 45440
rect 174120 45440 174280 45600
rect 174120 45600 174280 45760
rect 174120 45760 174280 45920
rect 174120 45920 174280 46080
rect 174120 46080 174280 46240
rect 174120 46240 174280 46400
rect 174120 46400 174280 46560
rect 174120 46560 174280 46720
rect 174120 46720 174280 46880
rect 174120 46880 174280 47040
rect 174120 47040 174280 47200
rect 174280 32640 174440 32800
rect 174280 32800 174440 32960
rect 174280 32960 174440 33120
rect 174280 33120 174440 33280
rect 174280 33280 174440 33440
rect 174280 33440 174440 33600
rect 174280 33600 174440 33760
rect 174280 33760 174440 33920
rect 174280 33920 174440 34080
rect 174280 34080 174440 34240
rect 174280 34240 174440 34400
rect 174280 34400 174440 34560
rect 174280 34560 174440 34720
rect 174280 34720 174440 34880
rect 174280 34880 174440 35040
rect 174280 35040 174440 35200
rect 174280 35200 174440 35360
rect 174280 35360 174440 35520
rect 174280 35520 174440 35680
rect 174280 35680 174440 35840
rect 174280 35840 174440 36000
rect 174280 36000 174440 36160
rect 174280 36160 174440 36320
rect 174280 36320 174440 36480
rect 174280 36480 174440 36640
rect 174280 36640 174440 36800
rect 174280 36800 174440 36960
rect 174280 36960 174440 37120
rect 174280 37120 174440 37280
rect 174280 37280 174440 37440
rect 174280 37440 174440 37600
rect 174280 37600 174440 37760
rect 174280 37760 174440 37920
rect 174280 37920 174440 38080
rect 174280 38080 174440 38240
rect 174280 38240 174440 38400
rect 174280 38400 174440 38560
rect 174280 38560 174440 38720
rect 174280 38720 174440 38880
rect 174280 38880 174440 39040
rect 174280 39040 174440 39200
rect 174280 39200 174440 39360
rect 174280 39360 174440 39520
rect 174280 39520 174440 39680
rect 174280 39680 174440 39840
rect 174280 39840 174440 40000
rect 174280 40000 174440 40160
rect 174280 40160 174440 40320
rect 174280 40320 174440 40480
rect 174280 40480 174440 40640
rect 174280 40640 174440 40800
rect 174280 40800 174440 40960
rect 174280 40960 174440 41120
rect 174280 41120 174440 41280
rect 174280 41280 174440 41440
rect 174280 41440 174440 41600
rect 174280 41600 174440 41760
rect 174280 41760 174440 41920
rect 174280 41920 174440 42080
rect 174280 42080 174440 42240
rect 174280 42240 174440 42400
rect 174280 42400 174440 42560
rect 174280 42560 174440 42720
rect 174280 42720 174440 42880
rect 174280 42880 174440 43040
rect 174280 43040 174440 43200
rect 174280 43200 174440 43360
rect 174280 43360 174440 43520
rect 174280 43520 174440 43680
rect 174280 43680 174440 43840
rect 174280 43840 174440 44000
rect 174280 44000 174440 44160
rect 174280 44160 174440 44320
rect 174280 44320 174440 44480
rect 174280 44480 174440 44640
rect 174280 44640 174440 44800
rect 174280 44800 174440 44960
rect 174280 44960 174440 45120
rect 174280 45120 174440 45280
rect 174280 45280 174440 45440
rect 174280 45440 174440 45600
rect 174280 45600 174440 45760
rect 174280 45760 174440 45920
rect 174280 45920 174440 46080
rect 174280 46080 174440 46240
rect 174280 46240 174440 46400
rect 174280 46400 174440 46560
rect 174440 31840 174600 32000
rect 174440 32000 174600 32160
rect 174440 32160 174600 32320
rect 174440 32320 174600 32480
rect 174440 32480 174600 32640
rect 174440 32640 174600 32800
rect 174440 32800 174600 32960
rect 174440 32960 174600 33120
rect 174440 33120 174600 33280
rect 174440 33280 174600 33440
rect 174440 33440 174600 33600
rect 174440 33600 174600 33760
rect 174440 33760 174600 33920
rect 174440 33920 174600 34080
rect 174440 34080 174600 34240
rect 174440 34240 174600 34400
rect 174440 34400 174600 34560
rect 174440 34560 174600 34720
rect 174440 34720 174600 34880
rect 174440 34880 174600 35040
rect 174440 35040 174600 35200
rect 174440 35200 174600 35360
rect 174440 35360 174600 35520
rect 174440 35520 174600 35680
rect 174440 35680 174600 35840
rect 174440 35840 174600 36000
rect 174440 36000 174600 36160
rect 174440 36160 174600 36320
rect 174440 36320 174600 36480
rect 174440 36480 174600 36640
rect 174440 36640 174600 36800
rect 174440 36800 174600 36960
rect 174440 36960 174600 37120
rect 174440 37120 174600 37280
rect 174440 37280 174600 37440
rect 174440 37440 174600 37600
rect 174440 37600 174600 37760
rect 174440 37760 174600 37920
rect 174440 37920 174600 38080
rect 174440 38080 174600 38240
rect 174440 38240 174600 38400
rect 174440 38400 174600 38560
rect 174440 38560 174600 38720
rect 174440 38720 174600 38880
rect 174440 38880 174600 39040
rect 174440 39040 174600 39200
rect 174440 39200 174600 39360
rect 174440 39360 174600 39520
rect 174440 39520 174600 39680
rect 174440 39680 174600 39840
rect 174440 39840 174600 40000
rect 174440 40000 174600 40160
rect 174440 40160 174600 40320
rect 174440 40320 174600 40480
rect 174440 40480 174600 40640
rect 174440 40640 174600 40800
rect 174440 40800 174600 40960
rect 174440 40960 174600 41120
rect 174440 41120 174600 41280
rect 174440 41280 174600 41440
rect 174440 41440 174600 41600
rect 174440 41600 174600 41760
rect 174440 41760 174600 41920
rect 174440 41920 174600 42080
rect 174440 42080 174600 42240
rect 174440 42240 174600 42400
rect 174440 42400 174600 42560
rect 174440 42560 174600 42720
rect 174440 42720 174600 42880
rect 174440 42880 174600 43040
rect 174440 43040 174600 43200
rect 174440 43200 174600 43360
rect 174440 43360 174600 43520
rect 174440 43520 174600 43680
rect 174440 43680 174600 43840
rect 174440 43840 174600 44000
rect 174440 44000 174600 44160
rect 174440 44160 174600 44320
rect 174440 44320 174600 44480
rect 174440 44480 174600 44640
rect 174440 44640 174600 44800
rect 174440 44800 174600 44960
rect 174440 44960 174600 45120
rect 174440 45120 174600 45280
rect 174440 45280 174600 45440
rect 174440 45440 174600 45600
rect 174440 45600 174600 45760
rect 174440 45760 174600 45920
rect 174440 45920 174600 46080
rect 174600 31200 174760 31360
rect 174600 31360 174760 31520
rect 174600 31520 174760 31680
rect 174600 31680 174760 31840
rect 174600 31840 174760 32000
rect 174600 32000 174760 32160
rect 174600 32160 174760 32320
rect 174600 32320 174760 32480
rect 174600 32480 174760 32640
rect 174600 32640 174760 32800
rect 174600 32800 174760 32960
rect 174600 32960 174760 33120
rect 174600 33120 174760 33280
rect 174600 33280 174760 33440
rect 174600 33440 174760 33600
rect 174600 33600 174760 33760
rect 174600 33760 174760 33920
rect 174600 33920 174760 34080
rect 174600 34080 174760 34240
rect 174600 34240 174760 34400
rect 174600 34400 174760 34560
rect 174600 34560 174760 34720
rect 174600 34720 174760 34880
rect 174600 34880 174760 35040
rect 174600 35040 174760 35200
rect 174600 35200 174760 35360
rect 174600 35360 174760 35520
rect 174600 35520 174760 35680
rect 174600 35680 174760 35840
rect 174600 35840 174760 36000
rect 174600 36000 174760 36160
rect 174600 36160 174760 36320
rect 174600 36320 174760 36480
rect 174600 36480 174760 36640
rect 174600 36640 174760 36800
rect 174600 36800 174760 36960
rect 174600 36960 174760 37120
rect 174600 37120 174760 37280
rect 174600 37280 174760 37440
rect 174600 37440 174760 37600
rect 174600 37600 174760 37760
rect 174600 37760 174760 37920
rect 174600 37920 174760 38080
rect 174600 38080 174760 38240
rect 174600 38240 174760 38400
rect 174600 38400 174760 38560
rect 174600 38560 174760 38720
rect 174600 38720 174760 38880
rect 174600 38880 174760 39040
rect 174600 39040 174760 39200
rect 174600 39200 174760 39360
rect 174600 39360 174760 39520
rect 174600 39520 174760 39680
rect 174600 39680 174760 39840
rect 174600 39840 174760 40000
rect 174600 40000 174760 40160
rect 174600 40160 174760 40320
rect 174600 40320 174760 40480
rect 174600 40480 174760 40640
rect 174600 40640 174760 40800
rect 174600 40800 174760 40960
rect 174600 40960 174760 41120
rect 174600 41120 174760 41280
rect 174600 41280 174760 41440
rect 174600 41440 174760 41600
rect 174600 41600 174760 41760
rect 174600 41760 174760 41920
rect 174600 41920 174760 42080
rect 174600 42080 174760 42240
rect 174600 42240 174760 42400
rect 174600 42400 174760 42560
rect 174600 42560 174760 42720
rect 174600 42720 174760 42880
rect 174600 42880 174760 43040
rect 174600 43040 174760 43200
rect 174600 43200 174760 43360
rect 174600 43360 174760 43520
rect 174600 43520 174760 43680
rect 174600 43680 174760 43840
rect 174600 43840 174760 44000
rect 174600 44000 174760 44160
rect 174600 44160 174760 44320
rect 174600 44320 174760 44480
rect 174600 44480 174760 44640
rect 174600 44640 174760 44800
rect 174600 44800 174760 44960
rect 174600 44960 174760 45120
rect 174600 45120 174760 45280
rect 174600 45280 174760 45440
rect 174760 30560 174920 30720
rect 174760 30720 174920 30880
rect 174760 30880 174920 31040
rect 174760 31040 174920 31200
rect 174760 31200 174920 31360
rect 174760 31360 174920 31520
rect 174760 31520 174920 31680
rect 174760 31680 174920 31840
rect 174760 31840 174920 32000
rect 174760 32000 174920 32160
rect 174760 32160 174920 32320
rect 174760 32320 174920 32480
rect 174760 32480 174920 32640
rect 174760 32640 174920 32800
rect 174760 32800 174920 32960
rect 174760 32960 174920 33120
rect 174760 33120 174920 33280
rect 174760 33280 174920 33440
rect 174760 33440 174920 33600
rect 174760 33600 174920 33760
rect 174760 33760 174920 33920
rect 174760 33920 174920 34080
rect 174760 34080 174920 34240
rect 174760 34240 174920 34400
rect 174760 34400 174920 34560
rect 174760 34560 174920 34720
rect 174760 34720 174920 34880
rect 174760 34880 174920 35040
rect 174760 35040 174920 35200
rect 174760 35200 174920 35360
rect 174760 35360 174920 35520
rect 174760 35520 174920 35680
rect 174760 35680 174920 35840
rect 174760 35840 174920 36000
rect 174760 36000 174920 36160
rect 174760 36160 174920 36320
rect 174760 36320 174920 36480
rect 174760 36480 174920 36640
rect 174760 36640 174920 36800
rect 174760 36800 174920 36960
rect 174760 36960 174920 37120
rect 174760 37120 174920 37280
rect 174760 37280 174920 37440
rect 174760 37440 174920 37600
rect 174760 37600 174920 37760
rect 174760 37760 174920 37920
rect 174760 37920 174920 38080
rect 174760 38080 174920 38240
rect 174760 38240 174920 38400
rect 174760 38400 174920 38560
rect 174760 38560 174920 38720
rect 174760 38720 174920 38880
rect 174760 38880 174920 39040
rect 174760 39040 174920 39200
rect 174760 39200 174920 39360
rect 174760 39360 174920 39520
rect 174760 39520 174920 39680
rect 174760 39680 174920 39840
rect 174760 39840 174920 40000
rect 174760 40000 174920 40160
rect 174760 40160 174920 40320
rect 174760 40320 174920 40480
rect 174760 40480 174920 40640
rect 174760 40640 174920 40800
rect 174760 40800 174920 40960
rect 174760 40960 174920 41120
rect 174760 41120 174920 41280
rect 174760 41280 174920 41440
rect 174760 41440 174920 41600
rect 174760 41600 174920 41760
rect 174760 41760 174920 41920
rect 174760 41920 174920 42080
rect 174760 42080 174920 42240
rect 174760 42240 174920 42400
rect 174760 42400 174920 42560
rect 174760 42560 174920 42720
rect 174760 42720 174920 42880
rect 174760 42880 174920 43040
rect 174760 43040 174920 43200
rect 174760 43200 174920 43360
rect 174760 43360 174920 43520
rect 174760 43520 174920 43680
rect 174760 43680 174920 43840
rect 174760 43840 174920 44000
rect 174760 44000 174920 44160
rect 174760 44160 174920 44320
rect 174760 44320 174920 44480
rect 174760 44480 174920 44640
rect 174760 44640 174920 44800
rect 174760 44800 174920 44960
rect 174920 29760 175080 29920
rect 174920 29920 175080 30080
rect 174920 30080 175080 30240
rect 174920 30240 175080 30400
rect 174920 30400 175080 30560
rect 174920 30560 175080 30720
rect 174920 30720 175080 30880
rect 174920 30880 175080 31040
rect 174920 31040 175080 31200
rect 174920 31200 175080 31360
rect 174920 31360 175080 31520
rect 174920 31520 175080 31680
rect 174920 31680 175080 31840
rect 174920 31840 175080 32000
rect 174920 32000 175080 32160
rect 174920 32160 175080 32320
rect 174920 32320 175080 32480
rect 174920 32480 175080 32640
rect 174920 32640 175080 32800
rect 174920 32800 175080 32960
rect 174920 32960 175080 33120
rect 174920 33120 175080 33280
rect 174920 33280 175080 33440
rect 174920 33440 175080 33600
rect 174920 33600 175080 33760
rect 174920 33760 175080 33920
rect 174920 33920 175080 34080
rect 174920 34080 175080 34240
rect 174920 34240 175080 34400
rect 174920 34400 175080 34560
rect 174920 34560 175080 34720
rect 174920 34720 175080 34880
rect 174920 34880 175080 35040
rect 174920 35040 175080 35200
rect 174920 35200 175080 35360
rect 174920 35360 175080 35520
rect 174920 35520 175080 35680
rect 174920 35680 175080 35840
rect 174920 35840 175080 36000
rect 174920 36000 175080 36160
rect 174920 36160 175080 36320
rect 174920 36320 175080 36480
rect 174920 36480 175080 36640
rect 174920 36640 175080 36800
rect 174920 36800 175080 36960
rect 174920 36960 175080 37120
rect 174920 37120 175080 37280
rect 174920 37280 175080 37440
rect 174920 37440 175080 37600
rect 174920 37600 175080 37760
rect 174920 37760 175080 37920
rect 174920 37920 175080 38080
rect 174920 38080 175080 38240
rect 174920 38240 175080 38400
rect 174920 38400 175080 38560
rect 174920 38560 175080 38720
rect 174920 38720 175080 38880
rect 174920 38880 175080 39040
rect 174920 39040 175080 39200
rect 174920 39200 175080 39360
rect 174920 39360 175080 39520
rect 174920 39520 175080 39680
rect 174920 39680 175080 39840
rect 174920 39840 175080 40000
rect 174920 40000 175080 40160
rect 174920 40160 175080 40320
rect 174920 40320 175080 40480
rect 174920 40480 175080 40640
rect 174920 40640 175080 40800
rect 174920 40800 175080 40960
rect 174920 40960 175080 41120
rect 174920 41120 175080 41280
rect 174920 41280 175080 41440
rect 174920 41440 175080 41600
rect 174920 41600 175080 41760
rect 174920 41760 175080 41920
rect 174920 41920 175080 42080
rect 174920 42080 175080 42240
rect 174920 42240 175080 42400
rect 174920 42400 175080 42560
rect 174920 42560 175080 42720
rect 174920 42720 175080 42880
rect 174920 42880 175080 43040
rect 174920 43040 175080 43200
rect 174920 43200 175080 43360
rect 174920 43360 175080 43520
rect 174920 43520 175080 43680
rect 174920 43680 175080 43840
rect 174920 43840 175080 44000
rect 174920 44000 175080 44160
rect 174920 44160 175080 44320
rect 175080 29120 175240 29280
rect 175080 29280 175240 29440
rect 175080 29440 175240 29600
rect 175080 29600 175240 29760
rect 175080 29760 175240 29920
rect 175080 29920 175240 30080
rect 175080 30080 175240 30240
rect 175080 30240 175240 30400
rect 175080 30400 175240 30560
rect 175080 30560 175240 30720
rect 175080 30720 175240 30880
rect 175080 30880 175240 31040
rect 175080 31040 175240 31200
rect 175080 31200 175240 31360
rect 175080 31360 175240 31520
rect 175080 31520 175240 31680
rect 175080 31680 175240 31840
rect 175080 31840 175240 32000
rect 175080 32000 175240 32160
rect 175080 32160 175240 32320
rect 175080 32320 175240 32480
rect 175080 32480 175240 32640
rect 175080 32640 175240 32800
rect 175080 32800 175240 32960
rect 175080 32960 175240 33120
rect 175080 33120 175240 33280
rect 175080 33280 175240 33440
rect 175080 33440 175240 33600
rect 175080 33600 175240 33760
rect 175080 33760 175240 33920
rect 175080 33920 175240 34080
rect 175080 34080 175240 34240
rect 175080 34240 175240 34400
rect 175080 34400 175240 34560
rect 175080 34560 175240 34720
rect 175080 34720 175240 34880
rect 175080 34880 175240 35040
rect 175080 35040 175240 35200
rect 175080 35200 175240 35360
rect 175080 35360 175240 35520
rect 175080 35520 175240 35680
rect 175080 35680 175240 35840
rect 175080 35840 175240 36000
rect 175080 36000 175240 36160
rect 175080 36160 175240 36320
rect 175080 36320 175240 36480
rect 175080 36480 175240 36640
rect 175080 36640 175240 36800
rect 175080 36800 175240 36960
rect 175080 36960 175240 37120
rect 175080 37120 175240 37280
rect 175080 37280 175240 37440
rect 175080 37440 175240 37600
rect 175080 37600 175240 37760
rect 175080 37760 175240 37920
rect 175080 37920 175240 38080
rect 175080 38080 175240 38240
rect 175080 38240 175240 38400
rect 175080 38400 175240 38560
rect 175080 38560 175240 38720
rect 175080 38720 175240 38880
rect 175080 38880 175240 39040
rect 175080 39040 175240 39200
rect 175080 39200 175240 39360
rect 175080 39360 175240 39520
rect 175080 39520 175240 39680
rect 175080 39680 175240 39840
rect 175080 39840 175240 40000
rect 175080 40000 175240 40160
rect 175080 40160 175240 40320
rect 175080 40320 175240 40480
rect 175080 40480 175240 40640
rect 175080 40640 175240 40800
rect 175080 40800 175240 40960
rect 175080 40960 175240 41120
rect 175080 41120 175240 41280
rect 175080 41280 175240 41440
rect 175080 41440 175240 41600
rect 175080 41600 175240 41760
rect 175080 41760 175240 41920
rect 175080 41920 175240 42080
rect 175080 42080 175240 42240
rect 175080 42240 175240 42400
rect 175080 42400 175240 42560
rect 175080 42560 175240 42720
rect 175080 42720 175240 42880
rect 175080 42880 175240 43040
rect 175080 43040 175240 43200
rect 175080 43200 175240 43360
rect 175080 43360 175240 43520
rect 175080 43520 175240 43680
rect 175240 28160 175400 28320
rect 175240 28320 175400 28480
rect 175240 28480 175400 28640
rect 175240 28640 175400 28800
rect 175240 28800 175400 28960
rect 175240 28960 175400 29120
rect 175240 29120 175400 29280
rect 175240 29280 175400 29440
rect 175240 29440 175400 29600
rect 175240 29600 175400 29760
rect 175240 29760 175400 29920
rect 175240 29920 175400 30080
rect 175240 30080 175400 30240
rect 175240 30240 175400 30400
rect 175240 30400 175400 30560
rect 175240 30560 175400 30720
rect 175240 30720 175400 30880
rect 175240 30880 175400 31040
rect 175240 31040 175400 31200
rect 175240 31200 175400 31360
rect 175240 31360 175400 31520
rect 175240 31520 175400 31680
rect 175240 31680 175400 31840
rect 175240 31840 175400 32000
rect 175240 32000 175400 32160
rect 175240 32160 175400 32320
rect 175240 32320 175400 32480
rect 175240 32480 175400 32640
rect 175240 32640 175400 32800
rect 175240 32800 175400 32960
rect 175240 32960 175400 33120
rect 175240 33120 175400 33280
rect 175240 33280 175400 33440
rect 175240 33440 175400 33600
rect 175240 33600 175400 33760
rect 175240 33760 175400 33920
rect 175240 33920 175400 34080
rect 175240 34080 175400 34240
rect 175240 34240 175400 34400
rect 175240 34400 175400 34560
rect 175240 34560 175400 34720
rect 175240 34720 175400 34880
rect 175240 34880 175400 35040
rect 175240 35040 175400 35200
rect 175240 35200 175400 35360
rect 175240 35360 175400 35520
rect 175240 35520 175400 35680
rect 175240 35680 175400 35840
rect 175240 35840 175400 36000
rect 175240 36000 175400 36160
rect 175240 36160 175400 36320
rect 175240 36320 175400 36480
rect 175240 36480 175400 36640
rect 175240 36640 175400 36800
rect 175240 36800 175400 36960
rect 175240 36960 175400 37120
rect 175240 37120 175400 37280
rect 175240 37280 175400 37440
rect 175240 37440 175400 37600
rect 175240 37600 175400 37760
rect 175240 37760 175400 37920
rect 175240 37920 175400 38080
rect 175240 38080 175400 38240
rect 175240 38240 175400 38400
rect 175240 38400 175400 38560
rect 175240 38560 175400 38720
rect 175240 38720 175400 38880
rect 175240 38880 175400 39040
rect 175240 39040 175400 39200
rect 175240 39200 175400 39360
rect 175240 39360 175400 39520
rect 175240 39520 175400 39680
rect 175240 39680 175400 39840
rect 175240 39840 175400 40000
rect 175240 40000 175400 40160
rect 175240 40160 175400 40320
rect 175240 40320 175400 40480
rect 175240 40480 175400 40640
rect 175240 40640 175400 40800
rect 175240 40800 175400 40960
rect 175240 40960 175400 41120
rect 175240 41120 175400 41280
rect 175240 41280 175400 41440
rect 175240 41440 175400 41600
rect 175240 41600 175400 41760
rect 175240 41760 175400 41920
rect 175240 41920 175400 42080
rect 175240 42080 175400 42240
rect 175240 42240 175400 42400
rect 175240 42400 175400 42560
rect 175240 42560 175400 42720
rect 175240 42720 175400 42880
rect 175240 42880 175400 43040
rect 175400 27680 175560 27840
rect 175400 27840 175560 28000
rect 175400 28000 175560 28160
rect 175400 28160 175560 28320
rect 175400 28320 175560 28480
rect 175400 28480 175560 28640
rect 175400 28640 175560 28800
rect 175400 28800 175560 28960
rect 175400 28960 175560 29120
rect 175400 29120 175560 29280
rect 175400 29280 175560 29440
rect 175400 29440 175560 29600
rect 175400 29600 175560 29760
rect 175400 29760 175560 29920
rect 175400 29920 175560 30080
rect 175400 30080 175560 30240
rect 175400 30240 175560 30400
rect 175400 30400 175560 30560
rect 175400 30560 175560 30720
rect 175400 30720 175560 30880
rect 175400 30880 175560 31040
rect 175400 31040 175560 31200
rect 175400 31200 175560 31360
rect 175400 31360 175560 31520
rect 175400 31520 175560 31680
rect 175400 31680 175560 31840
rect 175400 31840 175560 32000
rect 175400 32000 175560 32160
rect 175400 32160 175560 32320
rect 175400 32320 175560 32480
rect 175400 32480 175560 32640
rect 175400 32640 175560 32800
rect 175400 32800 175560 32960
rect 175400 32960 175560 33120
rect 175400 33120 175560 33280
rect 175400 33280 175560 33440
rect 175400 33440 175560 33600
rect 175400 33600 175560 33760
rect 175400 33760 175560 33920
rect 175400 33920 175560 34080
rect 175400 34080 175560 34240
rect 175400 34240 175560 34400
rect 175400 34400 175560 34560
rect 175400 34560 175560 34720
rect 175400 34720 175560 34880
rect 175400 34880 175560 35040
rect 175400 35040 175560 35200
rect 175400 35200 175560 35360
rect 175400 35360 175560 35520
rect 175400 35520 175560 35680
rect 175400 35680 175560 35840
rect 175400 35840 175560 36000
rect 175400 36000 175560 36160
rect 175400 36160 175560 36320
rect 175400 36320 175560 36480
rect 175400 36480 175560 36640
rect 175400 36640 175560 36800
rect 175400 36800 175560 36960
rect 175400 36960 175560 37120
rect 175400 37120 175560 37280
rect 175400 37280 175560 37440
rect 175400 37440 175560 37600
rect 175400 37600 175560 37760
rect 175400 37760 175560 37920
rect 175400 37920 175560 38080
rect 175400 38080 175560 38240
rect 175400 38240 175560 38400
rect 175400 38400 175560 38560
rect 175400 38560 175560 38720
rect 175400 38720 175560 38880
rect 175400 38880 175560 39040
rect 175400 39040 175560 39200
rect 175400 39200 175560 39360
rect 175400 39360 175560 39520
rect 175400 39520 175560 39680
rect 175400 39680 175560 39840
rect 175400 39840 175560 40000
rect 175400 40000 175560 40160
rect 175400 40160 175560 40320
rect 175400 40320 175560 40480
rect 175400 40480 175560 40640
rect 175400 40640 175560 40800
rect 175400 40800 175560 40960
rect 175400 40960 175560 41120
rect 175400 41120 175560 41280
rect 175400 41280 175560 41440
rect 175400 41440 175560 41600
rect 175400 41600 175560 41760
rect 175400 41760 175560 41920
rect 175400 41920 175560 42080
rect 175400 42080 175560 42240
rect 175400 42240 175560 42400
rect 175560 27520 175720 27680
rect 175560 27680 175720 27840
rect 175560 27840 175720 28000
rect 175560 28000 175720 28160
rect 175560 28160 175720 28320
rect 175560 28320 175720 28480
rect 175560 28480 175720 28640
rect 175560 28640 175720 28800
rect 175560 28800 175720 28960
rect 175560 28960 175720 29120
rect 175560 29120 175720 29280
rect 175560 29280 175720 29440
rect 175560 29440 175720 29600
rect 175560 29600 175720 29760
rect 175560 29760 175720 29920
rect 175560 29920 175720 30080
rect 175560 30080 175720 30240
rect 175560 30240 175720 30400
rect 175560 30400 175720 30560
rect 175560 30560 175720 30720
rect 175560 30720 175720 30880
rect 175560 30880 175720 31040
rect 175560 31040 175720 31200
rect 175560 31200 175720 31360
rect 175560 31360 175720 31520
rect 175560 31520 175720 31680
rect 175560 31680 175720 31840
rect 175560 31840 175720 32000
rect 175560 32000 175720 32160
rect 175560 32160 175720 32320
rect 175560 32320 175720 32480
rect 175560 32480 175720 32640
rect 175560 32640 175720 32800
rect 175560 32800 175720 32960
rect 175560 32960 175720 33120
rect 175560 33120 175720 33280
rect 175560 33280 175720 33440
rect 175560 33440 175720 33600
rect 175560 33600 175720 33760
rect 175560 33760 175720 33920
rect 175560 33920 175720 34080
rect 175560 34080 175720 34240
rect 175560 34240 175720 34400
rect 175560 34400 175720 34560
rect 175560 34560 175720 34720
rect 175560 34720 175720 34880
rect 175560 34880 175720 35040
rect 175560 35040 175720 35200
rect 175560 35200 175720 35360
rect 175560 35360 175720 35520
rect 175560 35520 175720 35680
rect 175560 35680 175720 35840
rect 175560 35840 175720 36000
rect 175560 36000 175720 36160
rect 175560 36160 175720 36320
rect 175560 36320 175720 36480
rect 175560 36480 175720 36640
rect 175560 36640 175720 36800
rect 175560 36800 175720 36960
rect 175560 36960 175720 37120
rect 175560 37120 175720 37280
rect 175560 37280 175720 37440
rect 175560 37440 175720 37600
rect 175560 37600 175720 37760
rect 175560 37760 175720 37920
rect 175560 37920 175720 38080
rect 175560 38080 175720 38240
rect 175560 38240 175720 38400
rect 175560 38400 175720 38560
rect 175560 38560 175720 38720
rect 175560 38720 175720 38880
rect 175560 38880 175720 39040
rect 175560 39040 175720 39200
rect 175560 39200 175720 39360
rect 175560 39360 175720 39520
rect 175560 39520 175720 39680
rect 175560 39680 175720 39840
rect 175560 39840 175720 40000
rect 175560 40000 175720 40160
rect 175560 40160 175720 40320
rect 175560 40320 175720 40480
rect 175560 40480 175720 40640
rect 175560 40640 175720 40800
rect 175560 40800 175720 40960
rect 175560 40960 175720 41120
rect 175560 41120 175720 41280
rect 175560 41280 175720 41440
rect 175560 41440 175720 41600
rect 175720 27200 175880 27360
rect 175720 27360 175880 27520
rect 175720 27520 175880 27680
rect 175720 27680 175880 27840
rect 175720 27840 175880 28000
rect 175720 28000 175880 28160
rect 175720 28160 175880 28320
rect 175720 28320 175880 28480
rect 175720 28480 175880 28640
rect 175720 28640 175880 28800
rect 175720 28800 175880 28960
rect 175720 28960 175880 29120
rect 175720 29120 175880 29280
rect 175720 29280 175880 29440
rect 175720 29440 175880 29600
rect 175720 29600 175880 29760
rect 175720 29760 175880 29920
rect 175720 29920 175880 30080
rect 175720 30080 175880 30240
rect 175720 30240 175880 30400
rect 175720 30400 175880 30560
rect 175720 30560 175880 30720
rect 175720 30720 175880 30880
rect 175720 30880 175880 31040
rect 175720 31040 175880 31200
rect 175720 31200 175880 31360
rect 175720 31360 175880 31520
rect 175720 31520 175880 31680
rect 175720 31680 175880 31840
rect 175720 31840 175880 32000
rect 175720 32000 175880 32160
rect 175720 32160 175880 32320
rect 175720 32320 175880 32480
rect 175720 32480 175880 32640
rect 175720 32640 175880 32800
rect 175720 32800 175880 32960
rect 175720 32960 175880 33120
rect 175720 33120 175880 33280
rect 175720 33280 175880 33440
rect 175720 33440 175880 33600
rect 175720 33600 175880 33760
rect 175720 33760 175880 33920
rect 175720 33920 175880 34080
rect 175720 34080 175880 34240
rect 175720 34240 175880 34400
rect 175720 34400 175880 34560
rect 175720 34560 175880 34720
rect 175720 34720 175880 34880
rect 175720 34880 175880 35040
rect 175720 35040 175880 35200
rect 175720 35200 175880 35360
rect 175720 35360 175880 35520
rect 175720 35520 175880 35680
rect 175720 35680 175880 35840
rect 175720 35840 175880 36000
rect 175720 36000 175880 36160
rect 175720 36160 175880 36320
rect 175720 36320 175880 36480
rect 175720 36480 175880 36640
rect 175720 36640 175880 36800
rect 175720 36800 175880 36960
rect 175720 36960 175880 37120
rect 175720 37120 175880 37280
rect 175720 37280 175880 37440
rect 175720 37440 175880 37600
rect 175720 37600 175880 37760
rect 175720 37760 175880 37920
rect 175720 37920 175880 38080
rect 175720 38080 175880 38240
rect 175720 38240 175880 38400
rect 175720 38400 175880 38560
rect 175720 38560 175880 38720
rect 175720 38720 175880 38880
rect 175720 38880 175880 39040
rect 175720 39040 175880 39200
rect 175720 39200 175880 39360
rect 175720 39360 175880 39520
rect 175720 39520 175880 39680
rect 175720 39680 175880 39840
rect 175720 39840 175880 40000
rect 175720 40000 175880 40160
rect 175720 40160 175880 40320
rect 175720 40320 175880 40480
rect 175720 40480 175880 40640
rect 175720 40640 175880 40800
rect 175720 40800 175880 40960
rect 175880 27200 176040 27360
rect 175880 27360 176040 27520
rect 175880 27520 176040 27680
rect 175880 27680 176040 27840
rect 175880 27840 176040 28000
rect 175880 28000 176040 28160
rect 175880 28160 176040 28320
rect 175880 28320 176040 28480
rect 175880 28480 176040 28640
rect 175880 28640 176040 28800
rect 175880 28800 176040 28960
rect 175880 28960 176040 29120
rect 175880 29120 176040 29280
rect 175880 29280 176040 29440
rect 175880 29440 176040 29600
rect 175880 29600 176040 29760
rect 175880 29760 176040 29920
rect 175880 29920 176040 30080
rect 175880 30080 176040 30240
rect 175880 30240 176040 30400
rect 175880 30400 176040 30560
rect 175880 30560 176040 30720
rect 175880 30720 176040 30880
rect 175880 30880 176040 31040
rect 175880 31040 176040 31200
rect 175880 31200 176040 31360
rect 175880 31360 176040 31520
rect 175880 31520 176040 31680
rect 175880 31680 176040 31840
rect 175880 31840 176040 32000
rect 175880 32000 176040 32160
rect 175880 32160 176040 32320
rect 175880 32320 176040 32480
rect 175880 32480 176040 32640
rect 175880 32640 176040 32800
rect 175880 32800 176040 32960
rect 175880 32960 176040 33120
rect 175880 33120 176040 33280
rect 175880 33280 176040 33440
rect 175880 33440 176040 33600
rect 175880 33600 176040 33760
rect 175880 33760 176040 33920
rect 175880 33920 176040 34080
rect 175880 34080 176040 34240
rect 175880 34240 176040 34400
rect 175880 34400 176040 34560
rect 175880 34560 176040 34720
rect 175880 34720 176040 34880
rect 175880 34880 176040 35040
rect 175880 35040 176040 35200
rect 175880 35200 176040 35360
rect 175880 35360 176040 35520
rect 175880 35520 176040 35680
rect 175880 35680 176040 35840
rect 175880 35840 176040 36000
rect 175880 36000 176040 36160
rect 175880 36160 176040 36320
rect 175880 36320 176040 36480
rect 175880 36480 176040 36640
rect 175880 36640 176040 36800
rect 175880 36800 176040 36960
rect 175880 36960 176040 37120
rect 175880 37120 176040 37280
rect 175880 37280 176040 37440
rect 175880 37440 176040 37600
rect 175880 37600 176040 37760
rect 175880 37760 176040 37920
rect 175880 37920 176040 38080
rect 175880 38080 176040 38240
rect 175880 38240 176040 38400
rect 175880 38400 176040 38560
rect 175880 38560 176040 38720
rect 175880 38720 176040 38880
rect 175880 38880 176040 39040
rect 175880 39040 176040 39200
rect 175880 39200 176040 39360
rect 175880 39360 176040 39520
rect 175880 39520 176040 39680
rect 175880 39680 176040 39840
rect 175880 39840 176040 40000
rect 175880 40000 176040 40160
rect 175880 40160 176040 40320
rect 176040 27040 176200 27200
rect 176040 27200 176200 27360
rect 176040 27360 176200 27520
rect 176040 27520 176200 27680
rect 176040 27680 176200 27840
rect 176040 27840 176200 28000
rect 176040 28000 176200 28160
rect 176040 28160 176200 28320
rect 176040 28320 176200 28480
rect 176040 28480 176200 28640
rect 176040 28640 176200 28800
rect 176040 28800 176200 28960
rect 176040 28960 176200 29120
rect 176040 29120 176200 29280
rect 176040 29280 176200 29440
rect 176040 29440 176200 29600
rect 176040 29600 176200 29760
rect 176040 29760 176200 29920
rect 176040 29920 176200 30080
rect 176040 30080 176200 30240
rect 176040 30240 176200 30400
rect 176040 30400 176200 30560
rect 176040 30560 176200 30720
rect 176040 30720 176200 30880
rect 176040 30880 176200 31040
rect 176040 31040 176200 31200
rect 176040 31200 176200 31360
rect 176040 31360 176200 31520
rect 176040 31520 176200 31680
rect 176040 31680 176200 31840
rect 176040 31840 176200 32000
rect 176040 32000 176200 32160
rect 176040 32160 176200 32320
rect 176040 32320 176200 32480
rect 176040 32480 176200 32640
rect 176040 32640 176200 32800
rect 176040 32800 176200 32960
rect 176040 32960 176200 33120
rect 176040 33120 176200 33280
rect 176040 33280 176200 33440
rect 176040 33440 176200 33600
rect 176040 33600 176200 33760
rect 176040 33760 176200 33920
rect 176040 33920 176200 34080
rect 176040 34080 176200 34240
rect 176040 34240 176200 34400
rect 176040 34400 176200 34560
rect 176040 34560 176200 34720
rect 176040 34720 176200 34880
rect 176040 34880 176200 35040
rect 176040 35040 176200 35200
rect 176040 35200 176200 35360
rect 176040 35360 176200 35520
rect 176040 35520 176200 35680
rect 176040 35680 176200 35840
rect 176040 35840 176200 36000
rect 176040 36000 176200 36160
rect 176040 36160 176200 36320
rect 176040 36320 176200 36480
rect 176040 36480 176200 36640
rect 176040 36640 176200 36800
rect 176040 36800 176200 36960
rect 176040 36960 176200 37120
rect 176040 37120 176200 37280
rect 176040 37280 176200 37440
rect 176040 37440 176200 37600
rect 176040 37600 176200 37760
rect 176040 37760 176200 37920
rect 176040 37920 176200 38080
rect 176040 38080 176200 38240
rect 176040 38240 176200 38400
rect 176040 38400 176200 38560
rect 176040 38560 176200 38720
rect 176040 38720 176200 38880
rect 176040 38880 176200 39040
rect 176040 39040 176200 39200
rect 176040 39200 176200 39360
rect 176040 39360 176200 39520
rect 176200 26880 176360 27040
rect 176200 27040 176360 27200
rect 176200 27200 176360 27360
rect 176200 27360 176360 27520
rect 176200 27520 176360 27680
rect 176200 27680 176360 27840
rect 176200 27840 176360 28000
rect 176200 28000 176360 28160
rect 176200 28160 176360 28320
rect 176200 28320 176360 28480
rect 176200 28480 176360 28640
rect 176200 28640 176360 28800
rect 176200 28800 176360 28960
rect 176200 28960 176360 29120
rect 176200 29120 176360 29280
rect 176200 29280 176360 29440
rect 176200 29440 176360 29600
rect 176200 29600 176360 29760
rect 176200 29760 176360 29920
rect 176200 29920 176360 30080
rect 176200 30080 176360 30240
rect 176200 30240 176360 30400
rect 176200 30400 176360 30560
rect 176200 30560 176360 30720
rect 176200 30720 176360 30880
rect 176200 30880 176360 31040
rect 176200 31040 176360 31200
rect 176200 31200 176360 31360
rect 176200 31360 176360 31520
rect 176200 31520 176360 31680
rect 176200 31680 176360 31840
rect 176200 31840 176360 32000
rect 176200 32000 176360 32160
rect 176200 32160 176360 32320
rect 176200 32320 176360 32480
rect 176200 32480 176360 32640
rect 176200 32640 176360 32800
rect 176200 32800 176360 32960
rect 176200 32960 176360 33120
rect 176200 33120 176360 33280
rect 176200 33280 176360 33440
rect 176200 33440 176360 33600
rect 176200 33600 176360 33760
rect 176200 33760 176360 33920
rect 176200 33920 176360 34080
rect 176200 34080 176360 34240
rect 176200 34240 176360 34400
rect 176200 34400 176360 34560
rect 176200 34560 176360 34720
rect 176200 34720 176360 34880
rect 176200 34880 176360 35040
rect 176200 35040 176360 35200
rect 176200 35200 176360 35360
rect 176200 35360 176360 35520
rect 176200 35520 176360 35680
rect 176200 35680 176360 35840
rect 176200 35840 176360 36000
rect 176200 36000 176360 36160
rect 176200 36160 176360 36320
rect 176200 36320 176360 36480
rect 176200 36480 176360 36640
rect 176200 36640 176360 36800
rect 176200 36800 176360 36960
rect 176200 36960 176360 37120
rect 176200 37120 176360 37280
rect 176200 37280 176360 37440
rect 176200 37440 176360 37600
rect 176200 37600 176360 37760
rect 176200 37760 176360 37920
rect 176200 37920 176360 38080
rect 176200 38080 176360 38240
rect 176200 38240 176360 38400
rect 176200 38400 176360 38560
rect 176200 38560 176360 38720
rect 176360 26880 176520 27040
rect 176360 27040 176520 27200
rect 176360 27200 176520 27360
rect 176360 27360 176520 27520
rect 176360 27520 176520 27680
rect 176360 27680 176520 27840
rect 176360 27840 176520 28000
rect 176360 28000 176520 28160
rect 176360 28160 176520 28320
rect 176360 28320 176520 28480
rect 176360 28480 176520 28640
rect 176360 28640 176520 28800
rect 176360 28800 176520 28960
rect 176360 28960 176520 29120
rect 176360 29120 176520 29280
rect 176360 29280 176520 29440
rect 176360 29440 176520 29600
rect 176360 29600 176520 29760
rect 176360 29760 176520 29920
rect 176360 29920 176520 30080
rect 176360 30080 176520 30240
rect 176360 30240 176520 30400
rect 176360 30400 176520 30560
rect 176360 30560 176520 30720
rect 176360 30720 176520 30880
rect 176360 30880 176520 31040
rect 176360 31040 176520 31200
rect 176360 31200 176520 31360
rect 176360 31360 176520 31520
rect 176360 31520 176520 31680
rect 176360 31680 176520 31840
rect 176360 31840 176520 32000
rect 176360 32000 176520 32160
rect 176360 32160 176520 32320
rect 176360 32320 176520 32480
rect 176360 32480 176520 32640
rect 176360 32640 176520 32800
rect 176360 32800 176520 32960
rect 176360 32960 176520 33120
rect 176360 33120 176520 33280
rect 176360 33280 176520 33440
rect 176360 33440 176520 33600
rect 176360 33600 176520 33760
rect 176360 33760 176520 33920
rect 176360 33920 176520 34080
rect 176360 34080 176520 34240
rect 176360 34240 176520 34400
rect 176360 34400 176520 34560
rect 176360 34560 176520 34720
rect 176360 34720 176520 34880
rect 176360 34880 176520 35040
rect 176360 35040 176520 35200
rect 176360 35200 176520 35360
rect 176360 35360 176520 35520
rect 176360 35520 176520 35680
rect 176360 35680 176520 35840
rect 176360 35840 176520 36000
rect 176360 36000 176520 36160
rect 176360 36160 176520 36320
rect 176360 36320 176520 36480
rect 176360 36480 176520 36640
rect 176360 36640 176520 36800
rect 176360 36800 176520 36960
rect 176360 36960 176520 37120
rect 176360 37120 176520 37280
rect 176360 37280 176520 37440
rect 176360 37440 176520 37600
rect 176360 37600 176520 37760
rect 176360 37760 176520 37920
rect 176360 37920 176520 38080
rect 176520 26880 176680 27040
rect 176520 27040 176680 27200
rect 176520 27200 176680 27360
rect 176520 27360 176680 27520
rect 176520 27520 176680 27680
rect 176520 27680 176680 27840
rect 176520 27840 176680 28000
rect 176520 28000 176680 28160
rect 176520 28160 176680 28320
rect 176520 28320 176680 28480
rect 176520 28480 176680 28640
rect 176520 28640 176680 28800
rect 176520 28800 176680 28960
rect 176520 28960 176680 29120
rect 176520 29120 176680 29280
rect 176520 29280 176680 29440
rect 176520 29440 176680 29600
rect 176520 29600 176680 29760
rect 176520 29760 176680 29920
rect 176520 29920 176680 30080
rect 176520 30080 176680 30240
rect 176520 30240 176680 30400
rect 176520 30400 176680 30560
rect 176520 30560 176680 30720
rect 176520 30720 176680 30880
rect 176520 30880 176680 31040
rect 176520 31040 176680 31200
rect 176520 31200 176680 31360
rect 176520 31360 176680 31520
rect 176520 31520 176680 31680
rect 176520 31680 176680 31840
rect 176520 31840 176680 32000
rect 176520 32000 176680 32160
rect 176520 32160 176680 32320
rect 176520 32320 176680 32480
rect 176520 32480 176680 32640
rect 176520 32640 176680 32800
rect 176520 32800 176680 32960
rect 176520 32960 176680 33120
rect 176520 33120 176680 33280
rect 176520 33280 176680 33440
rect 176520 33440 176680 33600
rect 176520 33600 176680 33760
rect 176520 33760 176680 33920
rect 176520 33920 176680 34080
rect 176520 34080 176680 34240
rect 176520 34240 176680 34400
rect 176520 34400 176680 34560
rect 176520 34560 176680 34720
rect 176520 34720 176680 34880
rect 176520 34880 176680 35040
rect 176520 35040 176680 35200
rect 176520 35200 176680 35360
rect 176520 35360 176680 35520
rect 176520 35520 176680 35680
rect 176520 35680 176680 35840
rect 176520 35840 176680 36000
rect 176520 36000 176680 36160
rect 176520 36160 176680 36320
rect 176520 36320 176680 36480
rect 176520 36480 176680 36640
rect 176520 36640 176680 36800
rect 176520 36800 176680 36960
rect 176520 36960 176680 37120
rect 176520 37120 176680 37280
rect 176680 26880 176840 27040
rect 176680 27040 176840 27200
rect 176680 27200 176840 27360
rect 176680 27360 176840 27520
rect 176680 27520 176840 27680
rect 176680 27680 176840 27840
rect 176680 27840 176840 28000
rect 176680 28000 176840 28160
rect 176680 28160 176840 28320
rect 176680 28320 176840 28480
rect 176680 28480 176840 28640
rect 176680 28640 176840 28800
rect 176680 28800 176840 28960
rect 176680 28960 176840 29120
rect 176680 29120 176840 29280
rect 176680 29280 176840 29440
rect 176680 29440 176840 29600
rect 176680 29600 176840 29760
rect 176680 29760 176840 29920
rect 176680 29920 176840 30080
rect 176680 30080 176840 30240
rect 176680 30240 176840 30400
rect 176680 30400 176840 30560
rect 176680 30560 176840 30720
rect 176680 30720 176840 30880
rect 176680 30880 176840 31040
rect 176680 31040 176840 31200
rect 176680 31200 176840 31360
rect 176680 31360 176840 31520
rect 176680 31520 176840 31680
rect 176680 31680 176840 31840
rect 176680 31840 176840 32000
rect 176680 32000 176840 32160
rect 176680 32160 176840 32320
rect 176680 32320 176840 32480
rect 176680 32480 176840 32640
rect 176680 32640 176840 32800
rect 176680 32800 176840 32960
rect 176680 32960 176840 33120
rect 176680 33120 176840 33280
rect 176680 33280 176840 33440
rect 176680 33440 176840 33600
rect 176680 33600 176840 33760
rect 176680 33760 176840 33920
rect 176680 33920 176840 34080
rect 176680 34080 176840 34240
rect 176680 34240 176840 34400
rect 176680 34400 176840 34560
rect 176680 34560 176840 34720
rect 176680 34720 176840 34880
rect 176680 34880 176840 35040
rect 176680 35040 176840 35200
rect 176680 35200 176840 35360
rect 176680 35360 176840 35520
rect 176680 35520 176840 35680
rect 176680 35680 176840 35840
rect 176680 35840 176840 36000
rect 176680 36000 176840 36160
rect 176680 36160 176840 36320
rect 176680 36320 176840 36480
rect 176680 36480 176840 36640
rect 176840 26720 177000 26880
rect 176840 26880 177000 27040
rect 176840 27040 177000 27200
rect 176840 27200 177000 27360
rect 176840 27360 177000 27520
rect 176840 27520 177000 27680
rect 176840 27680 177000 27840
rect 176840 27840 177000 28000
rect 176840 28000 177000 28160
rect 176840 28160 177000 28320
rect 176840 28320 177000 28480
rect 176840 28480 177000 28640
rect 176840 28640 177000 28800
rect 176840 28800 177000 28960
rect 176840 28960 177000 29120
rect 176840 29120 177000 29280
rect 176840 29280 177000 29440
rect 176840 29440 177000 29600
rect 176840 29600 177000 29760
rect 176840 29760 177000 29920
rect 176840 29920 177000 30080
rect 176840 30080 177000 30240
rect 176840 30240 177000 30400
rect 176840 30400 177000 30560
rect 176840 30560 177000 30720
rect 176840 30720 177000 30880
rect 176840 30880 177000 31040
rect 176840 31040 177000 31200
rect 176840 31200 177000 31360
rect 176840 31360 177000 31520
rect 176840 31520 177000 31680
rect 176840 31680 177000 31840
rect 176840 31840 177000 32000
rect 176840 32000 177000 32160
rect 176840 32160 177000 32320
rect 176840 32320 177000 32480
rect 176840 32480 177000 32640
rect 176840 32640 177000 32800
rect 176840 32800 177000 32960
rect 176840 32960 177000 33120
rect 176840 33120 177000 33280
rect 176840 33280 177000 33440
rect 176840 33440 177000 33600
rect 176840 33600 177000 33760
rect 176840 33760 177000 33920
rect 176840 33920 177000 34080
rect 176840 34080 177000 34240
rect 176840 34240 177000 34400
rect 176840 34400 177000 34560
rect 176840 34560 177000 34720
rect 176840 34720 177000 34880
rect 176840 34880 177000 35040
rect 176840 35040 177000 35200
rect 176840 35200 177000 35360
rect 176840 35360 177000 35520
rect 176840 35520 177000 35680
rect 176840 35680 177000 35840
rect 177000 26720 177160 26880
rect 177000 26880 177160 27040
rect 177000 27040 177160 27200
rect 177000 27200 177160 27360
rect 177000 27360 177160 27520
rect 177000 27520 177160 27680
rect 177000 27680 177160 27840
rect 177000 27840 177160 28000
rect 177000 28000 177160 28160
rect 177000 28160 177160 28320
rect 177000 28320 177160 28480
rect 177000 28480 177160 28640
rect 177000 28640 177160 28800
rect 177000 28800 177160 28960
rect 177000 28960 177160 29120
rect 177000 29120 177160 29280
rect 177000 29280 177160 29440
rect 177000 29440 177160 29600
rect 177000 29600 177160 29760
rect 177000 29760 177160 29920
rect 177000 29920 177160 30080
rect 177000 30080 177160 30240
rect 177000 30240 177160 30400
rect 177000 30400 177160 30560
rect 177000 30560 177160 30720
rect 177000 30720 177160 30880
rect 177000 30880 177160 31040
rect 177000 31040 177160 31200
rect 177000 31200 177160 31360
rect 177000 31360 177160 31520
rect 177000 31520 177160 31680
rect 177000 31680 177160 31840
rect 177000 31840 177160 32000
rect 177000 32000 177160 32160
rect 177000 32160 177160 32320
rect 177000 32320 177160 32480
rect 177000 32480 177160 32640
rect 177000 32640 177160 32800
rect 177000 32800 177160 32960
rect 177000 32960 177160 33120
rect 177000 33120 177160 33280
rect 177000 33280 177160 33440
rect 177000 33440 177160 33600
rect 177000 33600 177160 33760
rect 177000 33760 177160 33920
rect 177000 33920 177160 34080
rect 177000 34080 177160 34240
rect 177000 34240 177160 34400
rect 177000 34400 177160 34560
rect 177000 34560 177160 34720
rect 177000 34720 177160 34880
rect 177000 34880 177160 35040
rect 177000 35040 177160 35200
rect 177160 26720 177320 26880
rect 177160 26880 177320 27040
rect 177160 27040 177320 27200
rect 177160 27200 177320 27360
rect 177160 27360 177320 27520
rect 177160 27520 177320 27680
rect 177160 27680 177320 27840
rect 177160 27840 177320 28000
rect 177160 28000 177320 28160
rect 177160 28160 177320 28320
rect 177160 28320 177320 28480
rect 177160 28480 177320 28640
rect 177160 28640 177320 28800
rect 177160 28800 177320 28960
rect 177160 28960 177320 29120
rect 177160 29120 177320 29280
rect 177160 29280 177320 29440
rect 177160 29440 177320 29600
rect 177160 29600 177320 29760
rect 177160 29760 177320 29920
rect 177160 29920 177320 30080
rect 177160 30080 177320 30240
rect 177160 30240 177320 30400
rect 177160 30400 177320 30560
rect 177160 30560 177320 30720
rect 177160 30720 177320 30880
rect 177160 30880 177320 31040
rect 177160 31040 177320 31200
rect 177160 31200 177320 31360
rect 177160 31360 177320 31520
rect 177160 31520 177320 31680
rect 177160 31680 177320 31840
rect 177160 31840 177320 32000
rect 177160 32000 177320 32160
rect 177160 32160 177320 32320
rect 177160 32320 177320 32480
rect 177160 32480 177320 32640
rect 177160 32640 177320 32800
rect 177160 32800 177320 32960
rect 177160 32960 177320 33120
rect 177160 33120 177320 33280
rect 177160 33280 177320 33440
rect 177160 33440 177320 33600
rect 177160 33600 177320 33760
rect 177160 33760 177320 33920
rect 177160 33920 177320 34080
rect 177160 34080 177320 34240
rect 177160 34240 177320 34400
rect 177320 26720 177480 26880
rect 177320 26880 177480 27040
rect 177320 27040 177480 27200
rect 177320 27200 177480 27360
rect 177320 27360 177480 27520
rect 177320 27520 177480 27680
rect 177320 27680 177480 27840
rect 177320 27840 177480 28000
rect 177320 28000 177480 28160
rect 177320 28160 177480 28320
rect 177320 28320 177480 28480
rect 177320 28480 177480 28640
rect 177320 28640 177480 28800
rect 177320 28800 177480 28960
rect 177320 28960 177480 29120
rect 177320 29120 177480 29280
rect 177320 29280 177480 29440
rect 177320 29440 177480 29600
rect 177320 29600 177480 29760
rect 177320 29760 177480 29920
rect 177320 29920 177480 30080
rect 177320 30080 177480 30240
rect 177320 30240 177480 30400
rect 177320 30400 177480 30560
rect 177320 30560 177480 30720
rect 177320 30720 177480 30880
rect 177320 30880 177480 31040
rect 177320 31040 177480 31200
rect 177320 31200 177480 31360
rect 177320 31360 177480 31520
rect 177320 31520 177480 31680
rect 177320 31680 177480 31840
rect 177320 31840 177480 32000
rect 177320 32000 177480 32160
rect 177320 32160 177480 32320
rect 177320 32320 177480 32480
rect 177320 32480 177480 32640
rect 177320 32640 177480 32800
rect 177320 32800 177480 32960
rect 177320 32960 177480 33120
rect 177320 33120 177480 33280
rect 177320 33280 177480 33440
rect 177320 33440 177480 33600
rect 177320 33600 177480 33760
rect 177320 33760 177480 33920
rect 177320 33920 177480 34080
rect 177480 26720 177640 26880
rect 177480 26880 177640 27040
rect 177480 27040 177640 27200
rect 177480 27200 177640 27360
rect 177480 27360 177640 27520
rect 177480 27520 177640 27680
rect 177480 27680 177640 27840
rect 177480 27840 177640 28000
rect 177480 28000 177640 28160
rect 177480 28160 177640 28320
rect 177480 28320 177640 28480
rect 177480 28480 177640 28640
rect 177480 28640 177640 28800
rect 177480 28800 177640 28960
rect 177480 28960 177640 29120
rect 177480 29120 177640 29280
rect 177480 29280 177640 29440
rect 177480 29440 177640 29600
rect 177480 29600 177640 29760
rect 177480 29760 177640 29920
rect 177480 29920 177640 30080
rect 177480 30080 177640 30240
rect 177480 30240 177640 30400
rect 177480 30400 177640 30560
rect 177480 30560 177640 30720
rect 177480 30720 177640 30880
rect 177480 30880 177640 31040
rect 177480 31040 177640 31200
rect 177480 31200 177640 31360
rect 177480 31360 177640 31520
rect 177480 31520 177640 31680
rect 177480 31680 177640 31840
rect 177480 31840 177640 32000
rect 177480 32000 177640 32160
rect 177480 32160 177640 32320
rect 177480 32320 177640 32480
rect 177480 32480 177640 32640
rect 177480 32640 177640 32800
rect 177480 32800 177640 32960
rect 177480 32960 177640 33120
rect 177480 33120 177640 33280
rect 177480 33280 177640 33440
rect 177480 33440 177640 33600
rect 177480 33600 177640 33760
rect 177480 33760 177640 33920
rect 177480 33920 177640 34080
rect 177480 34080 177640 34240
rect 177480 34240 177640 34400
rect 177640 26720 177800 26880
rect 177640 26880 177800 27040
rect 177640 27040 177800 27200
rect 177640 27200 177800 27360
rect 177640 27360 177800 27520
rect 177640 27520 177800 27680
rect 177640 27680 177800 27840
rect 177640 27840 177800 28000
rect 177640 28000 177800 28160
rect 177640 28160 177800 28320
rect 177640 28320 177800 28480
rect 177640 28480 177800 28640
rect 177640 28640 177800 28800
rect 177640 28800 177800 28960
rect 177640 28960 177800 29120
rect 177640 29120 177800 29280
rect 177640 29280 177800 29440
rect 177640 29440 177800 29600
rect 177640 29600 177800 29760
rect 177640 29760 177800 29920
rect 177640 29920 177800 30080
rect 177640 30080 177800 30240
rect 177640 30240 177800 30400
rect 177640 30400 177800 30560
rect 177640 30560 177800 30720
rect 177640 30720 177800 30880
rect 177640 30880 177800 31040
rect 177640 31040 177800 31200
rect 177640 31200 177800 31360
rect 177640 31360 177800 31520
rect 177640 31520 177800 31680
rect 177640 31680 177800 31840
rect 177640 31840 177800 32000
rect 177640 32000 177800 32160
rect 177640 32160 177800 32320
rect 177640 32320 177800 32480
rect 177640 32480 177800 32640
rect 177640 32640 177800 32800
rect 177640 32800 177800 32960
rect 177640 32960 177800 33120
rect 177640 33120 177800 33280
rect 177640 33280 177800 33440
rect 177640 33440 177800 33600
rect 177640 33600 177800 33760
rect 177640 33760 177800 33920
rect 177640 33920 177800 34080
rect 177640 34080 177800 34240
rect 177640 34240 177800 34400
rect 177640 34400 177800 34560
rect 177640 34560 177800 34720
rect 177640 34720 177800 34880
rect 177800 26720 177960 26880
rect 177800 26880 177960 27040
rect 177800 27040 177960 27200
rect 177800 27200 177960 27360
rect 177800 27360 177960 27520
rect 177800 27520 177960 27680
rect 177800 27680 177960 27840
rect 177800 27840 177960 28000
rect 177800 28000 177960 28160
rect 177800 28160 177960 28320
rect 177800 28320 177960 28480
rect 177800 28480 177960 28640
rect 177800 28640 177960 28800
rect 177800 28800 177960 28960
rect 177800 28960 177960 29120
rect 177800 29120 177960 29280
rect 177800 29280 177960 29440
rect 177800 29440 177960 29600
rect 177800 29600 177960 29760
rect 177800 29760 177960 29920
rect 177800 29920 177960 30080
rect 177800 30080 177960 30240
rect 177800 30240 177960 30400
rect 177800 30400 177960 30560
rect 177800 30560 177960 30720
rect 177800 30720 177960 30880
rect 177800 30880 177960 31040
rect 177800 31040 177960 31200
rect 177800 31200 177960 31360
rect 177800 31360 177960 31520
rect 177800 31520 177960 31680
rect 177800 31680 177960 31840
rect 177800 31840 177960 32000
rect 177800 32000 177960 32160
rect 177800 32160 177960 32320
rect 177800 32320 177960 32480
rect 177800 32480 177960 32640
rect 177800 32640 177960 32800
rect 177800 32800 177960 32960
rect 177800 32960 177960 33120
rect 177800 33120 177960 33280
rect 177800 33280 177960 33440
rect 177800 33440 177960 33600
rect 177800 33600 177960 33760
rect 177800 33760 177960 33920
rect 177800 33920 177960 34080
rect 177800 34080 177960 34240
rect 177800 34240 177960 34400
rect 177800 34400 177960 34560
rect 177800 34560 177960 34720
rect 177800 34720 177960 34880
rect 177800 34880 177960 35040
rect 177800 35040 177960 35200
rect 177960 26720 178120 26880
rect 177960 26880 178120 27040
rect 177960 27040 178120 27200
rect 177960 27200 178120 27360
rect 177960 27360 178120 27520
rect 177960 27520 178120 27680
rect 177960 27680 178120 27840
rect 177960 27840 178120 28000
rect 177960 28000 178120 28160
rect 177960 28160 178120 28320
rect 177960 28320 178120 28480
rect 177960 28480 178120 28640
rect 177960 28640 178120 28800
rect 177960 28800 178120 28960
rect 177960 28960 178120 29120
rect 177960 29120 178120 29280
rect 177960 29280 178120 29440
rect 177960 29440 178120 29600
rect 177960 29600 178120 29760
rect 177960 29760 178120 29920
rect 177960 29920 178120 30080
rect 177960 30080 178120 30240
rect 177960 30240 178120 30400
rect 177960 30400 178120 30560
rect 177960 30560 178120 30720
rect 177960 30720 178120 30880
rect 177960 30880 178120 31040
rect 177960 31040 178120 31200
rect 177960 31200 178120 31360
rect 177960 31360 178120 31520
rect 177960 31520 178120 31680
rect 177960 31680 178120 31840
rect 177960 31840 178120 32000
rect 177960 32000 178120 32160
rect 177960 32160 178120 32320
rect 177960 32320 178120 32480
rect 177960 32480 178120 32640
rect 177960 32640 178120 32800
rect 177960 32800 178120 32960
rect 177960 32960 178120 33120
rect 177960 33120 178120 33280
rect 177960 33280 178120 33440
rect 177960 33440 178120 33600
rect 177960 33600 178120 33760
rect 177960 33760 178120 33920
rect 177960 33920 178120 34080
rect 177960 34080 178120 34240
rect 177960 34240 178120 34400
rect 177960 34400 178120 34560
rect 177960 34560 178120 34720
rect 177960 34720 178120 34880
rect 177960 34880 178120 35040
rect 177960 35040 178120 35200
rect 177960 35200 178120 35360
rect 177960 35360 178120 35520
rect 178120 26880 178280 27040
rect 178120 27040 178280 27200
rect 178120 27200 178280 27360
rect 178120 27360 178280 27520
rect 178120 27520 178280 27680
rect 178120 27680 178280 27840
rect 178120 27840 178280 28000
rect 178120 28000 178280 28160
rect 178120 28160 178280 28320
rect 178120 28320 178280 28480
rect 178120 28480 178280 28640
rect 178120 28640 178280 28800
rect 178120 28800 178280 28960
rect 178120 28960 178280 29120
rect 178120 29120 178280 29280
rect 178120 29280 178280 29440
rect 178120 29440 178280 29600
rect 178120 29600 178280 29760
rect 178120 29760 178280 29920
rect 178120 29920 178280 30080
rect 178120 30080 178280 30240
rect 178120 30240 178280 30400
rect 178120 30400 178280 30560
rect 178120 30560 178280 30720
rect 178120 30720 178280 30880
rect 178120 30880 178280 31040
rect 178120 31040 178280 31200
rect 178120 31200 178280 31360
rect 178120 31360 178280 31520
rect 178120 31520 178280 31680
rect 178120 31680 178280 31840
rect 178120 31840 178280 32000
rect 178120 32000 178280 32160
rect 178120 32160 178280 32320
rect 178120 32320 178280 32480
rect 178120 32480 178280 32640
rect 178120 32640 178280 32800
rect 178120 32800 178280 32960
rect 178120 32960 178280 33120
rect 178120 33120 178280 33280
rect 178120 33280 178280 33440
rect 178120 33440 178280 33600
rect 178120 33600 178280 33760
rect 178120 33760 178280 33920
rect 178120 33920 178280 34080
rect 178120 34080 178280 34240
rect 178120 34240 178280 34400
rect 178120 34400 178280 34560
rect 178120 34560 178280 34720
rect 178120 34720 178280 34880
rect 178120 34880 178280 35040
rect 178120 35040 178280 35200
rect 178120 35200 178280 35360
rect 178120 35360 178280 35520
rect 178120 35520 178280 35680
rect 178120 35680 178280 35840
rect 178120 35840 178280 36000
rect 178280 26880 178440 27040
rect 178280 27040 178440 27200
rect 178280 27200 178440 27360
rect 178280 27360 178440 27520
rect 178280 27520 178440 27680
rect 178280 27680 178440 27840
rect 178280 27840 178440 28000
rect 178280 28000 178440 28160
rect 178280 28160 178440 28320
rect 178280 28320 178440 28480
rect 178280 28480 178440 28640
rect 178280 28640 178440 28800
rect 178280 28800 178440 28960
rect 178280 28960 178440 29120
rect 178280 29120 178440 29280
rect 178280 29280 178440 29440
rect 178280 29440 178440 29600
rect 178280 29600 178440 29760
rect 178280 29760 178440 29920
rect 178280 29920 178440 30080
rect 178280 30080 178440 30240
rect 178280 30240 178440 30400
rect 178280 30400 178440 30560
rect 178280 30560 178440 30720
rect 178280 30720 178440 30880
rect 178280 30880 178440 31040
rect 178280 31040 178440 31200
rect 178280 31200 178440 31360
rect 178280 31360 178440 31520
rect 178280 31520 178440 31680
rect 178280 31680 178440 31840
rect 178280 31840 178440 32000
rect 178280 32000 178440 32160
rect 178280 32160 178440 32320
rect 178280 32320 178440 32480
rect 178280 32480 178440 32640
rect 178280 32640 178440 32800
rect 178280 32800 178440 32960
rect 178280 32960 178440 33120
rect 178280 33120 178440 33280
rect 178280 33280 178440 33440
rect 178280 33440 178440 33600
rect 178280 33600 178440 33760
rect 178280 33760 178440 33920
rect 178280 33920 178440 34080
rect 178280 34080 178440 34240
rect 178280 34240 178440 34400
rect 178280 34400 178440 34560
rect 178280 34560 178440 34720
rect 178280 34720 178440 34880
rect 178280 34880 178440 35040
rect 178280 35040 178440 35200
rect 178280 35200 178440 35360
rect 178280 35360 178440 35520
rect 178280 35520 178440 35680
rect 178280 35680 178440 35840
rect 178280 35840 178440 36000
rect 178280 36000 178440 36160
rect 178280 36160 178440 36320
rect 178280 36320 178440 36480
rect 178440 26880 178600 27040
rect 178440 27040 178600 27200
rect 178440 27200 178600 27360
rect 178440 27360 178600 27520
rect 178440 27520 178600 27680
rect 178440 27680 178600 27840
rect 178440 27840 178600 28000
rect 178440 28000 178600 28160
rect 178440 28160 178600 28320
rect 178440 28320 178600 28480
rect 178440 28480 178600 28640
rect 178440 28640 178600 28800
rect 178440 28800 178600 28960
rect 178440 28960 178600 29120
rect 178440 29120 178600 29280
rect 178440 29280 178600 29440
rect 178440 29440 178600 29600
rect 178440 29600 178600 29760
rect 178440 29760 178600 29920
rect 178440 29920 178600 30080
rect 178440 30080 178600 30240
rect 178440 30240 178600 30400
rect 178440 30400 178600 30560
rect 178440 30560 178600 30720
rect 178440 30720 178600 30880
rect 178440 30880 178600 31040
rect 178440 31040 178600 31200
rect 178440 31200 178600 31360
rect 178440 31360 178600 31520
rect 178440 31520 178600 31680
rect 178440 31680 178600 31840
rect 178440 31840 178600 32000
rect 178440 32000 178600 32160
rect 178440 32160 178600 32320
rect 178440 32320 178600 32480
rect 178440 32480 178600 32640
rect 178440 32640 178600 32800
rect 178440 32800 178600 32960
rect 178440 32960 178600 33120
rect 178440 33120 178600 33280
rect 178440 33280 178600 33440
rect 178440 33440 178600 33600
rect 178440 33600 178600 33760
rect 178440 33760 178600 33920
rect 178440 33920 178600 34080
rect 178440 34080 178600 34240
rect 178440 34240 178600 34400
rect 178440 34400 178600 34560
rect 178440 34560 178600 34720
rect 178440 34720 178600 34880
rect 178440 34880 178600 35040
rect 178440 35040 178600 35200
rect 178440 35200 178600 35360
rect 178440 35360 178600 35520
rect 178440 35520 178600 35680
rect 178440 35680 178600 35840
rect 178440 35840 178600 36000
rect 178440 36000 178600 36160
rect 178440 36160 178600 36320
rect 178440 36320 178600 36480
rect 178440 36480 178600 36640
rect 178440 36640 178600 36800
rect 178600 27040 178760 27200
rect 178600 27200 178760 27360
rect 178600 27360 178760 27520
rect 178600 27520 178760 27680
rect 178600 27680 178760 27840
rect 178600 27840 178760 28000
rect 178600 28000 178760 28160
rect 178600 28160 178760 28320
rect 178600 28320 178760 28480
rect 178600 28480 178760 28640
rect 178600 28640 178760 28800
rect 178600 28800 178760 28960
rect 178600 28960 178760 29120
rect 178600 29120 178760 29280
rect 178600 29280 178760 29440
rect 178600 29440 178760 29600
rect 178600 29600 178760 29760
rect 178600 29760 178760 29920
rect 178600 29920 178760 30080
rect 178600 30080 178760 30240
rect 178600 30240 178760 30400
rect 178600 30400 178760 30560
rect 178600 30560 178760 30720
rect 178600 30720 178760 30880
rect 178600 30880 178760 31040
rect 178600 31040 178760 31200
rect 178600 31200 178760 31360
rect 178600 31360 178760 31520
rect 178600 31520 178760 31680
rect 178600 31680 178760 31840
rect 178600 31840 178760 32000
rect 178600 32000 178760 32160
rect 178600 32160 178760 32320
rect 178600 32320 178760 32480
rect 178600 32480 178760 32640
rect 178600 32640 178760 32800
rect 178600 32800 178760 32960
rect 178600 32960 178760 33120
rect 178600 33120 178760 33280
rect 178600 33280 178760 33440
rect 178600 33440 178760 33600
rect 178600 33600 178760 33760
rect 178600 33760 178760 33920
rect 178600 33920 178760 34080
rect 178600 34080 178760 34240
rect 178600 34240 178760 34400
rect 178600 34400 178760 34560
rect 178600 34560 178760 34720
rect 178600 34720 178760 34880
rect 178600 34880 178760 35040
rect 178600 35040 178760 35200
rect 178600 35200 178760 35360
rect 178600 35360 178760 35520
rect 178600 35520 178760 35680
rect 178600 35680 178760 35840
rect 178600 35840 178760 36000
rect 178600 36000 178760 36160
rect 178600 36160 178760 36320
rect 178600 36320 178760 36480
rect 178600 36480 178760 36640
rect 178600 36640 178760 36800
rect 178600 36800 178760 36960
rect 178600 36960 178760 37120
rect 178600 37120 178760 37280
rect 178760 27200 178920 27360
rect 178760 27360 178920 27520
rect 178760 27520 178920 27680
rect 178760 27680 178920 27840
rect 178760 27840 178920 28000
rect 178760 28000 178920 28160
rect 178760 28160 178920 28320
rect 178760 28320 178920 28480
rect 178760 28480 178920 28640
rect 178760 28640 178920 28800
rect 178760 28800 178920 28960
rect 178760 28960 178920 29120
rect 178760 29120 178920 29280
rect 178760 29280 178920 29440
rect 178760 29440 178920 29600
rect 178760 29600 178920 29760
rect 178760 29760 178920 29920
rect 178760 29920 178920 30080
rect 178760 30080 178920 30240
rect 178760 30240 178920 30400
rect 178760 30400 178920 30560
rect 178760 30560 178920 30720
rect 178760 30720 178920 30880
rect 178760 30880 178920 31040
rect 178760 31040 178920 31200
rect 178760 31200 178920 31360
rect 178760 31360 178920 31520
rect 178760 31520 178920 31680
rect 178760 31680 178920 31840
rect 178760 31840 178920 32000
rect 178760 32000 178920 32160
rect 178760 32160 178920 32320
rect 178760 32320 178920 32480
rect 178760 32480 178920 32640
rect 178760 32640 178920 32800
rect 178760 32800 178920 32960
rect 178760 32960 178920 33120
rect 178760 33120 178920 33280
rect 178760 33280 178920 33440
rect 178760 33440 178920 33600
rect 178760 33600 178920 33760
rect 178760 33760 178920 33920
rect 178760 33920 178920 34080
rect 178760 34080 178920 34240
rect 178760 34240 178920 34400
rect 178760 34400 178920 34560
rect 178760 34560 178920 34720
rect 178760 34720 178920 34880
rect 178760 34880 178920 35040
rect 178760 35040 178920 35200
rect 178760 35200 178920 35360
rect 178760 35360 178920 35520
rect 178760 35520 178920 35680
rect 178760 35680 178920 35840
rect 178760 35840 178920 36000
rect 178760 36000 178920 36160
rect 178760 36160 178920 36320
rect 178760 36320 178920 36480
rect 178760 36480 178920 36640
rect 178760 36640 178920 36800
rect 178760 36800 178920 36960
rect 178760 36960 178920 37120
rect 178760 37120 178920 37280
rect 178760 37280 178920 37440
rect 178760 37440 178920 37600
rect 178760 37600 178920 37760
rect 178920 27200 179080 27360
rect 178920 27360 179080 27520
rect 178920 27520 179080 27680
rect 178920 27680 179080 27840
rect 178920 27840 179080 28000
rect 178920 28000 179080 28160
rect 178920 28160 179080 28320
rect 178920 28320 179080 28480
rect 178920 28480 179080 28640
rect 178920 28640 179080 28800
rect 178920 28800 179080 28960
rect 178920 28960 179080 29120
rect 178920 29120 179080 29280
rect 178920 29280 179080 29440
rect 178920 29440 179080 29600
rect 178920 29600 179080 29760
rect 178920 29760 179080 29920
rect 178920 29920 179080 30080
rect 178920 30080 179080 30240
rect 178920 30240 179080 30400
rect 178920 30400 179080 30560
rect 178920 30560 179080 30720
rect 178920 30720 179080 30880
rect 178920 30880 179080 31040
rect 178920 31040 179080 31200
rect 178920 31200 179080 31360
rect 178920 31360 179080 31520
rect 178920 31520 179080 31680
rect 178920 31680 179080 31840
rect 178920 31840 179080 32000
rect 178920 32000 179080 32160
rect 178920 32160 179080 32320
rect 178920 32320 179080 32480
rect 178920 32480 179080 32640
rect 178920 32640 179080 32800
rect 178920 32800 179080 32960
rect 178920 32960 179080 33120
rect 178920 33120 179080 33280
rect 178920 33280 179080 33440
rect 178920 33440 179080 33600
rect 178920 33600 179080 33760
rect 178920 33760 179080 33920
rect 178920 33920 179080 34080
rect 178920 34080 179080 34240
rect 178920 34240 179080 34400
rect 178920 34400 179080 34560
rect 178920 34560 179080 34720
rect 178920 34720 179080 34880
rect 178920 34880 179080 35040
rect 178920 35040 179080 35200
rect 178920 35200 179080 35360
rect 178920 35360 179080 35520
rect 178920 35520 179080 35680
rect 178920 35680 179080 35840
rect 178920 35840 179080 36000
rect 178920 36000 179080 36160
rect 178920 36160 179080 36320
rect 178920 36320 179080 36480
rect 178920 36480 179080 36640
rect 178920 36640 179080 36800
rect 178920 36800 179080 36960
rect 178920 36960 179080 37120
rect 178920 37120 179080 37280
rect 178920 37280 179080 37440
rect 178920 37440 179080 37600
rect 178920 37600 179080 37760
rect 178920 37760 179080 37920
rect 178920 37920 179080 38080
rect 179080 27360 179240 27520
rect 179080 27520 179240 27680
rect 179080 27680 179240 27840
rect 179080 27840 179240 28000
rect 179080 28000 179240 28160
rect 179080 28160 179240 28320
rect 179080 28320 179240 28480
rect 179080 28480 179240 28640
rect 179080 28640 179240 28800
rect 179080 28800 179240 28960
rect 179080 28960 179240 29120
rect 179080 29120 179240 29280
rect 179080 29280 179240 29440
rect 179080 29440 179240 29600
rect 179080 29600 179240 29760
rect 179080 29760 179240 29920
rect 179080 29920 179240 30080
rect 179080 30080 179240 30240
rect 179080 30240 179240 30400
rect 179080 30400 179240 30560
rect 179080 30560 179240 30720
rect 179080 30720 179240 30880
rect 179080 30880 179240 31040
rect 179080 31040 179240 31200
rect 179080 31200 179240 31360
rect 179080 31360 179240 31520
rect 179080 31520 179240 31680
rect 179080 31680 179240 31840
rect 179080 31840 179240 32000
rect 179080 32000 179240 32160
rect 179080 32160 179240 32320
rect 179080 32320 179240 32480
rect 179080 32480 179240 32640
rect 179080 32640 179240 32800
rect 179080 32800 179240 32960
rect 179080 32960 179240 33120
rect 179080 33120 179240 33280
rect 179080 33280 179240 33440
rect 179080 33440 179240 33600
rect 179080 33600 179240 33760
rect 179080 33760 179240 33920
rect 179080 33920 179240 34080
rect 179080 34080 179240 34240
rect 179080 34240 179240 34400
rect 179080 34400 179240 34560
rect 179080 34560 179240 34720
rect 179080 34720 179240 34880
rect 179080 34880 179240 35040
rect 179080 35040 179240 35200
rect 179080 35200 179240 35360
rect 179080 35360 179240 35520
rect 179080 35520 179240 35680
rect 179080 35680 179240 35840
rect 179080 35840 179240 36000
rect 179080 36000 179240 36160
rect 179080 36160 179240 36320
rect 179080 36320 179240 36480
rect 179080 36480 179240 36640
rect 179080 36640 179240 36800
rect 179080 36800 179240 36960
rect 179080 36960 179240 37120
rect 179080 37120 179240 37280
rect 179080 37280 179240 37440
rect 179080 37440 179240 37600
rect 179080 37600 179240 37760
rect 179080 37760 179240 37920
rect 179080 37920 179240 38080
rect 179080 38080 179240 38240
rect 179080 38240 179240 38400
rect 179080 38400 179240 38560
rect 179240 27520 179400 27680
rect 179240 27680 179400 27840
rect 179240 27840 179400 28000
rect 179240 28000 179400 28160
rect 179240 28160 179400 28320
rect 179240 28320 179400 28480
rect 179240 28480 179400 28640
rect 179240 28640 179400 28800
rect 179240 28800 179400 28960
rect 179240 28960 179400 29120
rect 179240 29120 179400 29280
rect 179240 29280 179400 29440
rect 179240 29440 179400 29600
rect 179240 29600 179400 29760
rect 179240 29760 179400 29920
rect 179240 29920 179400 30080
rect 179240 30080 179400 30240
rect 179240 30240 179400 30400
rect 179240 30400 179400 30560
rect 179240 30560 179400 30720
rect 179240 30720 179400 30880
rect 179240 30880 179400 31040
rect 179240 31040 179400 31200
rect 179240 31200 179400 31360
rect 179240 31360 179400 31520
rect 179240 31520 179400 31680
rect 179240 31680 179400 31840
rect 179240 31840 179400 32000
rect 179240 32000 179400 32160
rect 179240 32160 179400 32320
rect 179240 32320 179400 32480
rect 179240 32480 179400 32640
rect 179240 32640 179400 32800
rect 179240 32800 179400 32960
rect 179240 32960 179400 33120
rect 179240 33120 179400 33280
rect 179240 33280 179400 33440
rect 179240 33440 179400 33600
rect 179240 33600 179400 33760
rect 179240 33760 179400 33920
rect 179240 33920 179400 34080
rect 179240 34080 179400 34240
rect 179240 34240 179400 34400
rect 179240 34400 179400 34560
rect 179240 34560 179400 34720
rect 179240 34720 179400 34880
rect 179240 34880 179400 35040
rect 179240 35040 179400 35200
rect 179240 35200 179400 35360
rect 179240 35360 179400 35520
rect 179240 35520 179400 35680
rect 179240 35680 179400 35840
rect 179240 35840 179400 36000
rect 179240 36000 179400 36160
rect 179240 36160 179400 36320
rect 179240 36320 179400 36480
rect 179240 36480 179400 36640
rect 179240 36640 179400 36800
rect 179240 36800 179400 36960
rect 179240 36960 179400 37120
rect 179240 37120 179400 37280
rect 179240 37280 179400 37440
rect 179240 37440 179400 37600
rect 179240 37600 179400 37760
rect 179240 37760 179400 37920
rect 179240 37920 179400 38080
rect 179240 38080 179400 38240
rect 179240 38240 179400 38400
rect 179240 38400 179400 38560
rect 179240 38560 179400 38720
rect 179240 38720 179400 38880
rect 179240 38880 179400 39040
rect 179400 27840 179560 28000
rect 179400 28000 179560 28160
rect 179400 28160 179560 28320
rect 179400 28320 179560 28480
rect 179400 28480 179560 28640
rect 179400 28640 179560 28800
rect 179400 28800 179560 28960
rect 179400 29600 179560 29760
rect 179400 29760 179560 29920
rect 179400 29920 179560 30080
rect 179400 30080 179560 30240
rect 179400 30240 179560 30400
rect 179400 30400 179560 30560
rect 179400 30560 179560 30720
rect 179400 30720 179560 30880
rect 179400 30880 179560 31040
rect 179400 31040 179560 31200
rect 179400 31200 179560 31360
rect 179400 31360 179560 31520
rect 179400 31520 179560 31680
rect 179400 31680 179560 31840
rect 179400 31840 179560 32000
rect 179400 32000 179560 32160
rect 179400 32160 179560 32320
rect 179400 32320 179560 32480
rect 179400 32480 179560 32640
rect 179400 32640 179560 32800
rect 179400 32800 179560 32960
rect 179400 32960 179560 33120
rect 179400 33120 179560 33280
rect 179400 33280 179560 33440
rect 179400 33440 179560 33600
rect 179400 33600 179560 33760
rect 179400 33760 179560 33920
rect 179400 33920 179560 34080
rect 179400 34080 179560 34240
rect 179400 34240 179560 34400
rect 179400 34400 179560 34560
rect 179400 34560 179560 34720
rect 179400 34720 179560 34880
rect 179400 34880 179560 35040
rect 179400 35040 179560 35200
rect 179400 35200 179560 35360
rect 179400 35360 179560 35520
rect 179400 35520 179560 35680
rect 179400 35680 179560 35840
rect 179400 35840 179560 36000
rect 179400 36000 179560 36160
rect 179400 36160 179560 36320
rect 179400 36320 179560 36480
rect 179400 36480 179560 36640
rect 179400 36640 179560 36800
rect 179400 36800 179560 36960
rect 179400 36960 179560 37120
rect 179400 37120 179560 37280
rect 179400 37280 179560 37440
rect 179400 37440 179560 37600
rect 179400 37600 179560 37760
rect 179400 37760 179560 37920
rect 179400 37920 179560 38080
rect 179400 38080 179560 38240
rect 179400 38240 179560 38400
rect 179400 38400 179560 38560
rect 179400 38560 179560 38720
rect 179400 38720 179560 38880
rect 179400 38880 179560 39040
rect 179400 39040 179560 39200
rect 179400 39200 179560 39360
rect 179400 39360 179560 39520
rect 179560 30080 179720 30240
rect 179560 30240 179720 30400
rect 179560 30400 179720 30560
rect 179560 30560 179720 30720
rect 179560 30720 179720 30880
rect 179560 30880 179720 31040
rect 179560 31040 179720 31200
rect 179560 31200 179720 31360
rect 179560 31360 179720 31520
rect 179560 31520 179720 31680
rect 179560 31680 179720 31840
rect 179560 31840 179720 32000
rect 179560 32000 179720 32160
rect 179560 32160 179720 32320
rect 179560 32320 179720 32480
rect 179560 32480 179720 32640
rect 179560 32640 179720 32800
rect 179560 32800 179720 32960
rect 179560 32960 179720 33120
rect 179560 33120 179720 33280
rect 179560 33280 179720 33440
rect 179560 33440 179720 33600
rect 179560 33600 179720 33760
rect 179560 33760 179720 33920
rect 179560 33920 179720 34080
rect 179560 34080 179720 34240
rect 179560 34240 179720 34400
rect 179560 34400 179720 34560
rect 179560 34560 179720 34720
rect 179560 34720 179720 34880
rect 179560 34880 179720 35040
rect 179560 35040 179720 35200
rect 179560 35200 179720 35360
rect 179560 35360 179720 35520
rect 179560 35520 179720 35680
rect 179560 35680 179720 35840
rect 179560 35840 179720 36000
rect 179560 36000 179720 36160
rect 179560 36160 179720 36320
rect 179560 36320 179720 36480
rect 179560 36480 179720 36640
rect 179560 36640 179720 36800
rect 179560 36800 179720 36960
rect 179560 36960 179720 37120
rect 179560 37120 179720 37280
rect 179560 37280 179720 37440
rect 179560 37440 179720 37600
rect 179560 37600 179720 37760
rect 179560 37760 179720 37920
rect 179560 37920 179720 38080
rect 179560 38080 179720 38240
rect 179560 38240 179720 38400
rect 179560 38400 179720 38560
rect 179560 38560 179720 38720
rect 179560 38720 179720 38880
rect 179560 38880 179720 39040
rect 179560 39040 179720 39200
rect 179560 39200 179720 39360
rect 179560 39360 179720 39520
rect 179560 39520 179720 39680
rect 179560 39680 179720 39840
rect 179560 39840 179720 40000
rect 179720 30720 179880 30880
rect 179720 30880 179880 31040
rect 179720 31040 179880 31200
rect 179720 31200 179880 31360
rect 179720 31360 179880 31520
rect 179720 31520 179880 31680
rect 179720 31680 179880 31840
rect 179720 31840 179880 32000
rect 179720 32000 179880 32160
rect 179720 32160 179880 32320
rect 179720 32320 179880 32480
rect 179720 32480 179880 32640
rect 179720 32640 179880 32800
rect 179720 32800 179880 32960
rect 179720 32960 179880 33120
rect 179720 33120 179880 33280
rect 179720 33280 179880 33440
rect 179720 33440 179880 33600
rect 179720 33600 179880 33760
rect 179720 33760 179880 33920
rect 179720 33920 179880 34080
rect 179720 34080 179880 34240
rect 179720 34240 179880 34400
rect 179720 34400 179880 34560
rect 179720 34560 179880 34720
rect 179720 34720 179880 34880
rect 179720 34880 179880 35040
rect 179720 35040 179880 35200
rect 179720 35200 179880 35360
rect 179720 35360 179880 35520
rect 179720 35520 179880 35680
rect 179720 35680 179880 35840
rect 179720 35840 179880 36000
rect 179720 36000 179880 36160
rect 179720 36160 179880 36320
rect 179720 36320 179880 36480
rect 179720 36480 179880 36640
rect 179720 36640 179880 36800
rect 179720 36800 179880 36960
rect 179720 36960 179880 37120
rect 179720 37120 179880 37280
rect 179720 37280 179880 37440
rect 179720 37440 179880 37600
rect 179720 37600 179880 37760
rect 179720 37760 179880 37920
rect 179720 37920 179880 38080
rect 179720 38080 179880 38240
rect 179720 38240 179880 38400
rect 179720 38400 179880 38560
rect 179720 38560 179880 38720
rect 179720 38720 179880 38880
rect 179720 38880 179880 39040
rect 179720 39040 179880 39200
rect 179720 39200 179880 39360
rect 179720 39360 179880 39520
rect 179720 39520 179880 39680
rect 179720 39680 179880 39840
rect 179720 39840 179880 40000
rect 179720 40000 179880 40160
rect 179720 40160 179880 40320
rect 179720 40320 179880 40480
rect 179880 31040 180040 31200
rect 179880 31200 180040 31360
rect 179880 31360 180040 31520
rect 179880 31520 180040 31680
rect 179880 31680 180040 31840
rect 179880 31840 180040 32000
rect 179880 32000 180040 32160
rect 179880 32160 180040 32320
rect 179880 32320 180040 32480
rect 179880 32480 180040 32640
rect 179880 32640 180040 32800
rect 179880 32800 180040 32960
rect 179880 32960 180040 33120
rect 179880 33120 180040 33280
rect 179880 33280 180040 33440
rect 179880 33440 180040 33600
rect 179880 33600 180040 33760
rect 179880 33760 180040 33920
rect 179880 33920 180040 34080
rect 179880 34080 180040 34240
rect 179880 34240 180040 34400
rect 179880 34400 180040 34560
rect 179880 34560 180040 34720
rect 179880 34720 180040 34880
rect 179880 34880 180040 35040
rect 179880 35040 180040 35200
rect 179880 35200 180040 35360
rect 179880 35360 180040 35520
rect 179880 35520 180040 35680
rect 179880 35680 180040 35840
rect 179880 35840 180040 36000
rect 179880 36000 180040 36160
rect 179880 36160 180040 36320
rect 179880 36320 180040 36480
rect 179880 36480 180040 36640
rect 179880 36640 180040 36800
rect 179880 36800 180040 36960
rect 179880 36960 180040 37120
rect 179880 37120 180040 37280
rect 179880 37280 180040 37440
rect 179880 37440 180040 37600
rect 179880 37600 180040 37760
rect 179880 37760 180040 37920
rect 179880 37920 180040 38080
rect 179880 38080 180040 38240
rect 179880 38240 180040 38400
rect 179880 38400 180040 38560
rect 179880 38560 180040 38720
rect 179880 38720 180040 38880
rect 179880 38880 180040 39040
rect 179880 39040 180040 39200
rect 179880 39200 180040 39360
rect 179880 39360 180040 39520
rect 179880 39520 180040 39680
rect 179880 39680 180040 39840
rect 179880 39840 180040 40000
rect 179880 40000 180040 40160
rect 179880 40160 180040 40320
rect 179880 40320 180040 40480
rect 179880 40480 180040 40640
rect 179880 40640 180040 40800
rect 179880 40800 180040 40960
rect 180040 31520 180200 31680
rect 180040 31680 180200 31840
rect 180040 31840 180200 32000
rect 180040 32000 180200 32160
rect 180040 32160 180200 32320
rect 180040 32320 180200 32480
rect 180040 32480 180200 32640
rect 180040 32640 180200 32800
rect 180040 32800 180200 32960
rect 180040 32960 180200 33120
rect 180040 33120 180200 33280
rect 180040 33280 180200 33440
rect 180040 33440 180200 33600
rect 180040 33600 180200 33760
rect 180040 33760 180200 33920
rect 180040 33920 180200 34080
rect 180040 34080 180200 34240
rect 180040 34240 180200 34400
rect 180040 34400 180200 34560
rect 180040 34560 180200 34720
rect 180040 34720 180200 34880
rect 180040 34880 180200 35040
rect 180040 35040 180200 35200
rect 180040 35200 180200 35360
rect 180040 35360 180200 35520
rect 180040 35520 180200 35680
rect 180040 35680 180200 35840
rect 180040 35840 180200 36000
rect 180040 36000 180200 36160
rect 180040 36160 180200 36320
rect 180040 36320 180200 36480
rect 180040 36480 180200 36640
rect 180040 36640 180200 36800
rect 180040 36800 180200 36960
rect 180040 36960 180200 37120
rect 180040 37120 180200 37280
rect 180040 37280 180200 37440
rect 180040 37440 180200 37600
rect 180040 37600 180200 37760
rect 180040 37760 180200 37920
rect 180040 37920 180200 38080
rect 180040 38080 180200 38240
rect 180040 38240 180200 38400
rect 180040 38400 180200 38560
rect 180040 38560 180200 38720
rect 180040 38720 180200 38880
rect 180040 38880 180200 39040
rect 180040 39040 180200 39200
rect 180040 39200 180200 39360
rect 180040 39360 180200 39520
rect 180040 39520 180200 39680
rect 180040 39680 180200 39840
rect 180040 39840 180200 40000
rect 180040 40000 180200 40160
rect 180040 40160 180200 40320
rect 180040 40320 180200 40480
rect 180040 40480 180200 40640
rect 180040 40640 180200 40800
rect 180040 40800 180200 40960
rect 180040 40960 180200 41120
rect 180040 41120 180200 41280
rect 180040 41280 180200 41440
rect 180200 32000 180360 32160
rect 180200 32160 180360 32320
rect 180200 32320 180360 32480
rect 180200 32480 180360 32640
rect 180200 32640 180360 32800
rect 180200 32800 180360 32960
rect 180200 32960 180360 33120
rect 180200 33120 180360 33280
rect 180200 33280 180360 33440
rect 180200 33440 180360 33600
rect 180200 33600 180360 33760
rect 180200 33760 180360 33920
rect 180200 33920 180360 34080
rect 180200 34080 180360 34240
rect 180200 34240 180360 34400
rect 180200 34400 180360 34560
rect 180200 34560 180360 34720
rect 180200 34720 180360 34880
rect 180200 34880 180360 35040
rect 180200 35040 180360 35200
rect 180200 35200 180360 35360
rect 180200 35360 180360 35520
rect 180200 35520 180360 35680
rect 180200 35680 180360 35840
rect 180200 35840 180360 36000
rect 180200 36000 180360 36160
rect 180200 36160 180360 36320
rect 180200 36320 180360 36480
rect 180200 36480 180360 36640
rect 180200 36640 180360 36800
rect 180200 36800 180360 36960
rect 180200 36960 180360 37120
rect 180200 37120 180360 37280
rect 180200 37280 180360 37440
rect 180200 37440 180360 37600
rect 180200 37600 180360 37760
rect 180200 37760 180360 37920
rect 180200 37920 180360 38080
rect 180200 38080 180360 38240
rect 180200 38240 180360 38400
rect 180200 38400 180360 38560
rect 180200 38560 180360 38720
rect 180200 38720 180360 38880
rect 180200 38880 180360 39040
rect 180200 39040 180360 39200
rect 180200 39200 180360 39360
rect 180200 39360 180360 39520
rect 180200 39520 180360 39680
rect 180200 39680 180360 39840
rect 180200 39840 180360 40000
rect 180200 40000 180360 40160
rect 180200 40160 180360 40320
rect 180200 40320 180360 40480
rect 180200 40480 180360 40640
rect 180200 40640 180360 40800
rect 180200 40800 180360 40960
rect 180200 40960 180360 41120
rect 180200 41120 180360 41280
rect 180200 41280 180360 41440
rect 180200 41440 180360 41600
rect 180200 41600 180360 41760
rect 180200 41760 180360 41920
rect 180360 32480 180520 32640
rect 180360 32640 180520 32800
rect 180360 32800 180520 32960
rect 180360 32960 180520 33120
rect 180360 33120 180520 33280
rect 180360 33280 180520 33440
rect 180360 33440 180520 33600
rect 180360 33600 180520 33760
rect 180360 33760 180520 33920
rect 180360 33920 180520 34080
rect 180360 34080 180520 34240
rect 180360 34240 180520 34400
rect 180360 34400 180520 34560
rect 180360 34560 180520 34720
rect 180360 34720 180520 34880
rect 180360 34880 180520 35040
rect 180360 35040 180520 35200
rect 180360 35200 180520 35360
rect 180360 35360 180520 35520
rect 180360 35520 180520 35680
rect 180360 35680 180520 35840
rect 180360 35840 180520 36000
rect 180360 36000 180520 36160
rect 180360 36160 180520 36320
rect 180360 36320 180520 36480
rect 180360 36480 180520 36640
rect 180360 36640 180520 36800
rect 180360 36800 180520 36960
rect 180360 36960 180520 37120
rect 180360 37120 180520 37280
rect 180360 37280 180520 37440
rect 180360 37440 180520 37600
rect 180360 37600 180520 37760
rect 180360 37760 180520 37920
rect 180360 37920 180520 38080
rect 180360 38080 180520 38240
rect 180360 38240 180520 38400
rect 180360 38400 180520 38560
rect 180360 38560 180520 38720
rect 180360 38720 180520 38880
rect 180360 38880 180520 39040
rect 180360 39040 180520 39200
rect 180360 39200 180520 39360
rect 180360 39360 180520 39520
rect 180360 39520 180520 39680
rect 180360 39680 180520 39840
rect 180360 39840 180520 40000
rect 180360 40000 180520 40160
rect 180360 40160 180520 40320
rect 180360 40320 180520 40480
rect 180360 40480 180520 40640
rect 180360 40640 180520 40800
rect 180360 40800 180520 40960
rect 180360 40960 180520 41120
rect 180360 41120 180520 41280
rect 180360 41280 180520 41440
rect 180360 41440 180520 41600
rect 180360 41600 180520 41760
rect 180360 41760 180520 41920
rect 180360 41920 180520 42080
rect 180360 42080 180520 42240
rect 180360 42240 180520 42400
rect 180360 42400 180520 42560
rect 180520 32960 180680 33120
rect 180520 33120 180680 33280
rect 180520 33280 180680 33440
rect 180520 33440 180680 33600
rect 180520 33600 180680 33760
rect 180520 33760 180680 33920
rect 180520 33920 180680 34080
rect 180520 34080 180680 34240
rect 180520 34240 180680 34400
rect 180520 34400 180680 34560
rect 180520 34560 180680 34720
rect 180520 34720 180680 34880
rect 180520 34880 180680 35040
rect 180520 35040 180680 35200
rect 180520 35200 180680 35360
rect 180520 35360 180680 35520
rect 180520 35520 180680 35680
rect 180520 35680 180680 35840
rect 180520 35840 180680 36000
rect 180520 36000 180680 36160
rect 180520 36160 180680 36320
rect 180520 36320 180680 36480
rect 180520 36480 180680 36640
rect 180520 36640 180680 36800
rect 180520 36800 180680 36960
rect 180520 36960 180680 37120
rect 180520 37120 180680 37280
rect 180520 37280 180680 37440
rect 180520 37440 180680 37600
rect 180520 37600 180680 37760
rect 180520 37760 180680 37920
rect 180520 37920 180680 38080
rect 180520 38080 180680 38240
rect 180520 38240 180680 38400
rect 180520 38400 180680 38560
rect 180520 38560 180680 38720
rect 180520 38720 180680 38880
rect 180520 38880 180680 39040
rect 180520 39040 180680 39200
rect 180520 39200 180680 39360
rect 180520 39360 180680 39520
rect 180520 39520 180680 39680
rect 180520 39680 180680 39840
rect 180520 39840 180680 40000
rect 180520 40000 180680 40160
rect 180520 40160 180680 40320
rect 180520 40320 180680 40480
rect 180520 40480 180680 40640
rect 180520 40640 180680 40800
rect 180520 40800 180680 40960
rect 180520 40960 180680 41120
rect 180520 41120 180680 41280
rect 180520 41280 180680 41440
rect 180520 41440 180680 41600
rect 180520 41600 180680 41760
rect 180520 41760 180680 41920
rect 180520 41920 180680 42080
rect 180520 42080 180680 42240
rect 180520 42240 180680 42400
rect 180520 42400 180680 42560
rect 180520 42560 180680 42720
rect 180520 42720 180680 42880
rect 180520 42880 180680 43040
rect 180680 33280 180840 33440
rect 180680 33440 180840 33600
rect 180680 33600 180840 33760
rect 180680 33760 180840 33920
rect 180680 33920 180840 34080
rect 180680 34080 180840 34240
rect 180680 34240 180840 34400
rect 180680 34400 180840 34560
rect 180680 34560 180840 34720
rect 180680 34720 180840 34880
rect 180680 34880 180840 35040
rect 180680 35040 180840 35200
rect 180680 35200 180840 35360
rect 180680 35360 180840 35520
rect 180680 35520 180840 35680
rect 180680 35680 180840 35840
rect 180680 35840 180840 36000
rect 180680 36000 180840 36160
rect 180680 36160 180840 36320
rect 180680 36320 180840 36480
rect 180680 36480 180840 36640
rect 180680 36640 180840 36800
rect 180680 36800 180840 36960
rect 180680 36960 180840 37120
rect 180680 37120 180840 37280
rect 180680 37280 180840 37440
rect 180680 37440 180840 37600
rect 180680 37600 180840 37760
rect 180680 37760 180840 37920
rect 180680 37920 180840 38080
rect 180680 38080 180840 38240
rect 180680 38240 180840 38400
rect 180680 38400 180840 38560
rect 180680 38560 180840 38720
rect 180680 38720 180840 38880
rect 180680 38880 180840 39040
rect 180680 39040 180840 39200
rect 180680 39200 180840 39360
rect 180680 39360 180840 39520
rect 180680 39520 180840 39680
rect 180680 39680 180840 39840
rect 180680 39840 180840 40000
rect 180680 40000 180840 40160
rect 180680 40160 180840 40320
rect 180680 40320 180840 40480
rect 180680 40480 180840 40640
rect 180680 40640 180840 40800
rect 180680 40800 180840 40960
rect 180680 40960 180840 41120
rect 180680 41120 180840 41280
rect 180680 41280 180840 41440
rect 180680 41440 180840 41600
rect 180680 41600 180840 41760
rect 180680 41760 180840 41920
rect 180680 41920 180840 42080
rect 180680 42080 180840 42240
rect 180680 42240 180840 42400
rect 180680 42400 180840 42560
rect 180680 42560 180840 42720
rect 180680 42720 180840 42880
rect 180680 42880 180840 43040
rect 180680 43040 180840 43200
rect 180680 43200 180840 43360
rect 180680 43360 180840 43520
rect 180840 33760 181000 33920
rect 180840 33920 181000 34080
rect 180840 34080 181000 34240
rect 180840 34240 181000 34400
rect 180840 34400 181000 34560
rect 180840 34560 181000 34720
rect 180840 34720 181000 34880
rect 180840 34880 181000 35040
rect 180840 35040 181000 35200
rect 180840 35200 181000 35360
rect 180840 35360 181000 35520
rect 180840 35520 181000 35680
rect 180840 35680 181000 35840
rect 180840 35840 181000 36000
rect 180840 36000 181000 36160
rect 180840 36160 181000 36320
rect 180840 36320 181000 36480
rect 180840 36480 181000 36640
rect 180840 36640 181000 36800
rect 180840 36800 181000 36960
rect 180840 36960 181000 37120
rect 180840 37120 181000 37280
rect 180840 37280 181000 37440
rect 180840 37440 181000 37600
rect 180840 37600 181000 37760
rect 180840 37760 181000 37920
rect 180840 37920 181000 38080
rect 180840 38080 181000 38240
rect 180840 38240 181000 38400
rect 180840 38400 181000 38560
rect 180840 38560 181000 38720
rect 180840 38720 181000 38880
rect 180840 38880 181000 39040
rect 180840 39040 181000 39200
rect 180840 39200 181000 39360
rect 180840 39360 181000 39520
rect 180840 39520 181000 39680
rect 180840 39680 181000 39840
rect 180840 39840 181000 40000
rect 180840 40000 181000 40160
rect 180840 40160 181000 40320
rect 180840 40320 181000 40480
rect 180840 40480 181000 40640
rect 180840 40640 181000 40800
rect 180840 40800 181000 40960
rect 180840 40960 181000 41120
rect 180840 41120 181000 41280
rect 180840 41280 181000 41440
rect 180840 41440 181000 41600
rect 180840 41600 181000 41760
rect 180840 41760 181000 41920
rect 180840 41920 181000 42080
rect 180840 42080 181000 42240
rect 180840 42240 181000 42400
rect 180840 42400 181000 42560
rect 180840 42560 181000 42720
rect 180840 42720 181000 42880
rect 180840 42880 181000 43040
rect 180840 43040 181000 43200
rect 180840 43200 181000 43360
rect 180840 43360 181000 43520
rect 180840 43520 181000 43680
rect 180840 43680 181000 43840
rect 180840 43840 181000 44000
rect 181000 34080 181160 34240
rect 181000 34240 181160 34400
rect 181000 34400 181160 34560
rect 181000 34560 181160 34720
rect 181000 34720 181160 34880
rect 181000 34880 181160 35040
rect 181000 35040 181160 35200
rect 181000 35200 181160 35360
rect 181000 35360 181160 35520
rect 181000 35520 181160 35680
rect 181000 35680 181160 35840
rect 181000 35840 181160 36000
rect 181000 36000 181160 36160
rect 181000 36160 181160 36320
rect 181000 36320 181160 36480
rect 181000 36480 181160 36640
rect 181000 36640 181160 36800
rect 181000 36800 181160 36960
rect 181000 36960 181160 37120
rect 181000 37120 181160 37280
rect 181000 37280 181160 37440
rect 181000 37440 181160 37600
rect 181000 37600 181160 37760
rect 181000 37760 181160 37920
rect 181000 37920 181160 38080
rect 181000 38080 181160 38240
rect 181000 38240 181160 38400
rect 181000 38400 181160 38560
rect 181000 38560 181160 38720
rect 181000 38720 181160 38880
rect 181000 38880 181160 39040
rect 181000 39040 181160 39200
rect 181000 39200 181160 39360
rect 181000 39360 181160 39520
rect 181000 39520 181160 39680
rect 181000 39680 181160 39840
rect 181000 39840 181160 40000
rect 181000 40000 181160 40160
rect 181000 40160 181160 40320
rect 181000 40320 181160 40480
rect 181000 40480 181160 40640
rect 181000 40640 181160 40800
rect 181000 40800 181160 40960
rect 181000 40960 181160 41120
rect 181000 41120 181160 41280
rect 181000 41280 181160 41440
rect 181000 41440 181160 41600
rect 181000 41600 181160 41760
rect 181000 41760 181160 41920
rect 181000 41920 181160 42080
rect 181000 42080 181160 42240
rect 181000 42240 181160 42400
rect 181000 42400 181160 42560
rect 181000 42560 181160 42720
rect 181000 42720 181160 42880
rect 181000 42880 181160 43040
rect 181000 43040 181160 43200
rect 181000 43200 181160 43360
rect 181000 43360 181160 43520
rect 181000 43520 181160 43680
rect 181000 43680 181160 43840
rect 181000 43840 181160 44000
rect 181000 44000 181160 44160
rect 181000 44160 181160 44320
rect 181000 44320 181160 44480
rect 181160 34400 181320 34560
rect 181160 34560 181320 34720
rect 181160 34720 181320 34880
rect 181160 34880 181320 35040
rect 181160 35040 181320 35200
rect 181160 35200 181320 35360
rect 181160 35360 181320 35520
rect 181160 35520 181320 35680
rect 181160 35680 181320 35840
rect 181160 35840 181320 36000
rect 181160 36000 181320 36160
rect 181160 36160 181320 36320
rect 181160 36320 181320 36480
rect 181160 36480 181320 36640
rect 181160 36640 181320 36800
rect 181160 36800 181320 36960
rect 181160 36960 181320 37120
rect 181160 37120 181320 37280
rect 181160 37280 181320 37440
rect 181160 37440 181320 37600
rect 181160 37600 181320 37760
rect 181160 37760 181320 37920
rect 181160 37920 181320 38080
rect 181160 38080 181320 38240
rect 181160 38240 181320 38400
rect 181160 38400 181320 38560
rect 181160 38560 181320 38720
rect 181160 38720 181320 38880
rect 181160 38880 181320 39040
rect 181160 39040 181320 39200
rect 181160 39200 181320 39360
rect 181160 39360 181320 39520
rect 181160 39520 181320 39680
rect 181160 39680 181320 39840
rect 181160 39840 181320 40000
rect 181160 40000 181320 40160
rect 181160 40160 181320 40320
rect 181160 40320 181320 40480
rect 181160 40480 181320 40640
rect 181160 40640 181320 40800
rect 181160 40800 181320 40960
rect 181160 40960 181320 41120
rect 181160 41120 181320 41280
rect 181160 41280 181320 41440
rect 181160 41440 181320 41600
rect 181160 41600 181320 41760
rect 181160 41760 181320 41920
rect 181160 41920 181320 42080
rect 181160 42080 181320 42240
rect 181160 42240 181320 42400
rect 181160 42400 181320 42560
rect 181160 42560 181320 42720
rect 181160 42720 181320 42880
rect 181160 42880 181320 43040
rect 181160 43040 181320 43200
rect 181160 43200 181320 43360
rect 181160 43360 181320 43520
rect 181160 43520 181320 43680
rect 181160 43680 181320 43840
rect 181160 43840 181320 44000
rect 181160 44000 181320 44160
rect 181160 44160 181320 44320
rect 181160 44320 181320 44480
rect 181160 44480 181320 44640
rect 181160 44640 181320 44800
rect 181160 44800 181320 44960
rect 181160 44960 181320 45120
rect 181320 34880 181480 35040
rect 181320 35040 181480 35200
rect 181320 35200 181480 35360
rect 181320 35360 181480 35520
rect 181320 35520 181480 35680
rect 181320 35680 181480 35840
rect 181320 35840 181480 36000
rect 181320 36000 181480 36160
rect 181320 36160 181480 36320
rect 181320 36320 181480 36480
rect 181320 36480 181480 36640
rect 181320 36640 181480 36800
rect 181320 36800 181480 36960
rect 181320 36960 181480 37120
rect 181320 37120 181480 37280
rect 181320 37280 181480 37440
rect 181320 37440 181480 37600
rect 181320 37600 181480 37760
rect 181320 37760 181480 37920
rect 181320 37920 181480 38080
rect 181320 38080 181480 38240
rect 181320 38240 181480 38400
rect 181320 38400 181480 38560
rect 181320 38560 181480 38720
rect 181320 38720 181480 38880
rect 181320 38880 181480 39040
rect 181320 39040 181480 39200
rect 181320 39200 181480 39360
rect 181320 39360 181480 39520
rect 181320 39520 181480 39680
rect 181320 39680 181480 39840
rect 181320 39840 181480 40000
rect 181320 40000 181480 40160
rect 181320 40160 181480 40320
rect 181320 40320 181480 40480
rect 181320 40480 181480 40640
rect 181320 40640 181480 40800
rect 181320 40800 181480 40960
rect 181320 40960 181480 41120
rect 181320 41120 181480 41280
rect 181320 41280 181480 41440
rect 181320 41440 181480 41600
rect 181320 41600 181480 41760
rect 181320 41760 181480 41920
rect 181320 41920 181480 42080
rect 181320 42080 181480 42240
rect 181320 42240 181480 42400
rect 181320 42400 181480 42560
rect 181320 42560 181480 42720
rect 181320 42720 181480 42880
rect 181320 42880 181480 43040
rect 181320 43040 181480 43200
rect 181320 43200 181480 43360
rect 181320 43360 181480 43520
rect 181320 43520 181480 43680
rect 181320 43680 181480 43840
rect 181320 43840 181480 44000
rect 181320 44000 181480 44160
rect 181320 44160 181480 44320
rect 181320 44320 181480 44480
rect 181320 44480 181480 44640
rect 181320 44640 181480 44800
rect 181320 44800 181480 44960
rect 181320 44960 181480 45120
rect 181320 45120 181480 45280
rect 181320 45280 181480 45440
rect 181320 45440 181480 45600
rect 181480 35200 181640 35360
rect 181480 35360 181640 35520
rect 181480 35520 181640 35680
rect 181480 35680 181640 35840
rect 181480 35840 181640 36000
rect 181480 36000 181640 36160
rect 181480 36160 181640 36320
rect 181480 36320 181640 36480
rect 181480 36480 181640 36640
rect 181480 36640 181640 36800
rect 181480 36800 181640 36960
rect 181480 36960 181640 37120
rect 181480 37120 181640 37280
rect 181480 37280 181640 37440
rect 181480 37440 181640 37600
rect 181480 37600 181640 37760
rect 181480 37760 181640 37920
rect 181480 37920 181640 38080
rect 181480 38080 181640 38240
rect 181480 38240 181640 38400
rect 181480 38400 181640 38560
rect 181480 38560 181640 38720
rect 181480 38720 181640 38880
rect 181480 38880 181640 39040
rect 181480 39040 181640 39200
rect 181480 39200 181640 39360
rect 181480 39360 181640 39520
rect 181480 39520 181640 39680
rect 181480 39680 181640 39840
rect 181480 39840 181640 40000
rect 181480 40000 181640 40160
rect 181480 40160 181640 40320
rect 181480 40320 181640 40480
rect 181480 40480 181640 40640
rect 181480 40640 181640 40800
rect 181480 40800 181640 40960
rect 181480 40960 181640 41120
rect 181480 41120 181640 41280
rect 181480 41280 181640 41440
rect 181480 41440 181640 41600
rect 181480 41600 181640 41760
rect 181480 41760 181640 41920
rect 181480 41920 181640 42080
rect 181480 42080 181640 42240
rect 181480 42240 181640 42400
rect 181480 42400 181640 42560
rect 181480 42560 181640 42720
rect 181480 42720 181640 42880
rect 181480 42880 181640 43040
rect 181480 43040 181640 43200
rect 181480 43200 181640 43360
rect 181480 43360 181640 43520
rect 181480 43520 181640 43680
rect 181480 43680 181640 43840
rect 181480 43840 181640 44000
rect 181480 44000 181640 44160
rect 181480 44160 181640 44320
rect 181480 44320 181640 44480
rect 181480 44480 181640 44640
rect 181480 44640 181640 44800
rect 181480 44800 181640 44960
rect 181480 44960 181640 45120
rect 181480 45120 181640 45280
rect 181480 45280 181640 45440
rect 181480 45440 181640 45600
rect 181480 45600 181640 45760
rect 181480 45760 181640 45920
rect 181480 45920 181640 46080
rect 181640 35520 181800 35680
rect 181640 35680 181800 35840
rect 181640 35840 181800 36000
rect 181640 36000 181800 36160
rect 181640 36160 181800 36320
rect 181640 36320 181800 36480
rect 181640 36480 181800 36640
rect 181640 36640 181800 36800
rect 181640 36800 181800 36960
rect 181640 36960 181800 37120
rect 181640 37120 181800 37280
rect 181640 37280 181800 37440
rect 181640 37440 181800 37600
rect 181640 37600 181800 37760
rect 181640 37760 181800 37920
rect 181640 37920 181800 38080
rect 181640 38080 181800 38240
rect 181640 38240 181800 38400
rect 181640 38400 181800 38560
rect 181640 38560 181800 38720
rect 181640 38720 181800 38880
rect 181640 38880 181800 39040
rect 181640 39040 181800 39200
rect 181640 39200 181800 39360
rect 181640 39360 181800 39520
rect 181640 39520 181800 39680
rect 181640 39680 181800 39840
rect 181640 39840 181800 40000
rect 181640 40000 181800 40160
rect 181640 40160 181800 40320
rect 181640 40320 181800 40480
rect 181640 40480 181800 40640
rect 181640 40640 181800 40800
rect 181640 40800 181800 40960
rect 181640 40960 181800 41120
rect 181640 41120 181800 41280
rect 181640 41280 181800 41440
rect 181640 41440 181800 41600
rect 181640 41600 181800 41760
rect 181640 41760 181800 41920
rect 181640 41920 181800 42080
rect 181640 42080 181800 42240
rect 181640 42240 181800 42400
rect 181640 42400 181800 42560
rect 181640 42560 181800 42720
rect 181640 42720 181800 42880
rect 181640 42880 181800 43040
rect 181640 43040 181800 43200
rect 181640 43200 181800 43360
rect 181640 43360 181800 43520
rect 181640 43520 181800 43680
rect 181640 43680 181800 43840
rect 181640 43840 181800 44000
rect 181640 44000 181800 44160
rect 181640 44160 181800 44320
rect 181640 44320 181800 44480
rect 181640 44480 181800 44640
rect 181640 44640 181800 44800
rect 181640 44800 181800 44960
rect 181640 44960 181800 45120
rect 181640 45120 181800 45280
rect 181640 45280 181800 45440
rect 181640 45440 181800 45600
rect 181640 45600 181800 45760
rect 181640 45760 181800 45920
rect 181640 45920 181800 46080
rect 181640 46080 181800 46240
rect 181640 46240 181800 46400
rect 181640 46400 181800 46560
rect 181800 36000 181960 36160
rect 181800 36160 181960 36320
rect 181800 36320 181960 36480
rect 181800 36480 181960 36640
rect 181800 36640 181960 36800
rect 181800 36800 181960 36960
rect 181800 36960 181960 37120
rect 181800 37120 181960 37280
rect 181800 37280 181960 37440
rect 181800 37440 181960 37600
rect 181800 37600 181960 37760
rect 181800 37760 181960 37920
rect 181800 37920 181960 38080
rect 181800 38080 181960 38240
rect 181800 38240 181960 38400
rect 181800 38400 181960 38560
rect 181800 38560 181960 38720
rect 181800 38720 181960 38880
rect 181800 38880 181960 39040
rect 181800 39040 181960 39200
rect 181800 39200 181960 39360
rect 181800 39360 181960 39520
rect 181800 39520 181960 39680
rect 181800 39680 181960 39840
rect 181800 39840 181960 40000
rect 181800 40000 181960 40160
rect 181800 40160 181960 40320
rect 181800 40320 181960 40480
rect 181800 40480 181960 40640
rect 181800 40640 181960 40800
rect 181800 40800 181960 40960
rect 181800 40960 181960 41120
rect 181800 41120 181960 41280
rect 181800 41280 181960 41440
rect 181800 41440 181960 41600
rect 181800 41600 181960 41760
rect 181800 41760 181960 41920
rect 181800 41920 181960 42080
rect 181800 42080 181960 42240
rect 181800 42240 181960 42400
rect 181800 42400 181960 42560
rect 181800 42560 181960 42720
rect 181800 42720 181960 42880
rect 181800 42880 181960 43040
rect 181800 43040 181960 43200
rect 181800 43200 181960 43360
rect 181800 43360 181960 43520
rect 181800 43520 181960 43680
rect 181800 43680 181960 43840
rect 181800 43840 181960 44000
rect 181800 44000 181960 44160
rect 181800 44160 181960 44320
rect 181800 44320 181960 44480
rect 181800 44480 181960 44640
rect 181800 44640 181960 44800
rect 181800 44800 181960 44960
rect 181800 44960 181960 45120
rect 181800 45120 181960 45280
rect 181800 45280 181960 45440
rect 181800 45440 181960 45600
rect 181800 45600 181960 45760
rect 181800 45760 181960 45920
rect 181800 45920 181960 46080
rect 181800 46080 181960 46240
rect 181800 46240 181960 46400
rect 181800 46400 181960 46560
rect 181800 46560 181960 46720
rect 181800 46720 181960 46880
rect 181800 46880 181960 47040
rect 181960 36320 182120 36480
rect 181960 36480 182120 36640
rect 181960 36640 182120 36800
rect 181960 36800 182120 36960
rect 181960 36960 182120 37120
rect 181960 37120 182120 37280
rect 181960 37280 182120 37440
rect 181960 37440 182120 37600
rect 181960 37600 182120 37760
rect 181960 37760 182120 37920
rect 181960 37920 182120 38080
rect 181960 38080 182120 38240
rect 181960 38240 182120 38400
rect 181960 38400 182120 38560
rect 181960 38560 182120 38720
rect 181960 38720 182120 38880
rect 181960 38880 182120 39040
rect 181960 39040 182120 39200
rect 181960 39200 182120 39360
rect 181960 39360 182120 39520
rect 181960 39520 182120 39680
rect 181960 39680 182120 39840
rect 181960 39840 182120 40000
rect 181960 40000 182120 40160
rect 181960 40160 182120 40320
rect 181960 40320 182120 40480
rect 181960 40480 182120 40640
rect 181960 40640 182120 40800
rect 181960 40800 182120 40960
rect 181960 40960 182120 41120
rect 181960 41120 182120 41280
rect 181960 41280 182120 41440
rect 181960 41440 182120 41600
rect 181960 41600 182120 41760
rect 181960 41760 182120 41920
rect 181960 41920 182120 42080
rect 181960 42080 182120 42240
rect 181960 42240 182120 42400
rect 181960 42400 182120 42560
rect 181960 42560 182120 42720
rect 181960 42720 182120 42880
rect 181960 42880 182120 43040
rect 181960 43040 182120 43200
rect 181960 43200 182120 43360
rect 181960 43360 182120 43520
rect 181960 43520 182120 43680
rect 181960 43680 182120 43840
rect 181960 43840 182120 44000
rect 181960 44000 182120 44160
rect 181960 44160 182120 44320
rect 181960 44320 182120 44480
rect 181960 44480 182120 44640
rect 181960 44640 182120 44800
rect 181960 44800 182120 44960
rect 181960 44960 182120 45120
rect 181960 45120 182120 45280
rect 181960 45280 182120 45440
rect 181960 45440 182120 45600
rect 181960 45600 182120 45760
rect 181960 45760 182120 45920
rect 181960 45920 182120 46080
rect 181960 46080 182120 46240
rect 181960 46240 182120 46400
rect 181960 46400 182120 46560
rect 181960 46560 182120 46720
rect 181960 46720 182120 46880
rect 181960 46880 182120 47040
rect 181960 47040 182120 47200
rect 181960 47200 182120 47360
rect 181960 47360 182120 47520
rect 182120 36640 182280 36800
rect 182120 36800 182280 36960
rect 182120 36960 182280 37120
rect 182120 37120 182280 37280
rect 182120 37280 182280 37440
rect 182120 37440 182280 37600
rect 182120 37600 182280 37760
rect 182120 37760 182280 37920
rect 182120 37920 182280 38080
rect 182120 38080 182280 38240
rect 182120 38240 182280 38400
rect 182120 38400 182280 38560
rect 182120 38560 182280 38720
rect 182120 38720 182280 38880
rect 182120 38880 182280 39040
rect 182120 39040 182280 39200
rect 182120 39200 182280 39360
rect 182120 39360 182280 39520
rect 182120 39520 182280 39680
rect 182120 39680 182280 39840
rect 182120 39840 182280 40000
rect 182120 40000 182280 40160
rect 182120 40160 182280 40320
rect 182120 40320 182280 40480
rect 182120 40480 182280 40640
rect 182120 40640 182280 40800
rect 182120 40800 182280 40960
rect 182120 40960 182280 41120
rect 182120 41120 182280 41280
rect 182120 41280 182280 41440
rect 182120 41440 182280 41600
rect 182120 41600 182280 41760
rect 182120 41760 182280 41920
rect 182120 41920 182280 42080
rect 182120 42080 182280 42240
rect 182120 42240 182280 42400
rect 182120 42400 182280 42560
rect 182120 42560 182280 42720
rect 182120 42720 182280 42880
rect 182120 42880 182280 43040
rect 182120 43040 182280 43200
rect 182120 43200 182280 43360
rect 182120 43360 182280 43520
rect 182120 43520 182280 43680
rect 182120 43680 182280 43840
rect 182120 43840 182280 44000
rect 182120 44000 182280 44160
rect 182120 44160 182280 44320
rect 182120 44320 182280 44480
rect 182120 44480 182280 44640
rect 182120 44640 182280 44800
rect 182120 44800 182280 44960
rect 182120 44960 182280 45120
rect 182120 45120 182280 45280
rect 182120 45280 182280 45440
rect 182120 45440 182280 45600
rect 182120 45600 182280 45760
rect 182120 45760 182280 45920
rect 182120 45920 182280 46080
rect 182120 46080 182280 46240
rect 182120 46240 182280 46400
rect 182120 46400 182280 46560
rect 182120 46560 182280 46720
rect 182120 46720 182280 46880
rect 182120 46880 182280 47040
rect 182120 47040 182280 47200
rect 182120 47200 182280 47360
rect 182120 47360 182280 47520
rect 182120 47520 182280 47680
rect 182120 47680 182280 47840
rect 182120 47840 182280 48000
rect 182280 37120 182440 37280
rect 182280 37280 182440 37440
rect 182280 37440 182440 37600
rect 182280 37600 182440 37760
rect 182280 37760 182440 37920
rect 182280 37920 182440 38080
rect 182280 38080 182440 38240
rect 182280 38240 182440 38400
rect 182280 38400 182440 38560
rect 182280 38560 182440 38720
rect 182280 38720 182440 38880
rect 182280 38880 182440 39040
rect 182280 39040 182440 39200
rect 182280 39200 182440 39360
rect 182280 39360 182440 39520
rect 182280 39520 182440 39680
rect 182280 39680 182440 39840
rect 182280 39840 182440 40000
rect 182280 40000 182440 40160
rect 182280 40160 182440 40320
rect 182280 40320 182440 40480
rect 182280 40480 182440 40640
rect 182280 40640 182440 40800
rect 182280 40800 182440 40960
rect 182280 40960 182440 41120
rect 182280 41120 182440 41280
rect 182280 41280 182440 41440
rect 182280 41440 182440 41600
rect 182280 41600 182440 41760
rect 182280 41760 182440 41920
rect 182280 41920 182440 42080
rect 182280 42080 182440 42240
rect 182280 42240 182440 42400
rect 182280 42400 182440 42560
rect 182280 42560 182440 42720
rect 182280 42720 182440 42880
rect 182280 42880 182440 43040
rect 182280 43040 182440 43200
rect 182280 43200 182440 43360
rect 182280 43360 182440 43520
rect 182280 43520 182440 43680
rect 182280 43680 182440 43840
rect 182280 43840 182440 44000
rect 182280 44000 182440 44160
rect 182280 44160 182440 44320
rect 182280 44320 182440 44480
rect 182280 44480 182440 44640
rect 182280 44640 182440 44800
rect 182280 44800 182440 44960
rect 182280 44960 182440 45120
rect 182280 45120 182440 45280
rect 182280 45280 182440 45440
rect 182280 45440 182440 45600
rect 182280 45600 182440 45760
rect 182280 45760 182440 45920
rect 182280 45920 182440 46080
rect 182280 46080 182440 46240
rect 182280 46240 182440 46400
rect 182280 46400 182440 46560
rect 182280 46560 182440 46720
rect 182280 46720 182440 46880
rect 182280 46880 182440 47040
rect 182280 47040 182440 47200
rect 182280 47200 182440 47360
rect 182280 47360 182440 47520
rect 182280 47520 182440 47680
rect 182280 47680 182440 47840
rect 182280 47840 182440 48000
rect 182280 48000 182440 48160
rect 182280 48160 182440 48320
rect 182280 48320 182440 48480
rect 182440 37440 182600 37600
rect 182440 37600 182600 37760
rect 182440 37760 182600 37920
rect 182440 37920 182600 38080
rect 182440 38080 182600 38240
rect 182440 38240 182600 38400
rect 182440 38400 182600 38560
rect 182440 38560 182600 38720
rect 182440 38720 182600 38880
rect 182440 38880 182600 39040
rect 182440 39040 182600 39200
rect 182440 39200 182600 39360
rect 182440 39360 182600 39520
rect 182440 39520 182600 39680
rect 182440 39680 182600 39840
rect 182440 39840 182600 40000
rect 182440 40000 182600 40160
rect 182440 40160 182600 40320
rect 182440 40320 182600 40480
rect 182440 40480 182600 40640
rect 182440 40640 182600 40800
rect 182440 40800 182600 40960
rect 182440 40960 182600 41120
rect 182440 41120 182600 41280
rect 182440 41280 182600 41440
rect 182440 41440 182600 41600
rect 182440 41600 182600 41760
rect 182440 41760 182600 41920
rect 182440 41920 182600 42080
rect 182440 42080 182600 42240
rect 182440 42240 182600 42400
rect 182440 42400 182600 42560
rect 182440 42560 182600 42720
rect 182440 42720 182600 42880
rect 182440 42880 182600 43040
rect 182440 43040 182600 43200
rect 182440 43200 182600 43360
rect 182440 43360 182600 43520
rect 182440 43520 182600 43680
rect 182440 43680 182600 43840
rect 182440 43840 182600 44000
rect 182440 44000 182600 44160
rect 182440 44160 182600 44320
rect 182440 44320 182600 44480
rect 182440 44480 182600 44640
rect 182440 44640 182600 44800
rect 182440 44800 182600 44960
rect 182440 44960 182600 45120
rect 182440 45120 182600 45280
rect 182440 45280 182600 45440
rect 182440 45440 182600 45600
rect 182440 45600 182600 45760
rect 182440 45760 182600 45920
rect 182440 45920 182600 46080
rect 182440 46080 182600 46240
rect 182440 46240 182600 46400
rect 182440 46400 182600 46560
rect 182440 46560 182600 46720
rect 182440 46720 182600 46880
rect 182440 46880 182600 47040
rect 182440 47040 182600 47200
rect 182440 47200 182600 47360
rect 182440 47360 182600 47520
rect 182440 47520 182600 47680
rect 182440 47680 182600 47840
rect 182440 47840 182600 48000
rect 182440 48000 182600 48160
rect 182440 48160 182600 48320
rect 182440 48320 182600 48480
rect 182440 48480 182600 48640
rect 182440 48640 182600 48800
rect 182440 48800 182600 48960
rect 182600 37920 182760 38080
rect 182600 38080 182760 38240
rect 182600 38240 182760 38400
rect 182600 38400 182760 38560
rect 182600 38560 182760 38720
rect 182600 38720 182760 38880
rect 182600 38880 182760 39040
rect 182600 39040 182760 39200
rect 182600 39200 182760 39360
rect 182600 39360 182760 39520
rect 182600 39520 182760 39680
rect 182600 39680 182760 39840
rect 182600 39840 182760 40000
rect 182600 40000 182760 40160
rect 182600 40160 182760 40320
rect 182600 40320 182760 40480
rect 182600 40480 182760 40640
rect 182600 40640 182760 40800
rect 182600 40800 182760 40960
rect 182600 40960 182760 41120
rect 182600 41120 182760 41280
rect 182600 41280 182760 41440
rect 182600 41440 182760 41600
rect 182600 41600 182760 41760
rect 182600 41760 182760 41920
rect 182600 41920 182760 42080
rect 182600 42080 182760 42240
rect 182600 42240 182760 42400
rect 182600 42400 182760 42560
rect 182600 42560 182760 42720
rect 182600 42720 182760 42880
rect 182600 42880 182760 43040
rect 182600 43040 182760 43200
rect 182600 43200 182760 43360
rect 182600 43360 182760 43520
rect 182600 43520 182760 43680
rect 182600 43680 182760 43840
rect 182600 43840 182760 44000
rect 182600 44000 182760 44160
rect 182600 44160 182760 44320
rect 182600 44320 182760 44480
rect 182600 44480 182760 44640
rect 182600 44640 182760 44800
rect 182600 44800 182760 44960
rect 182600 44960 182760 45120
rect 182600 45120 182760 45280
rect 182600 45280 182760 45440
rect 182600 45440 182760 45600
rect 182600 45600 182760 45760
rect 182600 45760 182760 45920
rect 182600 45920 182760 46080
rect 182600 46080 182760 46240
rect 182600 46240 182760 46400
rect 182600 46400 182760 46560
rect 182600 46560 182760 46720
rect 182600 46720 182760 46880
rect 182600 46880 182760 47040
rect 182600 47040 182760 47200
rect 182600 47200 182760 47360
rect 182600 47360 182760 47520
rect 182600 47520 182760 47680
rect 182600 47680 182760 47840
rect 182600 47840 182760 48000
rect 182600 48000 182760 48160
rect 182600 48160 182760 48320
rect 182600 48320 182760 48480
rect 182600 48480 182760 48640
rect 182600 48640 182760 48800
rect 182600 48800 182760 48960
rect 182600 48960 182760 49120
rect 182600 49120 182760 49280
rect 182760 38240 182920 38400
rect 182760 38400 182920 38560
rect 182760 38560 182920 38720
rect 182760 38720 182920 38880
rect 182760 38880 182920 39040
rect 182760 39040 182920 39200
rect 182760 39200 182920 39360
rect 182760 39360 182920 39520
rect 182760 39520 182920 39680
rect 182760 39680 182920 39840
rect 182760 39840 182920 40000
rect 182760 40000 182920 40160
rect 182760 40160 182920 40320
rect 182760 40320 182920 40480
rect 182760 40480 182920 40640
rect 182760 40640 182920 40800
rect 182760 40800 182920 40960
rect 182760 40960 182920 41120
rect 182760 41120 182920 41280
rect 182760 41280 182920 41440
rect 182760 41440 182920 41600
rect 182760 41600 182920 41760
rect 182760 41760 182920 41920
rect 182760 41920 182920 42080
rect 182760 42080 182920 42240
rect 182760 42240 182920 42400
rect 182760 42400 182920 42560
rect 182760 42560 182920 42720
rect 182760 42720 182920 42880
rect 182760 42880 182920 43040
rect 182760 43040 182920 43200
rect 182760 43200 182920 43360
rect 182760 43360 182920 43520
rect 182760 43520 182920 43680
rect 182760 43680 182920 43840
rect 182760 43840 182920 44000
rect 182760 44000 182920 44160
rect 182760 44160 182920 44320
rect 182760 44320 182920 44480
rect 182760 44480 182920 44640
rect 182760 44640 182920 44800
rect 182760 44800 182920 44960
rect 182760 44960 182920 45120
rect 182760 45120 182920 45280
rect 182760 45280 182920 45440
rect 182760 45440 182920 45600
rect 182760 45600 182920 45760
rect 182760 45760 182920 45920
rect 182760 45920 182920 46080
rect 182760 46080 182920 46240
rect 182760 46240 182920 46400
rect 182760 46400 182920 46560
rect 182760 46560 182920 46720
rect 182760 46720 182920 46880
rect 182760 46880 182920 47040
rect 182760 47040 182920 47200
rect 182760 47200 182920 47360
rect 182760 47360 182920 47520
rect 182760 47520 182920 47680
rect 182760 47680 182920 47840
rect 182760 47840 182920 48000
rect 182760 48000 182920 48160
rect 182760 48160 182920 48320
rect 182760 48320 182920 48480
rect 182760 48480 182920 48640
rect 182760 48640 182920 48800
rect 182760 48800 182920 48960
rect 182760 48960 182920 49120
rect 182760 49120 182920 49280
rect 182760 49280 182920 49440
rect 182760 49440 182920 49600
rect 182920 38720 183080 38880
rect 182920 38880 183080 39040
rect 182920 39040 183080 39200
rect 182920 39200 183080 39360
rect 182920 39360 183080 39520
rect 182920 39520 183080 39680
rect 182920 39680 183080 39840
rect 182920 39840 183080 40000
rect 182920 40000 183080 40160
rect 182920 40160 183080 40320
rect 182920 40320 183080 40480
rect 182920 40480 183080 40640
rect 182920 40640 183080 40800
rect 182920 40800 183080 40960
rect 182920 40960 183080 41120
rect 182920 41120 183080 41280
rect 182920 41280 183080 41440
rect 182920 41440 183080 41600
rect 182920 41600 183080 41760
rect 182920 41760 183080 41920
rect 182920 41920 183080 42080
rect 182920 42080 183080 42240
rect 182920 42240 183080 42400
rect 182920 42400 183080 42560
rect 182920 42560 183080 42720
rect 182920 42720 183080 42880
rect 182920 42880 183080 43040
rect 182920 43040 183080 43200
rect 182920 43200 183080 43360
rect 182920 43360 183080 43520
rect 182920 43520 183080 43680
rect 182920 43680 183080 43840
rect 182920 43840 183080 44000
rect 182920 44000 183080 44160
rect 182920 44160 183080 44320
rect 182920 44320 183080 44480
rect 182920 44480 183080 44640
rect 182920 44640 183080 44800
rect 182920 44800 183080 44960
rect 182920 44960 183080 45120
rect 182920 45120 183080 45280
rect 182920 45280 183080 45440
rect 182920 45440 183080 45600
rect 182920 45600 183080 45760
rect 182920 45760 183080 45920
rect 182920 45920 183080 46080
rect 182920 46080 183080 46240
rect 182920 46240 183080 46400
rect 182920 46400 183080 46560
rect 182920 46560 183080 46720
rect 182920 46720 183080 46880
rect 182920 46880 183080 47040
rect 182920 47040 183080 47200
rect 182920 47200 183080 47360
rect 182920 47360 183080 47520
rect 182920 47520 183080 47680
rect 182920 47680 183080 47840
rect 182920 47840 183080 48000
rect 182920 48000 183080 48160
rect 182920 48160 183080 48320
rect 182920 48320 183080 48480
rect 182920 48480 183080 48640
rect 182920 48640 183080 48800
rect 182920 48800 183080 48960
rect 182920 48960 183080 49120
rect 182920 49120 183080 49280
rect 182920 49280 183080 49440
rect 182920 49440 183080 49600
rect 182920 49600 183080 49760
rect 182920 49760 183080 49920
rect 182920 49920 183080 50080
rect 183080 39200 183240 39360
rect 183080 39360 183240 39520
rect 183080 39520 183240 39680
rect 183080 39680 183240 39840
rect 183080 39840 183240 40000
rect 183080 40000 183240 40160
rect 183080 40160 183240 40320
rect 183080 40320 183240 40480
rect 183080 40480 183240 40640
rect 183080 40640 183240 40800
rect 183080 40800 183240 40960
rect 183080 40960 183240 41120
rect 183080 41120 183240 41280
rect 183080 41280 183240 41440
rect 183080 41440 183240 41600
rect 183080 41600 183240 41760
rect 183080 41760 183240 41920
rect 183080 41920 183240 42080
rect 183080 42080 183240 42240
rect 183080 42240 183240 42400
rect 183080 42400 183240 42560
rect 183080 42560 183240 42720
rect 183080 42720 183240 42880
rect 183080 42880 183240 43040
rect 183080 43040 183240 43200
rect 183080 43200 183240 43360
rect 183080 43360 183240 43520
rect 183080 43520 183240 43680
rect 183080 43680 183240 43840
rect 183080 43840 183240 44000
rect 183080 44000 183240 44160
rect 183080 44160 183240 44320
rect 183080 44320 183240 44480
rect 183080 44480 183240 44640
rect 183080 44640 183240 44800
rect 183080 44800 183240 44960
rect 183080 44960 183240 45120
rect 183080 45120 183240 45280
rect 183080 45280 183240 45440
rect 183080 45440 183240 45600
rect 183080 45600 183240 45760
rect 183080 45760 183240 45920
rect 183080 45920 183240 46080
rect 183080 46080 183240 46240
rect 183080 46240 183240 46400
rect 183080 46400 183240 46560
rect 183080 46560 183240 46720
rect 183080 46720 183240 46880
rect 183080 46880 183240 47040
rect 183080 47040 183240 47200
rect 183080 47200 183240 47360
rect 183080 47360 183240 47520
rect 183080 47520 183240 47680
rect 183080 47680 183240 47840
rect 183080 47840 183240 48000
rect 183080 48000 183240 48160
rect 183080 48160 183240 48320
rect 183080 48320 183240 48480
rect 183080 48480 183240 48640
rect 183080 48640 183240 48800
rect 183080 48800 183240 48960
rect 183080 48960 183240 49120
rect 183080 49120 183240 49280
rect 183080 49280 183240 49440
rect 183080 49440 183240 49600
rect 183080 49600 183240 49760
rect 183080 49760 183240 49920
rect 183080 49920 183240 50080
rect 183080 50080 183240 50240
rect 183080 50240 183240 50400
rect 183240 39520 183400 39680
rect 183240 39680 183400 39840
rect 183240 39840 183400 40000
rect 183240 40000 183400 40160
rect 183240 40160 183400 40320
rect 183240 40320 183400 40480
rect 183240 40480 183400 40640
rect 183240 40640 183400 40800
rect 183240 40800 183400 40960
rect 183240 40960 183400 41120
rect 183240 41120 183400 41280
rect 183240 41280 183400 41440
rect 183240 41440 183400 41600
rect 183240 41600 183400 41760
rect 183240 41760 183400 41920
rect 183240 41920 183400 42080
rect 183240 42080 183400 42240
rect 183240 42240 183400 42400
rect 183240 42400 183400 42560
rect 183240 42560 183400 42720
rect 183240 42720 183400 42880
rect 183240 42880 183400 43040
rect 183240 43040 183400 43200
rect 183240 43200 183400 43360
rect 183240 43360 183400 43520
rect 183240 43520 183400 43680
rect 183240 43680 183400 43840
rect 183240 43840 183400 44000
rect 183240 44000 183400 44160
rect 183240 44160 183400 44320
rect 183240 44320 183400 44480
rect 183240 44480 183400 44640
rect 183240 44640 183400 44800
rect 183240 44800 183400 44960
rect 183240 44960 183400 45120
rect 183240 45120 183400 45280
rect 183240 45280 183400 45440
rect 183240 45440 183400 45600
rect 183240 45600 183400 45760
rect 183240 45760 183400 45920
rect 183240 45920 183400 46080
rect 183240 46080 183400 46240
rect 183240 46240 183400 46400
rect 183240 46400 183400 46560
rect 183240 46560 183400 46720
rect 183240 46720 183400 46880
rect 183240 46880 183400 47040
rect 183240 47040 183400 47200
rect 183240 47200 183400 47360
rect 183240 47360 183400 47520
rect 183240 47520 183400 47680
rect 183240 47680 183400 47840
rect 183240 47840 183400 48000
rect 183240 48000 183400 48160
rect 183240 48160 183400 48320
rect 183240 48320 183400 48480
rect 183240 48480 183400 48640
rect 183240 48640 183400 48800
rect 183240 48800 183400 48960
rect 183240 48960 183400 49120
rect 183240 49120 183400 49280
rect 183240 49280 183400 49440
rect 183240 49440 183400 49600
rect 183240 49600 183400 49760
rect 183240 49760 183400 49920
rect 183240 49920 183400 50080
rect 183240 50080 183400 50240
rect 183240 50240 183400 50400
rect 183240 50400 183400 50560
rect 183240 50560 183400 50720
rect 183400 40000 183560 40160
rect 183400 40160 183560 40320
rect 183400 40320 183560 40480
rect 183400 40480 183560 40640
rect 183400 40640 183560 40800
rect 183400 40800 183560 40960
rect 183400 40960 183560 41120
rect 183400 41120 183560 41280
rect 183400 41280 183560 41440
rect 183400 41440 183560 41600
rect 183400 41600 183560 41760
rect 183400 41760 183560 41920
rect 183400 41920 183560 42080
rect 183400 42080 183560 42240
rect 183400 42240 183560 42400
rect 183400 42400 183560 42560
rect 183400 42560 183560 42720
rect 183400 42720 183560 42880
rect 183400 42880 183560 43040
rect 183400 43040 183560 43200
rect 183400 43200 183560 43360
rect 183400 43360 183560 43520
rect 183400 43520 183560 43680
rect 183400 43680 183560 43840
rect 183400 43840 183560 44000
rect 183400 44000 183560 44160
rect 183400 44160 183560 44320
rect 183400 44320 183560 44480
rect 183400 44480 183560 44640
rect 183400 44640 183560 44800
rect 183400 44800 183560 44960
rect 183400 44960 183560 45120
rect 183400 45120 183560 45280
rect 183400 45280 183560 45440
rect 183400 45440 183560 45600
rect 183400 45600 183560 45760
rect 183400 45760 183560 45920
rect 183400 45920 183560 46080
rect 183400 46080 183560 46240
rect 183400 46240 183560 46400
rect 183400 46400 183560 46560
rect 183400 46560 183560 46720
rect 183400 46720 183560 46880
rect 183400 46880 183560 47040
rect 183400 47040 183560 47200
rect 183400 47200 183560 47360
rect 183400 47360 183560 47520
rect 183400 47520 183560 47680
rect 183400 47680 183560 47840
rect 183400 47840 183560 48000
rect 183400 48000 183560 48160
rect 183400 48160 183560 48320
rect 183400 48320 183560 48480
rect 183400 48480 183560 48640
rect 183400 48640 183560 48800
rect 183400 48800 183560 48960
rect 183400 48960 183560 49120
rect 183400 49120 183560 49280
rect 183400 49280 183560 49440
rect 183400 49440 183560 49600
rect 183400 49600 183560 49760
rect 183400 49760 183560 49920
rect 183400 49920 183560 50080
rect 183400 50080 183560 50240
rect 183400 50240 183560 50400
rect 183400 50400 183560 50560
rect 183400 50560 183560 50720
rect 183400 50720 183560 50880
rect 183560 40480 183720 40640
rect 183560 40640 183720 40800
rect 183560 40800 183720 40960
rect 183560 40960 183720 41120
rect 183560 41120 183720 41280
rect 183560 41280 183720 41440
rect 183560 41440 183720 41600
rect 183560 41600 183720 41760
rect 183560 41760 183720 41920
rect 183560 41920 183720 42080
rect 183560 42080 183720 42240
rect 183560 42240 183720 42400
rect 183560 42400 183720 42560
rect 183560 42560 183720 42720
rect 183560 42720 183720 42880
rect 183560 42880 183720 43040
rect 183560 43040 183720 43200
rect 183560 43200 183720 43360
rect 183560 43360 183720 43520
rect 183560 43520 183720 43680
rect 183560 43680 183720 43840
rect 183560 43840 183720 44000
rect 183560 44000 183720 44160
rect 183560 44160 183720 44320
rect 183560 44320 183720 44480
rect 183560 44480 183720 44640
rect 183560 44640 183720 44800
rect 183560 44800 183720 44960
rect 183560 44960 183720 45120
rect 183560 45120 183720 45280
rect 183560 45280 183720 45440
rect 183560 45440 183720 45600
rect 183560 45600 183720 45760
rect 183560 45760 183720 45920
rect 183560 45920 183720 46080
rect 183560 46080 183720 46240
rect 183560 46240 183720 46400
rect 183560 46400 183720 46560
rect 183560 46560 183720 46720
rect 183560 46720 183720 46880
rect 183560 46880 183720 47040
rect 183560 47040 183720 47200
rect 183560 47200 183720 47360
rect 183560 47360 183720 47520
rect 183560 47520 183720 47680
rect 183560 47680 183720 47840
rect 183560 47840 183720 48000
rect 183560 48000 183720 48160
rect 183560 48160 183720 48320
rect 183560 48320 183720 48480
rect 183560 48480 183720 48640
rect 183560 48640 183720 48800
rect 183560 48800 183720 48960
rect 183560 48960 183720 49120
rect 183560 49120 183720 49280
rect 183560 49280 183720 49440
rect 183560 49440 183720 49600
rect 183560 49600 183720 49760
rect 183560 49760 183720 49920
rect 183560 49920 183720 50080
rect 183560 50080 183720 50240
rect 183560 50240 183720 50400
rect 183560 50400 183720 50560
rect 183560 50560 183720 50720
rect 183560 50720 183720 50880
rect 183560 50880 183720 51040
rect 183560 51040 183720 51200
rect 183720 40960 183880 41120
rect 183720 41120 183880 41280
rect 183720 41280 183880 41440
rect 183720 41440 183880 41600
rect 183720 41600 183880 41760
rect 183720 41760 183880 41920
rect 183720 41920 183880 42080
rect 183720 42080 183880 42240
rect 183720 42240 183880 42400
rect 183720 42400 183880 42560
rect 183720 42560 183880 42720
rect 183720 42720 183880 42880
rect 183720 42880 183880 43040
rect 183720 43040 183880 43200
rect 183720 43200 183880 43360
rect 183720 43360 183880 43520
rect 183720 43520 183880 43680
rect 183720 43680 183880 43840
rect 183720 43840 183880 44000
rect 183720 44000 183880 44160
rect 183720 44160 183880 44320
rect 183720 44320 183880 44480
rect 183720 44480 183880 44640
rect 183720 44640 183880 44800
rect 183720 44800 183880 44960
rect 183720 44960 183880 45120
rect 183720 45120 183880 45280
rect 183720 45280 183880 45440
rect 183720 45440 183880 45600
rect 183720 45600 183880 45760
rect 183720 45760 183880 45920
rect 183720 45920 183880 46080
rect 183720 46080 183880 46240
rect 183720 46240 183880 46400
rect 183720 46400 183880 46560
rect 183720 46560 183880 46720
rect 183720 46720 183880 46880
rect 183720 46880 183880 47040
rect 183720 47040 183880 47200
rect 183720 47200 183880 47360
rect 183720 47360 183880 47520
rect 183720 47520 183880 47680
rect 183720 47680 183880 47840
rect 183720 47840 183880 48000
rect 183720 48000 183880 48160
rect 183720 48160 183880 48320
rect 183720 48320 183880 48480
rect 183720 48480 183880 48640
rect 183720 48640 183880 48800
rect 183720 48800 183880 48960
rect 183720 48960 183880 49120
rect 183720 49120 183880 49280
rect 183720 49280 183880 49440
rect 183720 49440 183880 49600
rect 183720 49600 183880 49760
rect 183720 49760 183880 49920
rect 183720 49920 183880 50080
rect 183720 50080 183880 50240
rect 183720 50240 183880 50400
rect 183720 50400 183880 50560
rect 183720 50560 183880 50720
rect 183720 50720 183880 50880
rect 183720 50880 183880 51040
rect 183720 51040 183880 51200
rect 183720 51200 183880 51360
rect 183720 51360 183880 51520
rect 183880 41440 184040 41600
rect 183880 41600 184040 41760
rect 183880 41760 184040 41920
rect 183880 41920 184040 42080
rect 183880 42080 184040 42240
rect 183880 42240 184040 42400
rect 183880 42400 184040 42560
rect 183880 42560 184040 42720
rect 183880 42720 184040 42880
rect 183880 42880 184040 43040
rect 183880 43040 184040 43200
rect 183880 43200 184040 43360
rect 183880 43360 184040 43520
rect 183880 43520 184040 43680
rect 183880 43680 184040 43840
rect 183880 43840 184040 44000
rect 183880 44000 184040 44160
rect 183880 44160 184040 44320
rect 183880 44320 184040 44480
rect 183880 44480 184040 44640
rect 183880 44640 184040 44800
rect 183880 44800 184040 44960
rect 183880 44960 184040 45120
rect 183880 45120 184040 45280
rect 183880 45280 184040 45440
rect 183880 45440 184040 45600
rect 183880 45600 184040 45760
rect 183880 45760 184040 45920
rect 183880 45920 184040 46080
rect 183880 46080 184040 46240
rect 183880 46240 184040 46400
rect 183880 46400 184040 46560
rect 183880 46560 184040 46720
rect 183880 46720 184040 46880
rect 183880 46880 184040 47040
rect 183880 47040 184040 47200
rect 183880 47200 184040 47360
rect 183880 47360 184040 47520
rect 183880 47520 184040 47680
rect 183880 47680 184040 47840
rect 183880 47840 184040 48000
rect 183880 48000 184040 48160
rect 183880 48160 184040 48320
rect 183880 48320 184040 48480
rect 183880 48480 184040 48640
rect 183880 48640 184040 48800
rect 183880 48800 184040 48960
rect 183880 48960 184040 49120
rect 183880 49120 184040 49280
rect 183880 49280 184040 49440
rect 183880 49440 184040 49600
rect 183880 49600 184040 49760
rect 183880 49760 184040 49920
rect 183880 49920 184040 50080
rect 183880 50080 184040 50240
rect 183880 50240 184040 50400
rect 183880 50400 184040 50560
rect 183880 50560 184040 50720
rect 183880 50720 184040 50880
rect 183880 50880 184040 51040
rect 183880 51040 184040 51200
rect 183880 51200 184040 51360
rect 183880 51360 184040 51520
rect 183880 51520 184040 51680
rect 184040 41920 184200 42080
rect 184040 42080 184200 42240
rect 184040 42240 184200 42400
rect 184040 42400 184200 42560
rect 184040 42560 184200 42720
rect 184040 42720 184200 42880
rect 184040 42880 184200 43040
rect 184040 43040 184200 43200
rect 184040 43200 184200 43360
rect 184040 43360 184200 43520
rect 184040 43520 184200 43680
rect 184040 43680 184200 43840
rect 184040 43840 184200 44000
rect 184040 44000 184200 44160
rect 184040 44160 184200 44320
rect 184040 44320 184200 44480
rect 184040 44480 184200 44640
rect 184040 44640 184200 44800
rect 184040 44800 184200 44960
rect 184040 44960 184200 45120
rect 184040 45120 184200 45280
rect 184040 45280 184200 45440
rect 184040 45440 184200 45600
rect 184040 45600 184200 45760
rect 184040 45760 184200 45920
rect 184040 45920 184200 46080
rect 184040 46080 184200 46240
rect 184040 46240 184200 46400
rect 184040 46400 184200 46560
rect 184040 46560 184200 46720
rect 184040 46720 184200 46880
rect 184040 46880 184200 47040
rect 184040 47040 184200 47200
rect 184040 47200 184200 47360
rect 184040 47360 184200 47520
rect 184040 47520 184200 47680
rect 184040 47680 184200 47840
rect 184040 47840 184200 48000
rect 184040 48000 184200 48160
rect 184040 48160 184200 48320
rect 184040 48320 184200 48480
rect 184040 48480 184200 48640
rect 184040 48640 184200 48800
rect 184040 48800 184200 48960
rect 184040 48960 184200 49120
rect 184040 49120 184200 49280
rect 184040 49280 184200 49440
rect 184040 49440 184200 49600
rect 184040 49600 184200 49760
rect 184040 49760 184200 49920
rect 184040 49920 184200 50080
rect 184040 50080 184200 50240
rect 184040 50240 184200 50400
rect 184040 50400 184200 50560
rect 184040 50560 184200 50720
rect 184040 50720 184200 50880
rect 184040 50880 184200 51040
rect 184040 51040 184200 51200
rect 184040 51200 184200 51360
rect 184040 51360 184200 51520
rect 184040 51520 184200 51680
rect 184040 51680 184200 51840
rect 184200 42560 184360 42720
rect 184200 42720 184360 42880
rect 184200 42880 184360 43040
rect 184200 43040 184360 43200
rect 184200 43200 184360 43360
rect 184200 43360 184360 43520
rect 184200 43520 184360 43680
rect 184200 43680 184360 43840
rect 184200 43840 184360 44000
rect 184200 44000 184360 44160
rect 184200 44160 184360 44320
rect 184200 44320 184360 44480
rect 184200 44480 184360 44640
rect 184200 44640 184360 44800
rect 184200 44800 184360 44960
rect 184200 44960 184360 45120
rect 184200 45120 184360 45280
rect 184200 45280 184360 45440
rect 184200 45440 184360 45600
rect 184200 45600 184360 45760
rect 184200 45760 184360 45920
rect 184200 45920 184360 46080
rect 184200 46080 184360 46240
rect 184200 46240 184360 46400
rect 184200 46400 184360 46560
rect 184200 46560 184360 46720
rect 184200 46720 184360 46880
rect 184200 46880 184360 47040
rect 184200 47040 184360 47200
rect 184200 47200 184360 47360
rect 184200 47360 184360 47520
rect 184200 47520 184360 47680
rect 184200 47680 184360 47840
rect 184200 47840 184360 48000
rect 184200 48000 184360 48160
rect 184200 48160 184360 48320
rect 184200 48320 184360 48480
rect 184200 48480 184360 48640
rect 184200 48640 184360 48800
rect 184200 48800 184360 48960
rect 184200 48960 184360 49120
rect 184200 49120 184360 49280
rect 184200 49280 184360 49440
rect 184200 49440 184360 49600
rect 184200 49600 184360 49760
rect 184200 49760 184360 49920
rect 184200 49920 184360 50080
rect 184200 50080 184360 50240
rect 184200 50240 184360 50400
rect 184200 50400 184360 50560
rect 184200 50560 184360 50720
rect 184200 50720 184360 50880
rect 184200 50880 184360 51040
rect 184200 51040 184360 51200
rect 184200 51200 184360 51360
rect 184200 51360 184360 51520
rect 184200 51520 184360 51680
rect 184200 51680 184360 51840
rect 184200 51840 184360 52000
rect 184200 52000 184360 52160
rect 184360 43040 184520 43200
rect 184360 43200 184520 43360
rect 184360 43360 184520 43520
rect 184360 43520 184520 43680
rect 184360 43680 184520 43840
rect 184360 43840 184520 44000
rect 184360 44000 184520 44160
rect 184360 44160 184520 44320
rect 184360 44320 184520 44480
rect 184360 44480 184520 44640
rect 184360 44640 184520 44800
rect 184360 44800 184520 44960
rect 184360 44960 184520 45120
rect 184360 45120 184520 45280
rect 184360 45280 184520 45440
rect 184360 45440 184520 45600
rect 184360 45600 184520 45760
rect 184360 45760 184520 45920
rect 184360 45920 184520 46080
rect 184360 46080 184520 46240
rect 184360 46240 184520 46400
rect 184360 46400 184520 46560
rect 184360 46560 184520 46720
rect 184360 46720 184520 46880
rect 184360 46880 184520 47040
rect 184360 47040 184520 47200
rect 184360 47200 184520 47360
rect 184360 47360 184520 47520
rect 184360 47520 184520 47680
rect 184360 47680 184520 47840
rect 184360 47840 184520 48000
rect 184360 48000 184520 48160
rect 184360 48160 184520 48320
rect 184360 48320 184520 48480
rect 184360 48480 184520 48640
rect 184360 48640 184520 48800
rect 184360 48800 184520 48960
rect 184360 48960 184520 49120
rect 184360 49120 184520 49280
rect 184360 49280 184520 49440
rect 184360 49440 184520 49600
rect 184360 49600 184520 49760
rect 184360 49760 184520 49920
rect 184360 49920 184520 50080
rect 184360 50080 184520 50240
rect 184360 50240 184520 50400
rect 184360 50400 184520 50560
rect 184360 50560 184520 50720
rect 184360 50720 184520 50880
rect 184360 50880 184520 51040
rect 184360 51040 184520 51200
rect 184360 51200 184520 51360
rect 184360 51360 184520 51520
rect 184360 51520 184520 51680
rect 184360 51680 184520 51840
rect 184360 51840 184520 52000
rect 184360 52000 184520 52160
rect 184360 52160 184520 52320
rect 184520 43520 184680 43680
rect 184520 43680 184680 43840
rect 184520 43840 184680 44000
rect 184520 44000 184680 44160
rect 184520 44160 184680 44320
rect 184520 44320 184680 44480
rect 184520 44480 184680 44640
rect 184520 44640 184680 44800
rect 184520 44800 184680 44960
rect 184520 44960 184680 45120
rect 184520 45120 184680 45280
rect 184520 45280 184680 45440
rect 184520 45440 184680 45600
rect 184520 45600 184680 45760
rect 184520 45760 184680 45920
rect 184520 45920 184680 46080
rect 184520 46080 184680 46240
rect 184520 46240 184680 46400
rect 184520 46400 184680 46560
rect 184520 46560 184680 46720
rect 184520 46720 184680 46880
rect 184520 46880 184680 47040
rect 184520 47040 184680 47200
rect 184520 47200 184680 47360
rect 184520 47360 184680 47520
rect 184520 47520 184680 47680
rect 184520 47680 184680 47840
rect 184520 47840 184680 48000
rect 184520 48000 184680 48160
rect 184520 48160 184680 48320
rect 184520 48320 184680 48480
rect 184520 48480 184680 48640
rect 184520 48640 184680 48800
rect 184520 48800 184680 48960
rect 184520 48960 184680 49120
rect 184520 49120 184680 49280
rect 184520 49280 184680 49440
rect 184520 49440 184680 49600
rect 184520 49600 184680 49760
rect 184520 49760 184680 49920
rect 184520 49920 184680 50080
rect 184520 50080 184680 50240
rect 184520 50240 184680 50400
rect 184520 50400 184680 50560
rect 184520 50560 184680 50720
rect 184520 50720 184680 50880
rect 184520 50880 184680 51040
rect 184520 51040 184680 51200
rect 184520 51200 184680 51360
rect 184520 51360 184680 51520
rect 184520 51520 184680 51680
rect 184520 51680 184680 51840
rect 184520 51840 184680 52000
rect 184520 52000 184680 52160
rect 184520 52160 184680 52320
rect 184680 44160 184840 44320
rect 184680 44320 184840 44480
rect 184680 44480 184840 44640
rect 184680 44640 184840 44800
rect 184680 44800 184840 44960
rect 184680 44960 184840 45120
rect 184680 45120 184840 45280
rect 184680 45280 184840 45440
rect 184680 45440 184840 45600
rect 184680 45600 184840 45760
rect 184680 45760 184840 45920
rect 184680 45920 184840 46080
rect 184680 46080 184840 46240
rect 184680 46240 184840 46400
rect 184680 46400 184840 46560
rect 184680 46560 184840 46720
rect 184680 46720 184840 46880
rect 184680 46880 184840 47040
rect 184680 47040 184840 47200
rect 184680 47200 184840 47360
rect 184680 47360 184840 47520
rect 184680 47520 184840 47680
rect 184680 47680 184840 47840
rect 184680 47840 184840 48000
rect 184680 48000 184840 48160
rect 184680 48160 184840 48320
rect 184680 48320 184840 48480
rect 184680 48480 184840 48640
rect 184680 48640 184840 48800
rect 184680 48800 184840 48960
rect 184680 48960 184840 49120
rect 184680 49120 184840 49280
rect 184680 49280 184840 49440
rect 184680 49440 184840 49600
rect 184680 49600 184840 49760
rect 184680 49760 184840 49920
rect 184680 49920 184840 50080
rect 184680 50080 184840 50240
rect 184680 50240 184840 50400
rect 184680 50400 184840 50560
rect 184680 50560 184840 50720
rect 184680 50720 184840 50880
rect 184680 50880 184840 51040
rect 184680 51040 184840 51200
rect 184680 51200 184840 51360
rect 184680 51360 184840 51520
rect 184680 51520 184840 51680
rect 184680 51680 184840 51840
rect 184680 51840 184840 52000
rect 184680 52000 184840 52160
rect 184680 52160 184840 52320
rect 184680 52320 184840 52480
rect 184840 44640 185000 44800
rect 184840 44800 185000 44960
rect 184840 44960 185000 45120
rect 184840 45120 185000 45280
rect 184840 45280 185000 45440
rect 184840 45440 185000 45600
rect 184840 45600 185000 45760
rect 184840 45760 185000 45920
rect 184840 45920 185000 46080
rect 184840 46080 185000 46240
rect 184840 46240 185000 46400
rect 184840 46400 185000 46560
rect 184840 46560 185000 46720
rect 184840 46720 185000 46880
rect 184840 46880 185000 47040
rect 184840 47040 185000 47200
rect 184840 47200 185000 47360
rect 184840 47360 185000 47520
rect 184840 47520 185000 47680
rect 184840 47680 185000 47840
rect 184840 47840 185000 48000
rect 184840 48000 185000 48160
rect 184840 48160 185000 48320
rect 184840 48320 185000 48480
rect 184840 48480 185000 48640
rect 184840 48640 185000 48800
rect 184840 48800 185000 48960
rect 184840 48960 185000 49120
rect 184840 49120 185000 49280
rect 184840 49280 185000 49440
rect 184840 49440 185000 49600
rect 184840 49600 185000 49760
rect 184840 49760 185000 49920
rect 184840 49920 185000 50080
rect 184840 50080 185000 50240
rect 184840 50240 185000 50400
rect 184840 50400 185000 50560
rect 184840 50560 185000 50720
rect 184840 50720 185000 50880
rect 184840 50880 185000 51040
rect 184840 51040 185000 51200
rect 184840 51200 185000 51360
rect 184840 51360 185000 51520
rect 184840 51520 185000 51680
rect 184840 51680 185000 51840
rect 184840 51840 185000 52000
rect 184840 52000 185000 52160
rect 184840 52160 185000 52320
rect 184840 52320 185000 52480
rect 184840 52480 185000 52640
rect 185000 45280 185160 45440
rect 185000 45440 185160 45600
rect 185000 45600 185160 45760
rect 185000 45760 185160 45920
rect 185000 45920 185160 46080
rect 185000 46080 185160 46240
rect 185000 46240 185160 46400
rect 185000 46400 185160 46560
rect 185000 46560 185160 46720
rect 185000 46720 185160 46880
rect 185000 46880 185160 47040
rect 185000 47040 185160 47200
rect 185000 47200 185160 47360
rect 185000 47360 185160 47520
rect 185000 47520 185160 47680
rect 185000 47680 185160 47840
rect 185000 47840 185160 48000
rect 185000 48000 185160 48160
rect 185000 48160 185160 48320
rect 185000 48320 185160 48480
rect 185000 48480 185160 48640
rect 185000 48640 185160 48800
rect 185000 48800 185160 48960
rect 185000 48960 185160 49120
rect 185000 49120 185160 49280
rect 185000 49280 185160 49440
rect 185000 49440 185160 49600
rect 185000 49600 185160 49760
rect 185000 49760 185160 49920
rect 185000 49920 185160 50080
rect 185000 50080 185160 50240
rect 185000 50240 185160 50400
rect 185000 50400 185160 50560
rect 185000 50560 185160 50720
rect 185000 50720 185160 50880
rect 185000 50880 185160 51040
rect 185000 51040 185160 51200
rect 185000 51200 185160 51360
rect 185000 51360 185160 51520
rect 185000 51520 185160 51680
rect 185000 51680 185160 51840
rect 185000 51840 185160 52000
rect 185000 52000 185160 52160
rect 185000 52160 185160 52320
rect 185000 52320 185160 52480
rect 185000 52480 185160 52640
rect 185160 44640 185320 44800
rect 185160 44800 185320 44960
rect 185160 44960 185320 45120
rect 185160 45120 185320 45280
rect 185160 45280 185320 45440
rect 185160 45440 185320 45600
rect 185160 45600 185320 45760
rect 185160 45760 185320 45920
rect 185160 45920 185320 46080
rect 185160 46080 185320 46240
rect 185160 46240 185320 46400
rect 185160 46400 185320 46560
rect 185160 46560 185320 46720
rect 185160 46720 185320 46880
rect 185160 46880 185320 47040
rect 185160 47040 185320 47200
rect 185160 47200 185320 47360
rect 185160 47360 185320 47520
rect 185160 47520 185320 47680
rect 185160 47680 185320 47840
rect 185160 47840 185320 48000
rect 185160 48000 185320 48160
rect 185160 48160 185320 48320
rect 185160 48320 185320 48480
rect 185160 48480 185320 48640
rect 185160 48640 185320 48800
rect 185160 48800 185320 48960
rect 185160 48960 185320 49120
rect 185160 49120 185320 49280
rect 185160 49280 185320 49440
rect 185160 49440 185320 49600
rect 185160 49600 185320 49760
rect 185160 49760 185320 49920
rect 185160 49920 185320 50080
rect 185160 50080 185320 50240
rect 185160 50240 185320 50400
rect 185160 50400 185320 50560
rect 185160 50560 185320 50720
rect 185160 50720 185320 50880
rect 185160 50880 185320 51040
rect 185160 51040 185320 51200
rect 185160 51200 185320 51360
rect 185160 51360 185320 51520
rect 185160 51520 185320 51680
rect 185160 51680 185320 51840
rect 185160 51840 185320 52000
rect 185160 52000 185320 52160
rect 185160 52160 185320 52320
rect 185160 52320 185320 52480
rect 185160 52480 185320 52640
rect 185160 52640 185320 52800
rect 185320 43520 185480 43680
rect 185320 43680 185480 43840
rect 185320 43840 185480 44000
rect 185320 44000 185480 44160
rect 185320 44160 185480 44320
rect 185320 44320 185480 44480
rect 185320 44480 185480 44640
rect 185320 44640 185480 44800
rect 185320 44800 185480 44960
rect 185320 44960 185480 45120
rect 185320 45120 185480 45280
rect 185320 45280 185480 45440
rect 185320 45440 185480 45600
rect 185320 45600 185480 45760
rect 185320 45760 185480 45920
rect 185320 45920 185480 46080
rect 185320 46080 185480 46240
rect 185320 46240 185480 46400
rect 185320 46400 185480 46560
rect 185320 46560 185480 46720
rect 185320 46720 185480 46880
rect 185320 46880 185480 47040
rect 185320 47040 185480 47200
rect 185320 47200 185480 47360
rect 185320 47360 185480 47520
rect 185320 47520 185480 47680
rect 185320 47680 185480 47840
rect 185320 47840 185480 48000
rect 185320 48000 185480 48160
rect 185320 48160 185480 48320
rect 185320 48320 185480 48480
rect 185320 48480 185480 48640
rect 185320 48640 185480 48800
rect 185320 48800 185480 48960
rect 185320 48960 185480 49120
rect 185320 49120 185480 49280
rect 185320 49280 185480 49440
rect 185320 49440 185480 49600
rect 185320 49600 185480 49760
rect 185320 49760 185480 49920
rect 185320 49920 185480 50080
rect 185320 50080 185480 50240
rect 185320 50240 185480 50400
rect 185320 50400 185480 50560
rect 185320 50560 185480 50720
rect 185320 50720 185480 50880
rect 185320 50880 185480 51040
rect 185320 51040 185480 51200
rect 185320 51200 185480 51360
rect 185320 51360 185480 51520
rect 185320 51520 185480 51680
rect 185320 51680 185480 51840
rect 185320 51840 185480 52000
rect 185320 52000 185480 52160
rect 185320 52160 185480 52320
rect 185320 52320 185480 52480
rect 185320 52480 185480 52640
rect 185320 52640 185480 52800
rect 185480 42400 185640 42560
rect 185480 42560 185640 42720
rect 185480 42720 185640 42880
rect 185480 42880 185640 43040
rect 185480 43040 185640 43200
rect 185480 43200 185640 43360
rect 185480 43360 185640 43520
rect 185480 43520 185640 43680
rect 185480 43680 185640 43840
rect 185480 43840 185640 44000
rect 185480 44000 185640 44160
rect 185480 44160 185640 44320
rect 185480 44320 185640 44480
rect 185480 44480 185640 44640
rect 185480 44640 185640 44800
rect 185480 44800 185640 44960
rect 185480 44960 185640 45120
rect 185480 45120 185640 45280
rect 185480 45280 185640 45440
rect 185480 45440 185640 45600
rect 185480 45600 185640 45760
rect 185480 45760 185640 45920
rect 185480 45920 185640 46080
rect 185480 46080 185640 46240
rect 185480 46240 185640 46400
rect 185480 46400 185640 46560
rect 185480 46560 185640 46720
rect 185480 46720 185640 46880
rect 185480 46880 185640 47040
rect 185480 47040 185640 47200
rect 185480 47200 185640 47360
rect 185480 47360 185640 47520
rect 185480 47520 185640 47680
rect 185480 47680 185640 47840
rect 185480 47840 185640 48000
rect 185480 48000 185640 48160
rect 185480 48160 185640 48320
rect 185480 48320 185640 48480
rect 185480 48480 185640 48640
rect 185480 48640 185640 48800
rect 185480 48800 185640 48960
rect 185480 48960 185640 49120
rect 185480 49120 185640 49280
rect 185480 49280 185640 49440
rect 185480 49440 185640 49600
rect 185480 49600 185640 49760
rect 185480 49760 185640 49920
rect 185480 49920 185640 50080
rect 185480 50080 185640 50240
rect 185480 50240 185640 50400
rect 185480 50400 185640 50560
rect 185480 50560 185640 50720
rect 185480 50720 185640 50880
rect 185480 50880 185640 51040
rect 185480 51040 185640 51200
rect 185480 51200 185640 51360
rect 185480 51360 185640 51520
rect 185480 51520 185640 51680
rect 185480 51680 185640 51840
rect 185480 51840 185640 52000
rect 185480 52000 185640 52160
rect 185480 52160 185640 52320
rect 185480 52320 185640 52480
rect 185480 52480 185640 52640
rect 185480 52640 185640 52800
rect 185640 41440 185800 41600
rect 185640 41600 185800 41760
rect 185640 41760 185800 41920
rect 185640 41920 185800 42080
rect 185640 42080 185800 42240
rect 185640 42240 185800 42400
rect 185640 42400 185800 42560
rect 185640 42560 185800 42720
rect 185640 42720 185800 42880
rect 185640 42880 185800 43040
rect 185640 43040 185800 43200
rect 185640 43200 185800 43360
rect 185640 43360 185800 43520
rect 185640 43520 185800 43680
rect 185640 43680 185800 43840
rect 185640 43840 185800 44000
rect 185640 44000 185800 44160
rect 185640 44160 185800 44320
rect 185640 44320 185800 44480
rect 185640 44480 185800 44640
rect 185640 44640 185800 44800
rect 185640 44800 185800 44960
rect 185640 44960 185800 45120
rect 185640 45120 185800 45280
rect 185640 45280 185800 45440
rect 185640 45440 185800 45600
rect 185640 45600 185800 45760
rect 185640 45760 185800 45920
rect 185640 45920 185800 46080
rect 185640 46080 185800 46240
rect 185640 46240 185800 46400
rect 185640 46400 185800 46560
rect 185640 46560 185800 46720
rect 185640 46720 185800 46880
rect 185640 46880 185800 47040
rect 185640 47040 185800 47200
rect 185640 47200 185800 47360
rect 185640 47360 185800 47520
rect 185640 47520 185800 47680
rect 185640 47680 185800 47840
rect 185640 47840 185800 48000
rect 185640 48000 185800 48160
rect 185640 48160 185800 48320
rect 185640 48320 185800 48480
rect 185640 48480 185800 48640
rect 185640 48640 185800 48800
rect 185640 48800 185800 48960
rect 185640 48960 185800 49120
rect 185640 49120 185800 49280
rect 185640 49280 185800 49440
rect 185640 49440 185800 49600
rect 185640 49600 185800 49760
rect 185640 49760 185800 49920
rect 185640 49920 185800 50080
rect 185640 50080 185800 50240
rect 185640 50240 185800 50400
rect 185640 50400 185800 50560
rect 185640 50560 185800 50720
rect 185640 50720 185800 50880
rect 185640 50880 185800 51040
rect 185640 51040 185800 51200
rect 185640 51200 185800 51360
rect 185640 51360 185800 51520
rect 185640 51520 185800 51680
rect 185640 51680 185800 51840
rect 185640 51840 185800 52000
rect 185640 52000 185800 52160
rect 185640 52160 185800 52320
rect 185640 52320 185800 52480
rect 185640 52480 185800 52640
rect 185640 52640 185800 52800
rect 185800 40480 185960 40640
rect 185800 40640 185960 40800
rect 185800 40800 185960 40960
rect 185800 40960 185960 41120
rect 185800 41120 185960 41280
rect 185800 41280 185960 41440
rect 185800 41440 185960 41600
rect 185800 41600 185960 41760
rect 185800 41760 185960 41920
rect 185800 41920 185960 42080
rect 185800 42080 185960 42240
rect 185800 42240 185960 42400
rect 185800 42400 185960 42560
rect 185800 42560 185960 42720
rect 185800 42720 185960 42880
rect 185800 42880 185960 43040
rect 185800 43040 185960 43200
rect 185800 43200 185960 43360
rect 185800 43360 185960 43520
rect 185800 43520 185960 43680
rect 185800 43680 185960 43840
rect 185800 43840 185960 44000
rect 185800 44000 185960 44160
rect 185800 44160 185960 44320
rect 185800 44320 185960 44480
rect 185800 44480 185960 44640
rect 185800 44640 185960 44800
rect 185800 44800 185960 44960
rect 185800 44960 185960 45120
rect 185800 45120 185960 45280
rect 185800 45280 185960 45440
rect 185800 45440 185960 45600
rect 185800 45600 185960 45760
rect 185800 45760 185960 45920
rect 185800 45920 185960 46080
rect 185800 46080 185960 46240
rect 185800 46240 185960 46400
rect 185800 46400 185960 46560
rect 185800 46560 185960 46720
rect 185800 46720 185960 46880
rect 185800 46880 185960 47040
rect 185800 47040 185960 47200
rect 185800 47200 185960 47360
rect 185800 47360 185960 47520
rect 185800 47520 185960 47680
rect 185800 47680 185960 47840
rect 185800 47840 185960 48000
rect 185800 48000 185960 48160
rect 185800 48160 185960 48320
rect 185800 48320 185960 48480
rect 185800 48480 185960 48640
rect 185800 48640 185960 48800
rect 185800 48800 185960 48960
rect 185800 48960 185960 49120
rect 185800 49120 185960 49280
rect 185800 49280 185960 49440
rect 185800 49440 185960 49600
rect 185800 49600 185960 49760
rect 185800 49760 185960 49920
rect 185800 49920 185960 50080
rect 185800 50080 185960 50240
rect 185800 50240 185960 50400
rect 185800 50400 185960 50560
rect 185800 50560 185960 50720
rect 185800 50720 185960 50880
rect 185800 50880 185960 51040
rect 185800 51040 185960 51200
rect 185800 51200 185960 51360
rect 185800 51360 185960 51520
rect 185800 51520 185960 51680
rect 185800 51680 185960 51840
rect 185800 51840 185960 52000
rect 185800 52000 185960 52160
rect 185800 52160 185960 52320
rect 185800 52320 185960 52480
rect 185800 52480 185960 52640
rect 185800 52640 185960 52800
rect 185960 39680 186120 39840
rect 185960 39840 186120 40000
rect 185960 40000 186120 40160
rect 185960 40160 186120 40320
rect 185960 40320 186120 40480
rect 185960 40480 186120 40640
rect 185960 40640 186120 40800
rect 185960 40800 186120 40960
rect 185960 40960 186120 41120
rect 185960 41120 186120 41280
rect 185960 41280 186120 41440
rect 185960 41440 186120 41600
rect 185960 41600 186120 41760
rect 185960 41760 186120 41920
rect 185960 41920 186120 42080
rect 185960 42080 186120 42240
rect 185960 42240 186120 42400
rect 185960 42400 186120 42560
rect 185960 42560 186120 42720
rect 185960 42720 186120 42880
rect 185960 42880 186120 43040
rect 185960 43040 186120 43200
rect 185960 43200 186120 43360
rect 185960 43360 186120 43520
rect 185960 43520 186120 43680
rect 185960 43680 186120 43840
rect 185960 43840 186120 44000
rect 185960 44000 186120 44160
rect 185960 44160 186120 44320
rect 185960 44320 186120 44480
rect 185960 44480 186120 44640
rect 185960 44640 186120 44800
rect 185960 44800 186120 44960
rect 185960 44960 186120 45120
rect 185960 45120 186120 45280
rect 185960 45280 186120 45440
rect 185960 45440 186120 45600
rect 185960 45600 186120 45760
rect 185960 45760 186120 45920
rect 185960 45920 186120 46080
rect 185960 46080 186120 46240
rect 185960 46240 186120 46400
rect 185960 46400 186120 46560
rect 185960 46560 186120 46720
rect 185960 46720 186120 46880
rect 185960 46880 186120 47040
rect 185960 47040 186120 47200
rect 185960 47200 186120 47360
rect 185960 47360 186120 47520
rect 185960 47520 186120 47680
rect 185960 47680 186120 47840
rect 185960 47840 186120 48000
rect 185960 48000 186120 48160
rect 185960 48160 186120 48320
rect 185960 48320 186120 48480
rect 185960 48480 186120 48640
rect 185960 48640 186120 48800
rect 185960 48800 186120 48960
rect 185960 48960 186120 49120
rect 185960 49120 186120 49280
rect 185960 49280 186120 49440
rect 185960 49440 186120 49600
rect 185960 49600 186120 49760
rect 185960 49760 186120 49920
rect 185960 49920 186120 50080
rect 185960 50080 186120 50240
rect 185960 50240 186120 50400
rect 185960 50400 186120 50560
rect 185960 50560 186120 50720
rect 185960 50720 186120 50880
rect 185960 50880 186120 51040
rect 185960 51040 186120 51200
rect 185960 51200 186120 51360
rect 185960 51360 186120 51520
rect 185960 51520 186120 51680
rect 185960 51680 186120 51840
rect 185960 51840 186120 52000
rect 185960 52000 186120 52160
rect 185960 52160 186120 52320
rect 185960 52320 186120 52480
rect 185960 52480 186120 52640
rect 186120 38720 186280 38880
rect 186120 38880 186280 39040
rect 186120 39040 186280 39200
rect 186120 39200 186280 39360
rect 186120 39360 186280 39520
rect 186120 39520 186280 39680
rect 186120 39680 186280 39840
rect 186120 39840 186280 40000
rect 186120 40000 186280 40160
rect 186120 40160 186280 40320
rect 186120 40320 186280 40480
rect 186120 40480 186280 40640
rect 186120 40640 186280 40800
rect 186120 40800 186280 40960
rect 186120 40960 186280 41120
rect 186120 41120 186280 41280
rect 186120 41280 186280 41440
rect 186120 41440 186280 41600
rect 186120 41600 186280 41760
rect 186120 41760 186280 41920
rect 186120 41920 186280 42080
rect 186120 42080 186280 42240
rect 186120 42240 186280 42400
rect 186120 42400 186280 42560
rect 186120 42560 186280 42720
rect 186120 42720 186280 42880
rect 186120 42880 186280 43040
rect 186120 43040 186280 43200
rect 186120 43200 186280 43360
rect 186120 43360 186280 43520
rect 186120 43520 186280 43680
rect 186120 43680 186280 43840
rect 186120 43840 186280 44000
rect 186120 44000 186280 44160
rect 186120 44160 186280 44320
rect 186120 44320 186280 44480
rect 186120 44480 186280 44640
rect 186120 44640 186280 44800
rect 186120 44800 186280 44960
rect 186120 44960 186280 45120
rect 186120 45120 186280 45280
rect 186120 45280 186280 45440
rect 186120 45440 186280 45600
rect 186120 45600 186280 45760
rect 186120 45760 186280 45920
rect 186120 45920 186280 46080
rect 186120 46080 186280 46240
rect 186120 46240 186280 46400
rect 186120 46400 186280 46560
rect 186120 46560 186280 46720
rect 186120 46720 186280 46880
rect 186120 46880 186280 47040
rect 186120 47040 186280 47200
rect 186120 47200 186280 47360
rect 186120 47360 186280 47520
rect 186120 47520 186280 47680
rect 186120 47680 186280 47840
rect 186120 47840 186280 48000
rect 186120 48000 186280 48160
rect 186120 48160 186280 48320
rect 186120 48320 186280 48480
rect 186120 48480 186280 48640
rect 186120 48640 186280 48800
rect 186120 48800 186280 48960
rect 186120 48960 186280 49120
rect 186120 49120 186280 49280
rect 186120 49280 186280 49440
rect 186120 49440 186280 49600
rect 186120 49600 186280 49760
rect 186120 49760 186280 49920
rect 186120 49920 186280 50080
rect 186120 50080 186280 50240
rect 186120 50240 186280 50400
rect 186120 50400 186280 50560
rect 186120 50560 186280 50720
rect 186120 50720 186280 50880
rect 186120 50880 186280 51040
rect 186120 51040 186280 51200
rect 186120 51200 186280 51360
rect 186120 51360 186280 51520
rect 186120 51520 186280 51680
rect 186120 51680 186280 51840
rect 186120 51840 186280 52000
rect 186120 52000 186280 52160
rect 186120 52160 186280 52320
rect 186120 52320 186280 52480
rect 186120 52480 186280 52640
rect 186280 37920 186440 38080
rect 186280 38080 186440 38240
rect 186280 38240 186440 38400
rect 186280 38400 186440 38560
rect 186280 38560 186440 38720
rect 186280 38720 186440 38880
rect 186280 38880 186440 39040
rect 186280 39040 186440 39200
rect 186280 39200 186440 39360
rect 186280 39360 186440 39520
rect 186280 39520 186440 39680
rect 186280 39680 186440 39840
rect 186280 39840 186440 40000
rect 186280 40000 186440 40160
rect 186280 40160 186440 40320
rect 186280 40320 186440 40480
rect 186280 40480 186440 40640
rect 186280 40640 186440 40800
rect 186280 40800 186440 40960
rect 186280 40960 186440 41120
rect 186280 41120 186440 41280
rect 186280 41280 186440 41440
rect 186280 41440 186440 41600
rect 186280 41600 186440 41760
rect 186280 41760 186440 41920
rect 186280 41920 186440 42080
rect 186280 42080 186440 42240
rect 186280 42240 186440 42400
rect 186280 42400 186440 42560
rect 186280 42560 186440 42720
rect 186280 42720 186440 42880
rect 186280 42880 186440 43040
rect 186280 43040 186440 43200
rect 186280 43200 186440 43360
rect 186280 43360 186440 43520
rect 186280 43520 186440 43680
rect 186280 43680 186440 43840
rect 186280 43840 186440 44000
rect 186280 44000 186440 44160
rect 186280 44160 186440 44320
rect 186280 44320 186440 44480
rect 186280 44480 186440 44640
rect 186280 44640 186440 44800
rect 186280 44800 186440 44960
rect 186280 44960 186440 45120
rect 186280 45120 186440 45280
rect 186280 45280 186440 45440
rect 186280 45440 186440 45600
rect 186280 45600 186440 45760
rect 186280 45760 186440 45920
rect 186280 45920 186440 46080
rect 186280 46080 186440 46240
rect 186280 46240 186440 46400
rect 186280 46400 186440 46560
rect 186280 46560 186440 46720
rect 186280 46720 186440 46880
rect 186280 46880 186440 47040
rect 186280 47040 186440 47200
rect 186280 47200 186440 47360
rect 186280 47360 186440 47520
rect 186280 47520 186440 47680
rect 186280 47680 186440 47840
rect 186280 47840 186440 48000
rect 186280 48000 186440 48160
rect 186280 48160 186440 48320
rect 186280 48320 186440 48480
rect 186280 48480 186440 48640
rect 186280 48640 186440 48800
rect 186280 48800 186440 48960
rect 186280 48960 186440 49120
rect 186280 49120 186440 49280
rect 186280 49280 186440 49440
rect 186280 49440 186440 49600
rect 186280 49600 186440 49760
rect 186280 49760 186440 49920
rect 186280 49920 186440 50080
rect 186280 50080 186440 50240
rect 186280 50240 186440 50400
rect 186280 50400 186440 50560
rect 186280 50560 186440 50720
rect 186280 50720 186440 50880
rect 186280 50880 186440 51040
rect 186280 51040 186440 51200
rect 186280 51200 186440 51360
rect 186280 51360 186440 51520
rect 186280 51520 186440 51680
rect 186280 51680 186440 51840
rect 186280 51840 186440 52000
rect 186280 52000 186440 52160
rect 186280 52160 186440 52320
rect 186280 52320 186440 52480
rect 186280 52480 186440 52640
rect 186440 36960 186600 37120
rect 186440 37120 186600 37280
rect 186440 37280 186600 37440
rect 186440 37440 186600 37600
rect 186440 37600 186600 37760
rect 186440 37760 186600 37920
rect 186440 37920 186600 38080
rect 186440 38080 186600 38240
rect 186440 38240 186600 38400
rect 186440 38400 186600 38560
rect 186440 38560 186600 38720
rect 186440 38720 186600 38880
rect 186440 38880 186600 39040
rect 186440 39040 186600 39200
rect 186440 39200 186600 39360
rect 186440 39360 186600 39520
rect 186440 39520 186600 39680
rect 186440 39680 186600 39840
rect 186440 39840 186600 40000
rect 186440 40000 186600 40160
rect 186440 40160 186600 40320
rect 186440 40320 186600 40480
rect 186440 40480 186600 40640
rect 186440 40640 186600 40800
rect 186440 40800 186600 40960
rect 186440 40960 186600 41120
rect 186440 41120 186600 41280
rect 186440 41280 186600 41440
rect 186440 41440 186600 41600
rect 186440 41600 186600 41760
rect 186440 41760 186600 41920
rect 186440 41920 186600 42080
rect 186440 42080 186600 42240
rect 186440 42240 186600 42400
rect 186440 42400 186600 42560
rect 186440 42560 186600 42720
rect 186440 42720 186600 42880
rect 186440 42880 186600 43040
rect 186440 43040 186600 43200
rect 186440 43200 186600 43360
rect 186440 43360 186600 43520
rect 186440 43520 186600 43680
rect 186440 43680 186600 43840
rect 186440 43840 186600 44000
rect 186440 44000 186600 44160
rect 186440 44160 186600 44320
rect 186440 44320 186600 44480
rect 186440 44480 186600 44640
rect 186440 44640 186600 44800
rect 186440 44800 186600 44960
rect 186440 44960 186600 45120
rect 186440 45120 186600 45280
rect 186440 45280 186600 45440
rect 186440 45440 186600 45600
rect 186440 45600 186600 45760
rect 186440 45760 186600 45920
rect 186440 45920 186600 46080
rect 186440 46080 186600 46240
rect 186440 46240 186600 46400
rect 186440 46400 186600 46560
rect 186440 46560 186600 46720
rect 186440 46720 186600 46880
rect 186440 46880 186600 47040
rect 186440 47040 186600 47200
rect 186440 47200 186600 47360
rect 186440 47360 186600 47520
rect 186440 47520 186600 47680
rect 186440 47680 186600 47840
rect 186440 47840 186600 48000
rect 186440 48000 186600 48160
rect 186440 48160 186600 48320
rect 186440 48320 186600 48480
rect 186440 48480 186600 48640
rect 186440 48640 186600 48800
rect 186440 48800 186600 48960
rect 186440 48960 186600 49120
rect 186440 49120 186600 49280
rect 186440 49280 186600 49440
rect 186440 49440 186600 49600
rect 186440 49600 186600 49760
rect 186440 49760 186600 49920
rect 186440 49920 186600 50080
rect 186440 50080 186600 50240
rect 186440 50240 186600 50400
rect 186440 50400 186600 50560
rect 186440 50560 186600 50720
rect 186440 50720 186600 50880
rect 186440 50880 186600 51040
rect 186440 51040 186600 51200
rect 186440 51200 186600 51360
rect 186440 51360 186600 51520
rect 186440 51520 186600 51680
rect 186440 51680 186600 51840
rect 186440 51840 186600 52000
rect 186440 52000 186600 52160
rect 186440 52160 186600 52320
rect 186440 52320 186600 52480
rect 186600 36160 186760 36320
rect 186600 36320 186760 36480
rect 186600 36480 186760 36640
rect 186600 36640 186760 36800
rect 186600 36800 186760 36960
rect 186600 36960 186760 37120
rect 186600 37120 186760 37280
rect 186600 37280 186760 37440
rect 186600 37440 186760 37600
rect 186600 37600 186760 37760
rect 186600 37760 186760 37920
rect 186600 37920 186760 38080
rect 186600 38080 186760 38240
rect 186600 38240 186760 38400
rect 186600 38400 186760 38560
rect 186600 38560 186760 38720
rect 186600 38720 186760 38880
rect 186600 38880 186760 39040
rect 186600 39040 186760 39200
rect 186600 39200 186760 39360
rect 186600 39360 186760 39520
rect 186600 39520 186760 39680
rect 186600 39680 186760 39840
rect 186600 39840 186760 40000
rect 186600 40000 186760 40160
rect 186600 40160 186760 40320
rect 186600 40320 186760 40480
rect 186600 40480 186760 40640
rect 186600 40640 186760 40800
rect 186600 40800 186760 40960
rect 186600 40960 186760 41120
rect 186600 41120 186760 41280
rect 186600 41280 186760 41440
rect 186600 41440 186760 41600
rect 186600 41600 186760 41760
rect 186600 41760 186760 41920
rect 186600 41920 186760 42080
rect 186600 42080 186760 42240
rect 186600 42240 186760 42400
rect 186600 42400 186760 42560
rect 186600 42560 186760 42720
rect 186600 42720 186760 42880
rect 186600 42880 186760 43040
rect 186600 43040 186760 43200
rect 186600 43200 186760 43360
rect 186600 43360 186760 43520
rect 186600 43520 186760 43680
rect 186600 43680 186760 43840
rect 186600 43840 186760 44000
rect 186600 44000 186760 44160
rect 186600 44160 186760 44320
rect 186600 44320 186760 44480
rect 186600 44480 186760 44640
rect 186600 44640 186760 44800
rect 186600 44800 186760 44960
rect 186600 44960 186760 45120
rect 186600 45120 186760 45280
rect 186600 45280 186760 45440
rect 186600 45440 186760 45600
rect 186600 45600 186760 45760
rect 186600 45760 186760 45920
rect 186600 45920 186760 46080
rect 186600 46080 186760 46240
rect 186600 46240 186760 46400
rect 186600 46400 186760 46560
rect 186600 46560 186760 46720
rect 186600 46720 186760 46880
rect 186600 46880 186760 47040
rect 186600 47040 186760 47200
rect 186600 47200 186760 47360
rect 186600 47360 186760 47520
rect 186600 47520 186760 47680
rect 186600 47680 186760 47840
rect 186600 47840 186760 48000
rect 186600 48000 186760 48160
rect 186600 48160 186760 48320
rect 186600 48320 186760 48480
rect 186600 48480 186760 48640
rect 186600 48640 186760 48800
rect 186600 48800 186760 48960
rect 186600 48960 186760 49120
rect 186600 49120 186760 49280
rect 186600 49280 186760 49440
rect 186600 49440 186760 49600
rect 186600 49600 186760 49760
rect 186600 49760 186760 49920
rect 186600 49920 186760 50080
rect 186600 50080 186760 50240
rect 186600 50240 186760 50400
rect 186600 50400 186760 50560
rect 186600 50560 186760 50720
rect 186600 50720 186760 50880
rect 186600 50880 186760 51040
rect 186600 51040 186760 51200
rect 186600 51200 186760 51360
rect 186600 51360 186760 51520
rect 186600 51520 186760 51680
rect 186600 51680 186760 51840
rect 186600 51840 186760 52000
rect 186600 52000 186760 52160
rect 186600 52160 186760 52320
rect 186760 35360 186920 35520
rect 186760 35520 186920 35680
rect 186760 35680 186920 35840
rect 186760 35840 186920 36000
rect 186760 36000 186920 36160
rect 186760 36160 186920 36320
rect 186760 36320 186920 36480
rect 186760 36480 186920 36640
rect 186760 36640 186920 36800
rect 186760 36800 186920 36960
rect 186760 36960 186920 37120
rect 186760 37120 186920 37280
rect 186760 37280 186920 37440
rect 186760 37440 186920 37600
rect 186760 37600 186920 37760
rect 186760 37760 186920 37920
rect 186760 37920 186920 38080
rect 186760 38080 186920 38240
rect 186760 38240 186920 38400
rect 186760 38400 186920 38560
rect 186760 38560 186920 38720
rect 186760 38720 186920 38880
rect 186760 38880 186920 39040
rect 186760 39040 186920 39200
rect 186760 39200 186920 39360
rect 186760 39360 186920 39520
rect 186760 39520 186920 39680
rect 186760 39680 186920 39840
rect 186760 39840 186920 40000
rect 186760 40000 186920 40160
rect 186760 40160 186920 40320
rect 186760 40320 186920 40480
rect 186760 40480 186920 40640
rect 186760 40640 186920 40800
rect 186760 40800 186920 40960
rect 186760 40960 186920 41120
rect 186760 41120 186920 41280
rect 186760 41280 186920 41440
rect 186760 41440 186920 41600
rect 186760 41600 186920 41760
rect 186760 41760 186920 41920
rect 186760 41920 186920 42080
rect 186760 42080 186920 42240
rect 186760 42240 186920 42400
rect 186760 42400 186920 42560
rect 186760 42560 186920 42720
rect 186760 42720 186920 42880
rect 186760 42880 186920 43040
rect 186760 43040 186920 43200
rect 186760 43200 186920 43360
rect 186760 43360 186920 43520
rect 186760 43520 186920 43680
rect 186760 43680 186920 43840
rect 186760 43840 186920 44000
rect 186760 44000 186920 44160
rect 186760 44160 186920 44320
rect 186760 44320 186920 44480
rect 186760 44480 186920 44640
rect 186760 44640 186920 44800
rect 186760 44800 186920 44960
rect 186760 44960 186920 45120
rect 186760 45120 186920 45280
rect 186760 45280 186920 45440
rect 186760 45440 186920 45600
rect 186760 45600 186920 45760
rect 186760 45760 186920 45920
rect 186760 45920 186920 46080
rect 186760 46080 186920 46240
rect 186760 46240 186920 46400
rect 186760 46400 186920 46560
rect 186760 46560 186920 46720
rect 186760 46720 186920 46880
rect 186760 46880 186920 47040
rect 186760 47040 186920 47200
rect 186760 47200 186920 47360
rect 186760 47360 186920 47520
rect 186760 47520 186920 47680
rect 186760 47680 186920 47840
rect 186760 47840 186920 48000
rect 186760 48000 186920 48160
rect 186760 48160 186920 48320
rect 186760 48320 186920 48480
rect 186760 48480 186920 48640
rect 186760 48640 186920 48800
rect 186760 48800 186920 48960
rect 186760 48960 186920 49120
rect 186760 49120 186920 49280
rect 186760 49280 186920 49440
rect 186760 49440 186920 49600
rect 186760 49600 186920 49760
rect 186760 49760 186920 49920
rect 186760 49920 186920 50080
rect 186760 50080 186920 50240
rect 186760 50240 186920 50400
rect 186760 50400 186920 50560
rect 186760 50560 186920 50720
rect 186760 50720 186920 50880
rect 186760 50880 186920 51040
rect 186760 51040 186920 51200
rect 186760 51200 186920 51360
rect 186760 51360 186920 51520
rect 186760 51520 186920 51680
rect 186760 51680 186920 51840
rect 186760 51840 186920 52000
rect 186760 52000 186920 52160
rect 186920 34400 187080 34560
rect 186920 34560 187080 34720
rect 186920 34720 187080 34880
rect 186920 34880 187080 35040
rect 186920 35040 187080 35200
rect 186920 35200 187080 35360
rect 186920 35360 187080 35520
rect 186920 35520 187080 35680
rect 186920 35680 187080 35840
rect 186920 35840 187080 36000
rect 186920 36000 187080 36160
rect 186920 36160 187080 36320
rect 186920 36320 187080 36480
rect 186920 36480 187080 36640
rect 186920 36640 187080 36800
rect 186920 36800 187080 36960
rect 186920 36960 187080 37120
rect 186920 37120 187080 37280
rect 186920 37280 187080 37440
rect 186920 37440 187080 37600
rect 186920 37600 187080 37760
rect 186920 37760 187080 37920
rect 186920 37920 187080 38080
rect 186920 38080 187080 38240
rect 186920 38240 187080 38400
rect 186920 38400 187080 38560
rect 186920 38560 187080 38720
rect 186920 38720 187080 38880
rect 186920 38880 187080 39040
rect 186920 39040 187080 39200
rect 186920 39200 187080 39360
rect 186920 39360 187080 39520
rect 186920 39520 187080 39680
rect 186920 39680 187080 39840
rect 186920 39840 187080 40000
rect 186920 40000 187080 40160
rect 186920 40160 187080 40320
rect 186920 40320 187080 40480
rect 186920 40480 187080 40640
rect 186920 40640 187080 40800
rect 186920 40800 187080 40960
rect 186920 40960 187080 41120
rect 186920 41120 187080 41280
rect 186920 41280 187080 41440
rect 186920 41440 187080 41600
rect 186920 41600 187080 41760
rect 186920 41760 187080 41920
rect 186920 41920 187080 42080
rect 186920 42080 187080 42240
rect 186920 42240 187080 42400
rect 186920 42400 187080 42560
rect 186920 42560 187080 42720
rect 186920 42720 187080 42880
rect 186920 42880 187080 43040
rect 186920 43040 187080 43200
rect 186920 43200 187080 43360
rect 186920 43360 187080 43520
rect 186920 43520 187080 43680
rect 186920 43680 187080 43840
rect 186920 43840 187080 44000
rect 186920 44000 187080 44160
rect 186920 44160 187080 44320
rect 186920 44320 187080 44480
rect 186920 44480 187080 44640
rect 186920 44640 187080 44800
rect 186920 44800 187080 44960
rect 186920 44960 187080 45120
rect 186920 45120 187080 45280
rect 186920 45280 187080 45440
rect 186920 45440 187080 45600
rect 186920 45600 187080 45760
rect 186920 45760 187080 45920
rect 186920 45920 187080 46080
rect 186920 46080 187080 46240
rect 186920 46240 187080 46400
rect 186920 46400 187080 46560
rect 186920 46560 187080 46720
rect 186920 46720 187080 46880
rect 186920 46880 187080 47040
rect 186920 47040 187080 47200
rect 186920 47200 187080 47360
rect 186920 47360 187080 47520
rect 186920 47520 187080 47680
rect 186920 47680 187080 47840
rect 186920 47840 187080 48000
rect 186920 48000 187080 48160
rect 186920 48160 187080 48320
rect 186920 48320 187080 48480
rect 186920 48480 187080 48640
rect 186920 48640 187080 48800
rect 186920 48800 187080 48960
rect 186920 48960 187080 49120
rect 186920 49120 187080 49280
rect 186920 49280 187080 49440
rect 186920 49440 187080 49600
rect 186920 49600 187080 49760
rect 186920 49760 187080 49920
rect 186920 49920 187080 50080
rect 186920 50080 187080 50240
rect 186920 50240 187080 50400
rect 186920 50400 187080 50560
rect 186920 50560 187080 50720
rect 186920 50720 187080 50880
rect 186920 50880 187080 51040
rect 186920 51040 187080 51200
rect 186920 51200 187080 51360
rect 186920 51360 187080 51520
rect 186920 51520 187080 51680
rect 186920 51680 187080 51840
rect 186920 51840 187080 52000
rect 187080 33600 187240 33760
rect 187080 33760 187240 33920
rect 187080 33920 187240 34080
rect 187080 34080 187240 34240
rect 187080 34240 187240 34400
rect 187080 34400 187240 34560
rect 187080 34560 187240 34720
rect 187080 34720 187240 34880
rect 187080 34880 187240 35040
rect 187080 35040 187240 35200
rect 187080 35200 187240 35360
rect 187080 35360 187240 35520
rect 187080 35520 187240 35680
rect 187080 35680 187240 35840
rect 187080 35840 187240 36000
rect 187080 36000 187240 36160
rect 187080 36160 187240 36320
rect 187080 36320 187240 36480
rect 187080 36480 187240 36640
rect 187080 36640 187240 36800
rect 187080 36800 187240 36960
rect 187080 36960 187240 37120
rect 187080 37120 187240 37280
rect 187080 37280 187240 37440
rect 187080 37440 187240 37600
rect 187080 37600 187240 37760
rect 187080 37760 187240 37920
rect 187080 37920 187240 38080
rect 187080 38080 187240 38240
rect 187080 38240 187240 38400
rect 187080 38400 187240 38560
rect 187080 38560 187240 38720
rect 187080 38720 187240 38880
rect 187080 38880 187240 39040
rect 187080 39040 187240 39200
rect 187080 39200 187240 39360
rect 187080 39360 187240 39520
rect 187080 39520 187240 39680
rect 187080 39680 187240 39840
rect 187080 39840 187240 40000
rect 187080 40000 187240 40160
rect 187080 40160 187240 40320
rect 187080 40320 187240 40480
rect 187080 40480 187240 40640
rect 187080 40640 187240 40800
rect 187080 40800 187240 40960
rect 187080 40960 187240 41120
rect 187080 41120 187240 41280
rect 187080 41280 187240 41440
rect 187080 41440 187240 41600
rect 187080 41600 187240 41760
rect 187080 41760 187240 41920
rect 187080 41920 187240 42080
rect 187080 42080 187240 42240
rect 187080 42240 187240 42400
rect 187080 42400 187240 42560
rect 187080 42560 187240 42720
rect 187080 42720 187240 42880
rect 187080 42880 187240 43040
rect 187080 43040 187240 43200
rect 187080 43200 187240 43360
rect 187080 43360 187240 43520
rect 187080 43520 187240 43680
rect 187080 43680 187240 43840
rect 187080 43840 187240 44000
rect 187080 44000 187240 44160
rect 187080 44160 187240 44320
rect 187080 44320 187240 44480
rect 187080 44480 187240 44640
rect 187080 44640 187240 44800
rect 187080 44800 187240 44960
rect 187080 44960 187240 45120
rect 187080 45120 187240 45280
rect 187080 45280 187240 45440
rect 187080 45440 187240 45600
rect 187080 45600 187240 45760
rect 187080 45760 187240 45920
rect 187080 45920 187240 46080
rect 187080 46080 187240 46240
rect 187080 46240 187240 46400
rect 187080 46400 187240 46560
rect 187080 46560 187240 46720
rect 187080 46720 187240 46880
rect 187080 46880 187240 47040
rect 187080 47040 187240 47200
rect 187080 47200 187240 47360
rect 187080 47360 187240 47520
rect 187080 47520 187240 47680
rect 187080 47680 187240 47840
rect 187080 47840 187240 48000
rect 187080 48000 187240 48160
rect 187080 48160 187240 48320
rect 187080 48320 187240 48480
rect 187080 48480 187240 48640
rect 187080 48640 187240 48800
rect 187080 48800 187240 48960
rect 187080 48960 187240 49120
rect 187080 49120 187240 49280
rect 187080 49280 187240 49440
rect 187080 49440 187240 49600
rect 187080 49600 187240 49760
rect 187080 49760 187240 49920
rect 187080 49920 187240 50080
rect 187080 50080 187240 50240
rect 187080 50240 187240 50400
rect 187080 50400 187240 50560
rect 187080 50560 187240 50720
rect 187080 50720 187240 50880
rect 187080 50880 187240 51040
rect 187080 51040 187240 51200
rect 187080 51200 187240 51360
rect 187080 51360 187240 51520
rect 187080 51520 187240 51680
rect 187240 32640 187400 32800
rect 187240 32800 187400 32960
rect 187240 32960 187400 33120
rect 187240 33120 187400 33280
rect 187240 33280 187400 33440
rect 187240 33440 187400 33600
rect 187240 33600 187400 33760
rect 187240 33760 187400 33920
rect 187240 33920 187400 34080
rect 187240 34080 187400 34240
rect 187240 34240 187400 34400
rect 187240 34400 187400 34560
rect 187240 34560 187400 34720
rect 187240 34720 187400 34880
rect 187240 34880 187400 35040
rect 187240 35040 187400 35200
rect 187240 35200 187400 35360
rect 187240 35360 187400 35520
rect 187240 35520 187400 35680
rect 187240 35680 187400 35840
rect 187240 35840 187400 36000
rect 187240 36000 187400 36160
rect 187240 36160 187400 36320
rect 187240 36320 187400 36480
rect 187240 36480 187400 36640
rect 187240 36640 187400 36800
rect 187240 36800 187400 36960
rect 187240 36960 187400 37120
rect 187240 37120 187400 37280
rect 187240 37280 187400 37440
rect 187240 37440 187400 37600
rect 187240 37600 187400 37760
rect 187240 37760 187400 37920
rect 187240 37920 187400 38080
rect 187240 38080 187400 38240
rect 187240 38240 187400 38400
rect 187240 38400 187400 38560
rect 187240 38560 187400 38720
rect 187240 38720 187400 38880
rect 187240 38880 187400 39040
rect 187240 39040 187400 39200
rect 187240 39200 187400 39360
rect 187240 39360 187400 39520
rect 187240 39520 187400 39680
rect 187240 39680 187400 39840
rect 187240 39840 187400 40000
rect 187240 40000 187400 40160
rect 187240 40160 187400 40320
rect 187240 40320 187400 40480
rect 187240 40480 187400 40640
rect 187240 40640 187400 40800
rect 187240 40800 187400 40960
rect 187240 40960 187400 41120
rect 187240 41120 187400 41280
rect 187240 41280 187400 41440
rect 187240 41440 187400 41600
rect 187240 41600 187400 41760
rect 187240 41760 187400 41920
rect 187240 41920 187400 42080
rect 187240 42080 187400 42240
rect 187240 42240 187400 42400
rect 187240 42400 187400 42560
rect 187240 42560 187400 42720
rect 187240 42720 187400 42880
rect 187240 42880 187400 43040
rect 187240 43040 187400 43200
rect 187240 43200 187400 43360
rect 187240 43360 187400 43520
rect 187240 43520 187400 43680
rect 187240 43680 187400 43840
rect 187240 43840 187400 44000
rect 187240 44000 187400 44160
rect 187240 44160 187400 44320
rect 187240 44320 187400 44480
rect 187240 44480 187400 44640
rect 187240 44640 187400 44800
rect 187240 44800 187400 44960
rect 187240 44960 187400 45120
rect 187240 45120 187400 45280
rect 187240 45280 187400 45440
rect 187240 45440 187400 45600
rect 187240 45600 187400 45760
rect 187240 45760 187400 45920
rect 187240 45920 187400 46080
rect 187240 46080 187400 46240
rect 187240 46240 187400 46400
rect 187240 46400 187400 46560
rect 187240 46560 187400 46720
rect 187240 46720 187400 46880
rect 187240 46880 187400 47040
rect 187240 47040 187400 47200
rect 187240 47200 187400 47360
rect 187240 47360 187400 47520
rect 187240 47520 187400 47680
rect 187240 47680 187400 47840
rect 187240 47840 187400 48000
rect 187240 48000 187400 48160
rect 187240 48160 187400 48320
rect 187240 48320 187400 48480
rect 187240 48480 187400 48640
rect 187240 48640 187400 48800
rect 187240 48800 187400 48960
rect 187240 48960 187400 49120
rect 187240 49120 187400 49280
rect 187240 49280 187400 49440
rect 187240 49440 187400 49600
rect 187240 49600 187400 49760
rect 187240 49760 187400 49920
rect 187240 49920 187400 50080
rect 187240 50080 187400 50240
rect 187240 50240 187400 50400
rect 187240 50400 187400 50560
rect 187240 50560 187400 50720
rect 187240 50720 187400 50880
rect 187240 50880 187400 51040
rect 187240 51040 187400 51200
rect 187400 31840 187560 32000
rect 187400 32000 187560 32160
rect 187400 32160 187560 32320
rect 187400 32320 187560 32480
rect 187400 32480 187560 32640
rect 187400 32640 187560 32800
rect 187400 32800 187560 32960
rect 187400 32960 187560 33120
rect 187400 33120 187560 33280
rect 187400 33280 187560 33440
rect 187400 33440 187560 33600
rect 187400 33600 187560 33760
rect 187400 33760 187560 33920
rect 187400 33920 187560 34080
rect 187400 34080 187560 34240
rect 187400 34240 187560 34400
rect 187400 34400 187560 34560
rect 187400 34560 187560 34720
rect 187400 34720 187560 34880
rect 187400 34880 187560 35040
rect 187400 35040 187560 35200
rect 187400 35200 187560 35360
rect 187400 35360 187560 35520
rect 187400 35520 187560 35680
rect 187400 35680 187560 35840
rect 187400 35840 187560 36000
rect 187400 36000 187560 36160
rect 187400 36160 187560 36320
rect 187400 36320 187560 36480
rect 187400 36480 187560 36640
rect 187400 36640 187560 36800
rect 187400 36800 187560 36960
rect 187400 36960 187560 37120
rect 187400 37120 187560 37280
rect 187400 37280 187560 37440
rect 187400 37440 187560 37600
rect 187400 37600 187560 37760
rect 187400 37760 187560 37920
rect 187400 37920 187560 38080
rect 187400 38080 187560 38240
rect 187400 38240 187560 38400
rect 187400 38400 187560 38560
rect 187400 38560 187560 38720
rect 187400 38720 187560 38880
rect 187400 38880 187560 39040
rect 187400 39040 187560 39200
rect 187400 39200 187560 39360
rect 187400 39360 187560 39520
rect 187400 39520 187560 39680
rect 187400 39680 187560 39840
rect 187400 39840 187560 40000
rect 187400 40000 187560 40160
rect 187400 40160 187560 40320
rect 187400 40320 187560 40480
rect 187400 40480 187560 40640
rect 187400 40640 187560 40800
rect 187400 40800 187560 40960
rect 187400 40960 187560 41120
rect 187400 41120 187560 41280
rect 187400 41280 187560 41440
rect 187400 41440 187560 41600
rect 187400 41600 187560 41760
rect 187400 41760 187560 41920
rect 187400 41920 187560 42080
rect 187400 42080 187560 42240
rect 187400 42240 187560 42400
rect 187400 42400 187560 42560
rect 187400 42560 187560 42720
rect 187400 42720 187560 42880
rect 187400 42880 187560 43040
rect 187400 43040 187560 43200
rect 187400 43200 187560 43360
rect 187400 43360 187560 43520
rect 187400 43520 187560 43680
rect 187400 43680 187560 43840
rect 187400 43840 187560 44000
rect 187400 44000 187560 44160
rect 187400 44160 187560 44320
rect 187400 44320 187560 44480
rect 187400 44480 187560 44640
rect 187400 44640 187560 44800
rect 187400 44800 187560 44960
rect 187400 44960 187560 45120
rect 187400 45120 187560 45280
rect 187400 45280 187560 45440
rect 187400 45440 187560 45600
rect 187400 45600 187560 45760
rect 187400 45760 187560 45920
rect 187400 45920 187560 46080
rect 187400 46080 187560 46240
rect 187400 46240 187560 46400
rect 187400 46400 187560 46560
rect 187400 46560 187560 46720
rect 187400 46720 187560 46880
rect 187400 46880 187560 47040
rect 187400 47040 187560 47200
rect 187400 47200 187560 47360
rect 187400 47360 187560 47520
rect 187400 47520 187560 47680
rect 187400 47680 187560 47840
rect 187400 47840 187560 48000
rect 187400 48000 187560 48160
rect 187400 48160 187560 48320
rect 187400 48320 187560 48480
rect 187400 48480 187560 48640
rect 187400 48640 187560 48800
rect 187400 48800 187560 48960
rect 187400 48960 187560 49120
rect 187400 49120 187560 49280
rect 187400 49280 187560 49440
rect 187400 49440 187560 49600
rect 187400 49600 187560 49760
rect 187400 49760 187560 49920
rect 187400 49920 187560 50080
rect 187400 50080 187560 50240
rect 187400 50240 187560 50400
rect 187400 50400 187560 50560
rect 187400 50560 187560 50720
rect 187560 30880 187720 31040
rect 187560 31040 187720 31200
rect 187560 31200 187720 31360
rect 187560 31360 187720 31520
rect 187560 31520 187720 31680
rect 187560 31680 187720 31840
rect 187560 31840 187720 32000
rect 187560 32000 187720 32160
rect 187560 32160 187720 32320
rect 187560 32320 187720 32480
rect 187560 32480 187720 32640
rect 187560 32640 187720 32800
rect 187560 32800 187720 32960
rect 187560 32960 187720 33120
rect 187560 33120 187720 33280
rect 187560 33280 187720 33440
rect 187560 33440 187720 33600
rect 187560 33600 187720 33760
rect 187560 33760 187720 33920
rect 187560 33920 187720 34080
rect 187560 34080 187720 34240
rect 187560 34240 187720 34400
rect 187560 34400 187720 34560
rect 187560 34560 187720 34720
rect 187560 34720 187720 34880
rect 187560 34880 187720 35040
rect 187560 35040 187720 35200
rect 187560 35200 187720 35360
rect 187560 35360 187720 35520
rect 187560 35520 187720 35680
rect 187560 35680 187720 35840
rect 187560 35840 187720 36000
rect 187560 36000 187720 36160
rect 187560 36160 187720 36320
rect 187560 36320 187720 36480
rect 187560 36480 187720 36640
rect 187560 36640 187720 36800
rect 187560 36800 187720 36960
rect 187560 36960 187720 37120
rect 187560 37120 187720 37280
rect 187560 37280 187720 37440
rect 187560 37440 187720 37600
rect 187560 37600 187720 37760
rect 187560 37760 187720 37920
rect 187560 37920 187720 38080
rect 187560 38080 187720 38240
rect 187560 38240 187720 38400
rect 187560 38400 187720 38560
rect 187560 38560 187720 38720
rect 187560 38720 187720 38880
rect 187560 38880 187720 39040
rect 187560 39040 187720 39200
rect 187560 39200 187720 39360
rect 187560 39360 187720 39520
rect 187560 39520 187720 39680
rect 187560 39680 187720 39840
rect 187560 39840 187720 40000
rect 187560 40000 187720 40160
rect 187560 40160 187720 40320
rect 187560 40320 187720 40480
rect 187560 40480 187720 40640
rect 187560 40640 187720 40800
rect 187560 40800 187720 40960
rect 187560 40960 187720 41120
rect 187560 41120 187720 41280
rect 187560 41280 187720 41440
rect 187560 41440 187720 41600
rect 187560 41600 187720 41760
rect 187560 41760 187720 41920
rect 187560 41920 187720 42080
rect 187560 42080 187720 42240
rect 187560 42240 187720 42400
rect 187560 42400 187720 42560
rect 187560 42560 187720 42720
rect 187560 42720 187720 42880
rect 187560 42880 187720 43040
rect 187560 43040 187720 43200
rect 187560 43200 187720 43360
rect 187560 43360 187720 43520
rect 187560 43520 187720 43680
rect 187560 43680 187720 43840
rect 187560 43840 187720 44000
rect 187560 44000 187720 44160
rect 187560 44160 187720 44320
rect 187560 44320 187720 44480
rect 187560 44480 187720 44640
rect 187560 44640 187720 44800
rect 187560 44800 187720 44960
rect 187560 44960 187720 45120
rect 187560 45120 187720 45280
rect 187560 45280 187720 45440
rect 187560 45440 187720 45600
rect 187560 45600 187720 45760
rect 187560 45760 187720 45920
rect 187560 45920 187720 46080
rect 187560 46080 187720 46240
rect 187560 46240 187720 46400
rect 187560 46400 187720 46560
rect 187560 46560 187720 46720
rect 187560 46720 187720 46880
rect 187560 46880 187720 47040
rect 187560 47040 187720 47200
rect 187560 47200 187720 47360
rect 187560 47360 187720 47520
rect 187560 47520 187720 47680
rect 187560 47680 187720 47840
rect 187560 47840 187720 48000
rect 187560 48000 187720 48160
rect 187560 48160 187720 48320
rect 187560 48320 187720 48480
rect 187560 48480 187720 48640
rect 187560 48640 187720 48800
rect 187560 48800 187720 48960
rect 187560 48960 187720 49120
rect 187560 49120 187720 49280
rect 187560 49280 187720 49440
rect 187560 49440 187720 49600
rect 187560 49600 187720 49760
rect 187560 49760 187720 49920
rect 187720 30080 187880 30240
rect 187720 30240 187880 30400
rect 187720 30400 187880 30560
rect 187720 30560 187880 30720
rect 187720 30720 187880 30880
rect 187720 30880 187880 31040
rect 187720 31040 187880 31200
rect 187720 31200 187880 31360
rect 187720 31360 187880 31520
rect 187720 31520 187880 31680
rect 187720 31680 187880 31840
rect 187720 31840 187880 32000
rect 187720 32000 187880 32160
rect 187720 32160 187880 32320
rect 187720 32320 187880 32480
rect 187720 32480 187880 32640
rect 187720 32640 187880 32800
rect 187720 32800 187880 32960
rect 187720 32960 187880 33120
rect 187720 33120 187880 33280
rect 187720 33280 187880 33440
rect 187720 33440 187880 33600
rect 187720 33600 187880 33760
rect 187720 33760 187880 33920
rect 187720 33920 187880 34080
rect 187720 34080 187880 34240
rect 187720 34240 187880 34400
rect 187720 34400 187880 34560
rect 187720 34560 187880 34720
rect 187720 34720 187880 34880
rect 187720 34880 187880 35040
rect 187720 35040 187880 35200
rect 187720 35200 187880 35360
rect 187720 35360 187880 35520
rect 187720 35520 187880 35680
rect 187720 35680 187880 35840
rect 187720 35840 187880 36000
rect 187720 36000 187880 36160
rect 187720 36160 187880 36320
rect 187720 36320 187880 36480
rect 187720 36480 187880 36640
rect 187720 36640 187880 36800
rect 187720 36800 187880 36960
rect 187720 36960 187880 37120
rect 187720 37120 187880 37280
rect 187720 37280 187880 37440
rect 187720 37440 187880 37600
rect 187720 37600 187880 37760
rect 187720 37760 187880 37920
rect 187720 37920 187880 38080
rect 187720 38080 187880 38240
rect 187720 38240 187880 38400
rect 187720 38400 187880 38560
rect 187720 38560 187880 38720
rect 187720 38720 187880 38880
rect 187720 38880 187880 39040
rect 187720 39040 187880 39200
rect 187720 39200 187880 39360
rect 187720 39360 187880 39520
rect 187720 39520 187880 39680
rect 187720 39680 187880 39840
rect 187720 39840 187880 40000
rect 187720 40000 187880 40160
rect 187720 40160 187880 40320
rect 187720 40320 187880 40480
rect 187720 40480 187880 40640
rect 187720 40640 187880 40800
rect 187720 40800 187880 40960
rect 187720 40960 187880 41120
rect 187720 41120 187880 41280
rect 187720 41280 187880 41440
rect 187720 41440 187880 41600
rect 187720 41600 187880 41760
rect 187720 41760 187880 41920
rect 187720 41920 187880 42080
rect 187720 42080 187880 42240
rect 187720 42240 187880 42400
rect 187720 42400 187880 42560
rect 187720 42560 187880 42720
rect 187720 42720 187880 42880
rect 187720 42880 187880 43040
rect 187720 43040 187880 43200
rect 187720 43200 187880 43360
rect 187720 43360 187880 43520
rect 187720 43520 187880 43680
rect 187720 43680 187880 43840
rect 187720 43840 187880 44000
rect 187720 44000 187880 44160
rect 187720 44160 187880 44320
rect 187720 44320 187880 44480
rect 187720 44480 187880 44640
rect 187720 44640 187880 44800
rect 187720 44800 187880 44960
rect 187720 44960 187880 45120
rect 187720 45120 187880 45280
rect 187720 45280 187880 45440
rect 187720 45440 187880 45600
rect 187720 45600 187880 45760
rect 187720 45760 187880 45920
rect 187720 45920 187880 46080
rect 187720 46080 187880 46240
rect 187720 46240 187880 46400
rect 187720 46400 187880 46560
rect 187720 46560 187880 46720
rect 187720 46720 187880 46880
rect 187720 46880 187880 47040
rect 187720 47040 187880 47200
rect 187720 47200 187880 47360
rect 187720 47360 187880 47520
rect 187720 47520 187880 47680
rect 187720 47680 187880 47840
rect 187720 47840 187880 48000
rect 187720 48000 187880 48160
rect 187720 48160 187880 48320
rect 187720 48320 187880 48480
rect 187720 48480 187880 48640
rect 187720 48640 187880 48800
rect 187720 48800 187880 48960
rect 187720 48960 187880 49120
rect 187880 29600 188040 29760
rect 187880 29760 188040 29920
rect 187880 29920 188040 30080
rect 187880 30080 188040 30240
rect 187880 30240 188040 30400
rect 187880 30400 188040 30560
rect 187880 30560 188040 30720
rect 187880 30720 188040 30880
rect 187880 30880 188040 31040
rect 187880 31040 188040 31200
rect 187880 31200 188040 31360
rect 187880 31360 188040 31520
rect 187880 31520 188040 31680
rect 187880 31680 188040 31840
rect 187880 31840 188040 32000
rect 187880 32000 188040 32160
rect 187880 32160 188040 32320
rect 187880 32320 188040 32480
rect 187880 32480 188040 32640
rect 187880 32640 188040 32800
rect 187880 32800 188040 32960
rect 187880 32960 188040 33120
rect 187880 33120 188040 33280
rect 187880 33280 188040 33440
rect 187880 33440 188040 33600
rect 187880 33600 188040 33760
rect 187880 33760 188040 33920
rect 187880 33920 188040 34080
rect 187880 34080 188040 34240
rect 187880 34240 188040 34400
rect 187880 34400 188040 34560
rect 187880 34560 188040 34720
rect 187880 34720 188040 34880
rect 187880 34880 188040 35040
rect 187880 35040 188040 35200
rect 187880 35200 188040 35360
rect 187880 35360 188040 35520
rect 187880 35520 188040 35680
rect 187880 35680 188040 35840
rect 187880 35840 188040 36000
rect 187880 36000 188040 36160
rect 187880 36160 188040 36320
rect 187880 36320 188040 36480
rect 187880 36480 188040 36640
rect 187880 36640 188040 36800
rect 187880 36800 188040 36960
rect 187880 36960 188040 37120
rect 187880 37120 188040 37280
rect 187880 37280 188040 37440
rect 187880 37440 188040 37600
rect 187880 37600 188040 37760
rect 187880 37760 188040 37920
rect 187880 37920 188040 38080
rect 187880 38080 188040 38240
rect 187880 38240 188040 38400
rect 187880 38400 188040 38560
rect 187880 38560 188040 38720
rect 187880 38720 188040 38880
rect 187880 38880 188040 39040
rect 187880 39040 188040 39200
rect 187880 39200 188040 39360
rect 187880 39360 188040 39520
rect 187880 39520 188040 39680
rect 187880 39680 188040 39840
rect 187880 39840 188040 40000
rect 187880 40000 188040 40160
rect 187880 40160 188040 40320
rect 187880 40320 188040 40480
rect 187880 40480 188040 40640
rect 187880 40640 188040 40800
rect 187880 40800 188040 40960
rect 187880 40960 188040 41120
rect 187880 41120 188040 41280
rect 187880 41280 188040 41440
rect 187880 41440 188040 41600
rect 187880 41600 188040 41760
rect 187880 41760 188040 41920
rect 187880 41920 188040 42080
rect 187880 42080 188040 42240
rect 187880 42240 188040 42400
rect 187880 42400 188040 42560
rect 187880 42560 188040 42720
rect 187880 42720 188040 42880
rect 187880 42880 188040 43040
rect 187880 43040 188040 43200
rect 187880 43200 188040 43360
rect 187880 43360 188040 43520
rect 187880 43520 188040 43680
rect 187880 43680 188040 43840
rect 187880 43840 188040 44000
rect 187880 44000 188040 44160
rect 187880 44160 188040 44320
rect 187880 44320 188040 44480
rect 187880 44480 188040 44640
rect 187880 44640 188040 44800
rect 187880 44800 188040 44960
rect 187880 44960 188040 45120
rect 187880 45120 188040 45280
rect 187880 45280 188040 45440
rect 187880 45440 188040 45600
rect 187880 45600 188040 45760
rect 187880 45760 188040 45920
rect 187880 45920 188040 46080
rect 187880 46080 188040 46240
rect 187880 46240 188040 46400
rect 187880 46400 188040 46560
rect 187880 46560 188040 46720
rect 187880 46720 188040 46880
rect 187880 46880 188040 47040
rect 187880 47040 188040 47200
rect 187880 47200 188040 47360
rect 187880 47360 188040 47520
rect 187880 47520 188040 47680
rect 187880 47680 188040 47840
rect 187880 47840 188040 48000
rect 187880 48000 188040 48160
rect 188040 29120 188200 29280
rect 188040 29280 188200 29440
rect 188040 29440 188200 29600
rect 188040 29600 188200 29760
rect 188040 29760 188200 29920
rect 188040 29920 188200 30080
rect 188040 30080 188200 30240
rect 188040 30240 188200 30400
rect 188040 30400 188200 30560
rect 188040 30560 188200 30720
rect 188040 30720 188200 30880
rect 188040 30880 188200 31040
rect 188040 31040 188200 31200
rect 188040 31200 188200 31360
rect 188040 31360 188200 31520
rect 188040 31520 188200 31680
rect 188040 31680 188200 31840
rect 188040 31840 188200 32000
rect 188040 32000 188200 32160
rect 188040 32160 188200 32320
rect 188040 32320 188200 32480
rect 188040 32480 188200 32640
rect 188040 32640 188200 32800
rect 188040 32800 188200 32960
rect 188040 32960 188200 33120
rect 188040 33120 188200 33280
rect 188040 33280 188200 33440
rect 188040 33440 188200 33600
rect 188040 33600 188200 33760
rect 188040 33760 188200 33920
rect 188040 33920 188200 34080
rect 188040 34080 188200 34240
rect 188040 34240 188200 34400
rect 188040 34400 188200 34560
rect 188040 34560 188200 34720
rect 188040 34720 188200 34880
rect 188040 34880 188200 35040
rect 188040 35040 188200 35200
rect 188040 35200 188200 35360
rect 188040 35360 188200 35520
rect 188040 35520 188200 35680
rect 188040 35680 188200 35840
rect 188040 35840 188200 36000
rect 188040 36000 188200 36160
rect 188040 36160 188200 36320
rect 188040 36320 188200 36480
rect 188040 36480 188200 36640
rect 188040 36640 188200 36800
rect 188040 36800 188200 36960
rect 188040 36960 188200 37120
rect 188040 37120 188200 37280
rect 188040 37280 188200 37440
rect 188040 37440 188200 37600
rect 188040 37600 188200 37760
rect 188040 37760 188200 37920
rect 188040 37920 188200 38080
rect 188040 38080 188200 38240
rect 188040 38240 188200 38400
rect 188040 38400 188200 38560
rect 188040 38560 188200 38720
rect 188040 38720 188200 38880
rect 188040 38880 188200 39040
rect 188040 39040 188200 39200
rect 188040 39200 188200 39360
rect 188040 39360 188200 39520
rect 188040 39520 188200 39680
rect 188040 39680 188200 39840
rect 188040 39840 188200 40000
rect 188040 40000 188200 40160
rect 188040 40160 188200 40320
rect 188040 40320 188200 40480
rect 188040 40480 188200 40640
rect 188040 40640 188200 40800
rect 188040 40800 188200 40960
rect 188040 40960 188200 41120
rect 188040 41120 188200 41280
rect 188040 41280 188200 41440
rect 188040 41440 188200 41600
rect 188040 41600 188200 41760
rect 188040 41760 188200 41920
rect 188040 41920 188200 42080
rect 188040 42080 188200 42240
rect 188040 42240 188200 42400
rect 188040 42400 188200 42560
rect 188040 42560 188200 42720
rect 188040 42720 188200 42880
rect 188040 42880 188200 43040
rect 188040 43040 188200 43200
rect 188040 43200 188200 43360
rect 188040 43360 188200 43520
rect 188040 43520 188200 43680
rect 188040 43680 188200 43840
rect 188040 43840 188200 44000
rect 188040 44000 188200 44160
rect 188040 44160 188200 44320
rect 188040 44320 188200 44480
rect 188040 44480 188200 44640
rect 188040 44640 188200 44800
rect 188040 44800 188200 44960
rect 188040 44960 188200 45120
rect 188040 45120 188200 45280
rect 188040 45280 188200 45440
rect 188040 45440 188200 45600
rect 188040 45600 188200 45760
rect 188040 45760 188200 45920
rect 188040 45920 188200 46080
rect 188040 46080 188200 46240
rect 188040 46240 188200 46400
rect 188040 46400 188200 46560
rect 188040 46560 188200 46720
rect 188040 46720 188200 46880
rect 188040 46880 188200 47040
rect 188200 28640 188360 28800
rect 188200 28800 188360 28960
rect 188200 28960 188360 29120
rect 188200 29120 188360 29280
rect 188200 29280 188360 29440
rect 188200 29440 188360 29600
rect 188200 29600 188360 29760
rect 188200 29760 188360 29920
rect 188200 29920 188360 30080
rect 188200 30080 188360 30240
rect 188200 30240 188360 30400
rect 188200 30400 188360 30560
rect 188200 30560 188360 30720
rect 188200 30720 188360 30880
rect 188200 30880 188360 31040
rect 188200 31040 188360 31200
rect 188200 31200 188360 31360
rect 188200 31360 188360 31520
rect 188200 31520 188360 31680
rect 188200 31680 188360 31840
rect 188200 31840 188360 32000
rect 188200 32000 188360 32160
rect 188200 32160 188360 32320
rect 188200 32320 188360 32480
rect 188200 32480 188360 32640
rect 188200 32640 188360 32800
rect 188200 32800 188360 32960
rect 188200 32960 188360 33120
rect 188200 33120 188360 33280
rect 188200 33280 188360 33440
rect 188200 33440 188360 33600
rect 188200 33600 188360 33760
rect 188200 33760 188360 33920
rect 188200 33920 188360 34080
rect 188200 34080 188360 34240
rect 188200 34240 188360 34400
rect 188200 34400 188360 34560
rect 188200 34560 188360 34720
rect 188200 34720 188360 34880
rect 188200 34880 188360 35040
rect 188200 35040 188360 35200
rect 188200 35200 188360 35360
rect 188200 35360 188360 35520
rect 188200 35520 188360 35680
rect 188200 35680 188360 35840
rect 188200 35840 188360 36000
rect 188200 36000 188360 36160
rect 188200 36160 188360 36320
rect 188200 36320 188360 36480
rect 188200 36480 188360 36640
rect 188200 36640 188360 36800
rect 188200 36800 188360 36960
rect 188200 36960 188360 37120
rect 188200 37120 188360 37280
rect 188200 37280 188360 37440
rect 188200 37440 188360 37600
rect 188200 37600 188360 37760
rect 188200 37760 188360 37920
rect 188200 37920 188360 38080
rect 188200 38080 188360 38240
rect 188200 38240 188360 38400
rect 188200 38400 188360 38560
rect 188200 38560 188360 38720
rect 188200 38720 188360 38880
rect 188200 38880 188360 39040
rect 188200 39040 188360 39200
rect 188200 39200 188360 39360
rect 188200 39360 188360 39520
rect 188200 39520 188360 39680
rect 188200 39680 188360 39840
rect 188200 39840 188360 40000
rect 188200 40000 188360 40160
rect 188200 40160 188360 40320
rect 188200 40320 188360 40480
rect 188200 40480 188360 40640
rect 188200 40640 188360 40800
rect 188200 40800 188360 40960
rect 188200 40960 188360 41120
rect 188200 41120 188360 41280
rect 188200 41280 188360 41440
rect 188200 41440 188360 41600
rect 188200 41600 188360 41760
rect 188200 41760 188360 41920
rect 188200 41920 188360 42080
rect 188200 42080 188360 42240
rect 188200 42240 188360 42400
rect 188200 42400 188360 42560
rect 188200 42560 188360 42720
rect 188200 42720 188360 42880
rect 188200 42880 188360 43040
rect 188200 43040 188360 43200
rect 188200 43200 188360 43360
rect 188200 43360 188360 43520
rect 188200 43520 188360 43680
rect 188200 43680 188360 43840
rect 188200 43840 188360 44000
rect 188200 44000 188360 44160
rect 188200 44160 188360 44320
rect 188200 44320 188360 44480
rect 188200 44480 188360 44640
rect 188200 44640 188360 44800
rect 188200 44800 188360 44960
rect 188200 44960 188360 45120
rect 188200 45120 188360 45280
rect 188200 45280 188360 45440
rect 188200 45440 188360 45600
rect 188200 45600 188360 45760
rect 188360 28160 188520 28320
rect 188360 28320 188520 28480
rect 188360 28480 188520 28640
rect 188360 28640 188520 28800
rect 188360 28800 188520 28960
rect 188360 28960 188520 29120
rect 188360 29120 188520 29280
rect 188360 29280 188520 29440
rect 188360 29440 188520 29600
rect 188360 29600 188520 29760
rect 188360 29760 188520 29920
rect 188360 29920 188520 30080
rect 188360 30080 188520 30240
rect 188360 30240 188520 30400
rect 188360 30400 188520 30560
rect 188360 30560 188520 30720
rect 188360 30720 188520 30880
rect 188360 30880 188520 31040
rect 188360 31040 188520 31200
rect 188360 31200 188520 31360
rect 188360 31360 188520 31520
rect 188360 31520 188520 31680
rect 188360 31680 188520 31840
rect 188360 31840 188520 32000
rect 188360 32000 188520 32160
rect 188360 32160 188520 32320
rect 188360 32320 188520 32480
rect 188360 32480 188520 32640
rect 188360 32640 188520 32800
rect 188360 32800 188520 32960
rect 188360 32960 188520 33120
rect 188360 33120 188520 33280
rect 188360 33280 188520 33440
rect 188360 33440 188520 33600
rect 188360 33600 188520 33760
rect 188360 33760 188520 33920
rect 188360 33920 188520 34080
rect 188360 34080 188520 34240
rect 188360 34240 188520 34400
rect 188360 34400 188520 34560
rect 188360 34560 188520 34720
rect 188360 34720 188520 34880
rect 188360 34880 188520 35040
rect 188360 35040 188520 35200
rect 188360 35200 188520 35360
rect 188360 35360 188520 35520
rect 188360 35520 188520 35680
rect 188360 35680 188520 35840
rect 188360 35840 188520 36000
rect 188360 36000 188520 36160
rect 188360 36160 188520 36320
rect 188360 36320 188520 36480
rect 188360 36480 188520 36640
rect 188360 36640 188520 36800
rect 188360 36800 188520 36960
rect 188360 36960 188520 37120
rect 188360 37120 188520 37280
rect 188360 37280 188520 37440
rect 188360 37440 188520 37600
rect 188360 37600 188520 37760
rect 188360 37760 188520 37920
rect 188360 37920 188520 38080
rect 188360 38080 188520 38240
rect 188360 38240 188520 38400
rect 188360 38400 188520 38560
rect 188360 38560 188520 38720
rect 188360 38720 188520 38880
rect 188360 38880 188520 39040
rect 188360 39040 188520 39200
rect 188360 39200 188520 39360
rect 188360 39360 188520 39520
rect 188360 39520 188520 39680
rect 188360 39680 188520 39840
rect 188360 39840 188520 40000
rect 188360 40000 188520 40160
rect 188360 40160 188520 40320
rect 188360 40320 188520 40480
rect 188360 40480 188520 40640
rect 188360 40640 188520 40800
rect 188360 40800 188520 40960
rect 188360 40960 188520 41120
rect 188360 41120 188520 41280
rect 188360 41280 188520 41440
rect 188360 41440 188520 41600
rect 188360 41600 188520 41760
rect 188360 41760 188520 41920
rect 188360 41920 188520 42080
rect 188360 42080 188520 42240
rect 188360 42240 188520 42400
rect 188360 42400 188520 42560
rect 188360 42560 188520 42720
rect 188360 42720 188520 42880
rect 188360 42880 188520 43040
rect 188360 43040 188520 43200
rect 188360 43200 188520 43360
rect 188360 43360 188520 43520
rect 188360 43520 188520 43680
rect 188360 43680 188520 43840
rect 188360 43840 188520 44000
rect 188360 44000 188520 44160
rect 188360 44160 188520 44320
rect 188360 44320 188520 44480
rect 188520 27520 188680 27680
rect 188520 27680 188680 27840
rect 188520 27840 188680 28000
rect 188520 28000 188680 28160
rect 188520 28160 188680 28320
rect 188520 28320 188680 28480
rect 188520 28480 188680 28640
rect 188520 28640 188680 28800
rect 188520 28800 188680 28960
rect 188520 28960 188680 29120
rect 188520 29120 188680 29280
rect 188520 29280 188680 29440
rect 188520 29440 188680 29600
rect 188520 29600 188680 29760
rect 188520 29760 188680 29920
rect 188520 29920 188680 30080
rect 188520 30080 188680 30240
rect 188520 30240 188680 30400
rect 188520 30400 188680 30560
rect 188520 30560 188680 30720
rect 188520 30720 188680 30880
rect 188520 30880 188680 31040
rect 188520 31040 188680 31200
rect 188520 31200 188680 31360
rect 188520 31360 188680 31520
rect 188520 31520 188680 31680
rect 188520 31680 188680 31840
rect 188520 31840 188680 32000
rect 188520 32000 188680 32160
rect 188520 32160 188680 32320
rect 188520 32320 188680 32480
rect 188520 32480 188680 32640
rect 188520 32640 188680 32800
rect 188520 32800 188680 32960
rect 188520 32960 188680 33120
rect 188520 33120 188680 33280
rect 188520 33280 188680 33440
rect 188520 33440 188680 33600
rect 188520 33600 188680 33760
rect 188520 33760 188680 33920
rect 188520 33920 188680 34080
rect 188520 34080 188680 34240
rect 188520 34240 188680 34400
rect 188520 34400 188680 34560
rect 188520 34560 188680 34720
rect 188520 34720 188680 34880
rect 188520 34880 188680 35040
rect 188520 35040 188680 35200
rect 188520 35200 188680 35360
rect 188520 35360 188680 35520
rect 188520 35520 188680 35680
rect 188520 35680 188680 35840
rect 188520 35840 188680 36000
rect 188520 36000 188680 36160
rect 188520 36160 188680 36320
rect 188520 36320 188680 36480
rect 188520 36480 188680 36640
rect 188520 36640 188680 36800
rect 188520 36800 188680 36960
rect 188520 36960 188680 37120
rect 188520 37120 188680 37280
rect 188520 37280 188680 37440
rect 188520 37440 188680 37600
rect 188520 37600 188680 37760
rect 188520 37760 188680 37920
rect 188520 37920 188680 38080
rect 188520 38080 188680 38240
rect 188520 38240 188680 38400
rect 188520 38400 188680 38560
rect 188520 38560 188680 38720
rect 188520 38720 188680 38880
rect 188520 38880 188680 39040
rect 188520 39040 188680 39200
rect 188520 39200 188680 39360
rect 188520 39360 188680 39520
rect 188520 39520 188680 39680
rect 188520 39680 188680 39840
rect 188520 39840 188680 40000
rect 188520 40000 188680 40160
rect 188520 40160 188680 40320
rect 188520 40320 188680 40480
rect 188520 40480 188680 40640
rect 188520 40640 188680 40800
rect 188520 40800 188680 40960
rect 188520 40960 188680 41120
rect 188520 41120 188680 41280
rect 188520 41280 188680 41440
rect 188520 41440 188680 41600
rect 188520 41600 188680 41760
rect 188520 41760 188680 41920
rect 188520 41920 188680 42080
rect 188520 42080 188680 42240
rect 188520 42240 188680 42400
rect 188520 42400 188680 42560
rect 188520 42560 188680 42720
rect 188520 42720 188680 42880
rect 188520 42880 188680 43040
rect 188520 43040 188680 43200
rect 188520 43200 188680 43360
rect 188680 27040 188840 27200
rect 188680 27200 188840 27360
rect 188680 27360 188840 27520
rect 188680 27520 188840 27680
rect 188680 27680 188840 27840
rect 188680 27840 188840 28000
rect 188680 28000 188840 28160
rect 188680 28160 188840 28320
rect 188680 28320 188840 28480
rect 188680 28480 188840 28640
rect 188680 28640 188840 28800
rect 188680 28800 188840 28960
rect 188680 28960 188840 29120
rect 188680 29120 188840 29280
rect 188680 29280 188840 29440
rect 188680 29440 188840 29600
rect 188680 29600 188840 29760
rect 188680 29760 188840 29920
rect 188680 29920 188840 30080
rect 188680 30080 188840 30240
rect 188680 30240 188840 30400
rect 188680 30400 188840 30560
rect 188680 30560 188840 30720
rect 188680 30720 188840 30880
rect 188680 30880 188840 31040
rect 188680 31040 188840 31200
rect 188680 31200 188840 31360
rect 188680 31360 188840 31520
rect 188680 31520 188840 31680
rect 188680 31680 188840 31840
rect 188680 31840 188840 32000
rect 188680 32000 188840 32160
rect 188680 32160 188840 32320
rect 188680 32320 188840 32480
rect 188680 32480 188840 32640
rect 188680 32640 188840 32800
rect 188680 32800 188840 32960
rect 188680 32960 188840 33120
rect 188680 33120 188840 33280
rect 188680 33280 188840 33440
rect 188680 33440 188840 33600
rect 188680 33600 188840 33760
rect 188680 33760 188840 33920
rect 188680 33920 188840 34080
rect 188680 34080 188840 34240
rect 188680 34240 188840 34400
rect 188680 34400 188840 34560
rect 188680 34560 188840 34720
rect 188680 34720 188840 34880
rect 188680 34880 188840 35040
rect 188680 35040 188840 35200
rect 188680 35200 188840 35360
rect 188680 35360 188840 35520
rect 188680 35520 188840 35680
rect 188680 35680 188840 35840
rect 188680 35840 188840 36000
rect 188680 36000 188840 36160
rect 188680 36160 188840 36320
rect 188680 36320 188840 36480
rect 188680 36480 188840 36640
rect 188680 36640 188840 36800
rect 188680 36800 188840 36960
rect 188680 36960 188840 37120
rect 188680 37120 188840 37280
rect 188680 37280 188840 37440
rect 188680 37440 188840 37600
rect 188680 37600 188840 37760
rect 188680 37760 188840 37920
rect 188680 37920 188840 38080
rect 188680 38080 188840 38240
rect 188680 38240 188840 38400
rect 188680 38400 188840 38560
rect 188680 38560 188840 38720
rect 188680 38720 188840 38880
rect 188680 38880 188840 39040
rect 188680 39040 188840 39200
rect 188680 39200 188840 39360
rect 188680 39360 188840 39520
rect 188680 39520 188840 39680
rect 188680 39680 188840 39840
rect 188680 39840 188840 40000
rect 188680 40000 188840 40160
rect 188680 40160 188840 40320
rect 188680 40320 188840 40480
rect 188680 40480 188840 40640
rect 188680 40640 188840 40800
rect 188680 40800 188840 40960
rect 188680 40960 188840 41120
rect 188680 41120 188840 41280
rect 188680 41280 188840 41440
rect 188680 41440 188840 41600
rect 188680 41600 188840 41760
rect 188680 41760 188840 41920
rect 188680 41920 188840 42080
rect 188680 42080 188840 42240
rect 188680 42240 188840 42400
rect 188840 26880 189000 27040
rect 188840 27040 189000 27200
rect 188840 27200 189000 27360
rect 188840 27360 189000 27520
rect 188840 27520 189000 27680
rect 188840 27680 189000 27840
rect 188840 27840 189000 28000
rect 188840 28000 189000 28160
rect 188840 28160 189000 28320
rect 188840 28320 189000 28480
rect 188840 28480 189000 28640
rect 188840 28640 189000 28800
rect 188840 28800 189000 28960
rect 188840 28960 189000 29120
rect 188840 29120 189000 29280
rect 188840 29280 189000 29440
rect 188840 29440 189000 29600
rect 188840 29600 189000 29760
rect 188840 29760 189000 29920
rect 188840 29920 189000 30080
rect 188840 30080 189000 30240
rect 188840 30240 189000 30400
rect 188840 30400 189000 30560
rect 188840 30560 189000 30720
rect 188840 30720 189000 30880
rect 188840 30880 189000 31040
rect 188840 31040 189000 31200
rect 188840 31200 189000 31360
rect 188840 31360 189000 31520
rect 188840 31520 189000 31680
rect 188840 31680 189000 31840
rect 188840 31840 189000 32000
rect 188840 32000 189000 32160
rect 188840 32160 189000 32320
rect 188840 32320 189000 32480
rect 188840 32480 189000 32640
rect 188840 32640 189000 32800
rect 188840 32800 189000 32960
rect 188840 32960 189000 33120
rect 188840 33120 189000 33280
rect 188840 33280 189000 33440
rect 188840 33440 189000 33600
rect 188840 33600 189000 33760
rect 188840 33760 189000 33920
rect 188840 33920 189000 34080
rect 188840 34080 189000 34240
rect 188840 34240 189000 34400
rect 188840 34400 189000 34560
rect 188840 34560 189000 34720
rect 188840 34720 189000 34880
rect 188840 34880 189000 35040
rect 188840 35040 189000 35200
rect 188840 35200 189000 35360
rect 188840 35360 189000 35520
rect 188840 35520 189000 35680
rect 188840 35680 189000 35840
rect 188840 35840 189000 36000
rect 188840 36000 189000 36160
rect 188840 36160 189000 36320
rect 188840 36320 189000 36480
rect 188840 36480 189000 36640
rect 188840 36640 189000 36800
rect 188840 36800 189000 36960
rect 188840 36960 189000 37120
rect 188840 37120 189000 37280
rect 188840 37280 189000 37440
rect 188840 37440 189000 37600
rect 188840 37600 189000 37760
rect 188840 37760 189000 37920
rect 188840 37920 189000 38080
rect 188840 38080 189000 38240
rect 188840 38240 189000 38400
rect 188840 38400 189000 38560
rect 188840 38560 189000 38720
rect 188840 38720 189000 38880
rect 188840 38880 189000 39040
rect 188840 39040 189000 39200
rect 188840 39200 189000 39360
rect 188840 39360 189000 39520
rect 188840 39520 189000 39680
rect 188840 39680 189000 39840
rect 188840 39840 189000 40000
rect 188840 40000 189000 40160
rect 188840 40160 189000 40320
rect 188840 40320 189000 40480
rect 188840 40480 189000 40640
rect 188840 40640 189000 40800
rect 188840 40800 189000 40960
rect 188840 40960 189000 41120
rect 188840 41120 189000 41280
rect 188840 41280 189000 41440
rect 189000 26720 189160 26880
rect 189000 26880 189160 27040
rect 189000 27040 189160 27200
rect 189000 27200 189160 27360
rect 189000 27360 189160 27520
rect 189000 27520 189160 27680
rect 189000 27680 189160 27840
rect 189000 27840 189160 28000
rect 189000 28000 189160 28160
rect 189000 28160 189160 28320
rect 189000 28320 189160 28480
rect 189000 28480 189160 28640
rect 189000 28640 189160 28800
rect 189000 28800 189160 28960
rect 189000 28960 189160 29120
rect 189000 29120 189160 29280
rect 189000 29280 189160 29440
rect 189000 29440 189160 29600
rect 189000 29600 189160 29760
rect 189000 29760 189160 29920
rect 189000 29920 189160 30080
rect 189000 30080 189160 30240
rect 189000 30240 189160 30400
rect 189000 30400 189160 30560
rect 189000 30560 189160 30720
rect 189000 30720 189160 30880
rect 189000 30880 189160 31040
rect 189000 31040 189160 31200
rect 189000 31200 189160 31360
rect 189000 31360 189160 31520
rect 189000 31520 189160 31680
rect 189000 31680 189160 31840
rect 189000 31840 189160 32000
rect 189000 32000 189160 32160
rect 189000 32160 189160 32320
rect 189000 32320 189160 32480
rect 189000 32480 189160 32640
rect 189000 32640 189160 32800
rect 189000 32800 189160 32960
rect 189000 32960 189160 33120
rect 189000 33120 189160 33280
rect 189000 33280 189160 33440
rect 189000 33440 189160 33600
rect 189000 33600 189160 33760
rect 189000 33760 189160 33920
rect 189000 33920 189160 34080
rect 189000 34080 189160 34240
rect 189000 34240 189160 34400
rect 189000 34400 189160 34560
rect 189000 34560 189160 34720
rect 189000 34720 189160 34880
rect 189000 34880 189160 35040
rect 189000 35040 189160 35200
rect 189000 35200 189160 35360
rect 189000 35360 189160 35520
rect 189000 35520 189160 35680
rect 189000 35680 189160 35840
rect 189000 35840 189160 36000
rect 189000 36000 189160 36160
rect 189000 36160 189160 36320
rect 189000 36320 189160 36480
rect 189000 36480 189160 36640
rect 189000 36640 189160 36800
rect 189000 36800 189160 36960
rect 189000 36960 189160 37120
rect 189000 37120 189160 37280
rect 189000 37280 189160 37440
rect 189000 37440 189160 37600
rect 189000 37600 189160 37760
rect 189000 37760 189160 37920
rect 189000 37920 189160 38080
rect 189000 38080 189160 38240
rect 189000 38240 189160 38400
rect 189000 38400 189160 38560
rect 189000 38560 189160 38720
rect 189000 38720 189160 38880
rect 189000 38880 189160 39040
rect 189000 39040 189160 39200
rect 189000 39200 189160 39360
rect 189000 39360 189160 39520
rect 189000 39520 189160 39680
rect 189000 39680 189160 39840
rect 189000 39840 189160 40000
rect 189000 40000 189160 40160
rect 189000 40160 189160 40320
rect 189000 40320 189160 40480
rect 189160 26560 189320 26720
rect 189160 26720 189320 26880
rect 189160 26880 189320 27040
rect 189160 27040 189320 27200
rect 189160 27200 189320 27360
rect 189160 27360 189320 27520
rect 189160 27520 189320 27680
rect 189160 27680 189320 27840
rect 189160 27840 189320 28000
rect 189160 28000 189320 28160
rect 189160 28160 189320 28320
rect 189160 28320 189320 28480
rect 189160 28480 189320 28640
rect 189160 28640 189320 28800
rect 189160 28800 189320 28960
rect 189160 28960 189320 29120
rect 189160 29120 189320 29280
rect 189160 29280 189320 29440
rect 189160 29440 189320 29600
rect 189160 29600 189320 29760
rect 189160 29760 189320 29920
rect 189160 29920 189320 30080
rect 189160 30080 189320 30240
rect 189160 30240 189320 30400
rect 189160 30400 189320 30560
rect 189160 30560 189320 30720
rect 189160 30720 189320 30880
rect 189160 30880 189320 31040
rect 189160 31040 189320 31200
rect 189160 31200 189320 31360
rect 189160 31360 189320 31520
rect 189160 31520 189320 31680
rect 189160 31680 189320 31840
rect 189160 31840 189320 32000
rect 189160 32000 189320 32160
rect 189160 32160 189320 32320
rect 189160 32320 189320 32480
rect 189160 32480 189320 32640
rect 189160 32640 189320 32800
rect 189160 32800 189320 32960
rect 189160 32960 189320 33120
rect 189160 33120 189320 33280
rect 189160 33280 189320 33440
rect 189160 33440 189320 33600
rect 189160 33600 189320 33760
rect 189160 33760 189320 33920
rect 189160 33920 189320 34080
rect 189160 34080 189320 34240
rect 189160 34240 189320 34400
rect 189160 34400 189320 34560
rect 189160 34560 189320 34720
rect 189160 34720 189320 34880
rect 189160 34880 189320 35040
rect 189160 35040 189320 35200
rect 189160 35200 189320 35360
rect 189160 35360 189320 35520
rect 189160 35520 189320 35680
rect 189160 35680 189320 35840
rect 189160 35840 189320 36000
rect 189160 36000 189320 36160
rect 189160 36160 189320 36320
rect 189160 36320 189320 36480
rect 189160 36480 189320 36640
rect 189160 36640 189320 36800
rect 189160 36800 189320 36960
rect 189160 36960 189320 37120
rect 189160 37120 189320 37280
rect 189160 37280 189320 37440
rect 189160 37440 189320 37600
rect 189160 37600 189320 37760
rect 189160 37760 189320 37920
rect 189160 37920 189320 38080
rect 189160 38080 189320 38240
rect 189160 38240 189320 38400
rect 189160 38400 189320 38560
rect 189160 38560 189320 38720
rect 189160 38720 189320 38880
rect 189160 38880 189320 39040
rect 189160 39040 189320 39200
rect 189160 39200 189320 39360
rect 189160 39360 189320 39520
rect 189160 39520 189320 39680
rect 189320 26400 189480 26560
rect 189320 26560 189480 26720
rect 189320 26720 189480 26880
rect 189320 26880 189480 27040
rect 189320 27040 189480 27200
rect 189320 27200 189480 27360
rect 189320 27360 189480 27520
rect 189320 27520 189480 27680
rect 189320 27680 189480 27840
rect 189320 27840 189480 28000
rect 189320 28000 189480 28160
rect 189320 28160 189480 28320
rect 189320 28320 189480 28480
rect 189320 28480 189480 28640
rect 189320 28640 189480 28800
rect 189320 28800 189480 28960
rect 189320 28960 189480 29120
rect 189320 29120 189480 29280
rect 189320 29280 189480 29440
rect 189320 29440 189480 29600
rect 189320 29600 189480 29760
rect 189320 29760 189480 29920
rect 189320 29920 189480 30080
rect 189320 30080 189480 30240
rect 189320 30240 189480 30400
rect 189320 30400 189480 30560
rect 189320 30560 189480 30720
rect 189320 30720 189480 30880
rect 189320 30880 189480 31040
rect 189320 31040 189480 31200
rect 189320 31200 189480 31360
rect 189320 31360 189480 31520
rect 189320 31520 189480 31680
rect 189320 31680 189480 31840
rect 189320 31840 189480 32000
rect 189320 32000 189480 32160
rect 189320 32160 189480 32320
rect 189320 32320 189480 32480
rect 189320 32480 189480 32640
rect 189320 32640 189480 32800
rect 189320 32800 189480 32960
rect 189320 32960 189480 33120
rect 189320 33120 189480 33280
rect 189320 33280 189480 33440
rect 189320 33440 189480 33600
rect 189320 33600 189480 33760
rect 189320 33760 189480 33920
rect 189320 33920 189480 34080
rect 189320 34080 189480 34240
rect 189320 34240 189480 34400
rect 189320 34400 189480 34560
rect 189320 34560 189480 34720
rect 189320 34720 189480 34880
rect 189320 34880 189480 35040
rect 189320 35040 189480 35200
rect 189320 35200 189480 35360
rect 189320 35360 189480 35520
rect 189320 35520 189480 35680
rect 189320 35680 189480 35840
rect 189320 35840 189480 36000
rect 189320 36000 189480 36160
rect 189320 36160 189480 36320
rect 189320 36320 189480 36480
rect 189320 36480 189480 36640
rect 189320 36640 189480 36800
rect 189320 36800 189480 36960
rect 189320 36960 189480 37120
rect 189320 37120 189480 37280
rect 189320 37280 189480 37440
rect 189320 37440 189480 37600
rect 189320 37600 189480 37760
rect 189320 37760 189480 37920
rect 189320 37920 189480 38080
rect 189320 38080 189480 38240
rect 189320 38240 189480 38400
rect 189320 38400 189480 38560
rect 189320 38560 189480 38720
rect 189320 38720 189480 38880
rect 189480 26240 189640 26400
rect 189480 26400 189640 26560
rect 189480 26560 189640 26720
rect 189480 26720 189640 26880
rect 189480 26880 189640 27040
rect 189480 27040 189640 27200
rect 189480 27200 189640 27360
rect 189480 27360 189640 27520
rect 189480 27520 189640 27680
rect 189480 27680 189640 27840
rect 189480 27840 189640 28000
rect 189480 28000 189640 28160
rect 189480 28160 189640 28320
rect 189480 28320 189640 28480
rect 189480 28480 189640 28640
rect 189480 28640 189640 28800
rect 189480 28800 189640 28960
rect 189480 28960 189640 29120
rect 189480 29120 189640 29280
rect 189480 29280 189640 29440
rect 189480 29440 189640 29600
rect 189480 29600 189640 29760
rect 189480 29760 189640 29920
rect 189480 29920 189640 30080
rect 189480 30080 189640 30240
rect 189480 30240 189640 30400
rect 189480 30400 189640 30560
rect 189480 30560 189640 30720
rect 189480 30720 189640 30880
rect 189480 30880 189640 31040
rect 189480 31040 189640 31200
rect 189480 31200 189640 31360
rect 189480 31360 189640 31520
rect 189480 31520 189640 31680
rect 189480 31680 189640 31840
rect 189480 31840 189640 32000
rect 189480 32000 189640 32160
rect 189480 32160 189640 32320
rect 189480 32320 189640 32480
rect 189480 32480 189640 32640
rect 189480 32640 189640 32800
rect 189480 32800 189640 32960
rect 189480 32960 189640 33120
rect 189480 33120 189640 33280
rect 189480 33280 189640 33440
rect 189480 33440 189640 33600
rect 189480 33600 189640 33760
rect 189480 33760 189640 33920
rect 189480 33920 189640 34080
rect 189480 34080 189640 34240
rect 189480 34240 189640 34400
rect 189480 34400 189640 34560
rect 189480 34560 189640 34720
rect 189480 34720 189640 34880
rect 189480 34880 189640 35040
rect 189480 35040 189640 35200
rect 189480 35200 189640 35360
rect 189480 35360 189640 35520
rect 189480 35520 189640 35680
rect 189480 35680 189640 35840
rect 189480 35840 189640 36000
rect 189480 36000 189640 36160
rect 189480 36160 189640 36320
rect 189480 36320 189640 36480
rect 189480 36480 189640 36640
rect 189480 36640 189640 36800
rect 189480 36800 189640 36960
rect 189480 36960 189640 37120
rect 189480 37120 189640 37280
rect 189480 37280 189640 37440
rect 189480 37440 189640 37600
rect 189480 37600 189640 37760
rect 189480 37760 189640 37920
rect 189480 37920 189640 38080
rect 189640 26240 189800 26400
rect 189640 26400 189800 26560
rect 189640 26560 189800 26720
rect 189640 26720 189800 26880
rect 189640 26880 189800 27040
rect 189640 27040 189800 27200
rect 189640 27200 189800 27360
rect 189640 27360 189800 27520
rect 189640 27520 189800 27680
rect 189640 27680 189800 27840
rect 189640 27840 189800 28000
rect 189640 28000 189800 28160
rect 189640 28160 189800 28320
rect 189640 28320 189800 28480
rect 189640 28480 189800 28640
rect 189640 28640 189800 28800
rect 189640 28800 189800 28960
rect 189640 28960 189800 29120
rect 189640 29120 189800 29280
rect 189640 29280 189800 29440
rect 189640 29440 189800 29600
rect 189640 29600 189800 29760
rect 189640 29760 189800 29920
rect 189640 29920 189800 30080
rect 189640 30080 189800 30240
rect 189640 30240 189800 30400
rect 189640 30400 189800 30560
rect 189640 30560 189800 30720
rect 189640 30720 189800 30880
rect 189640 30880 189800 31040
rect 189640 31040 189800 31200
rect 189640 31200 189800 31360
rect 189640 31360 189800 31520
rect 189640 31520 189800 31680
rect 189640 31680 189800 31840
rect 189640 31840 189800 32000
rect 189640 32000 189800 32160
rect 189640 32160 189800 32320
rect 189640 32320 189800 32480
rect 189640 32480 189800 32640
rect 189640 32640 189800 32800
rect 189640 32800 189800 32960
rect 189640 32960 189800 33120
rect 189640 33120 189800 33280
rect 189640 33280 189800 33440
rect 189640 33440 189800 33600
rect 189640 33600 189800 33760
rect 189640 33760 189800 33920
rect 189640 33920 189800 34080
rect 189640 34080 189800 34240
rect 189640 34240 189800 34400
rect 189640 34400 189800 34560
rect 189640 34560 189800 34720
rect 189640 34720 189800 34880
rect 189640 34880 189800 35040
rect 189640 35040 189800 35200
rect 189640 35200 189800 35360
rect 189640 35360 189800 35520
rect 189640 35520 189800 35680
rect 189640 35680 189800 35840
rect 189640 35840 189800 36000
rect 189640 36000 189800 36160
rect 189640 36160 189800 36320
rect 189640 36320 189800 36480
rect 189640 36480 189800 36640
rect 189640 36640 189800 36800
rect 189640 36800 189800 36960
rect 189640 36960 189800 37120
rect 189640 37120 189800 37280
rect 189800 26240 189960 26400
rect 189800 26400 189960 26560
rect 189800 26560 189960 26720
rect 189800 26720 189960 26880
rect 189800 26880 189960 27040
rect 189800 27040 189960 27200
rect 189800 27200 189960 27360
rect 189800 27360 189960 27520
rect 189800 27520 189960 27680
rect 189800 27680 189960 27840
rect 189800 27840 189960 28000
rect 189800 28000 189960 28160
rect 189800 28160 189960 28320
rect 189800 28320 189960 28480
rect 189800 28480 189960 28640
rect 189800 28640 189960 28800
rect 189800 28800 189960 28960
rect 189800 28960 189960 29120
rect 189800 29120 189960 29280
rect 189800 29280 189960 29440
rect 189800 29440 189960 29600
rect 189800 29600 189960 29760
rect 189800 29760 189960 29920
rect 189800 29920 189960 30080
rect 189800 30080 189960 30240
rect 189800 30240 189960 30400
rect 189800 30400 189960 30560
rect 189800 30560 189960 30720
rect 189800 30720 189960 30880
rect 189800 30880 189960 31040
rect 189800 31040 189960 31200
rect 189800 31200 189960 31360
rect 189800 31360 189960 31520
rect 189800 31520 189960 31680
rect 189800 31680 189960 31840
rect 189800 31840 189960 32000
rect 189800 32000 189960 32160
rect 189800 32160 189960 32320
rect 189800 32320 189960 32480
rect 189800 32480 189960 32640
rect 189800 32640 189960 32800
rect 189800 32800 189960 32960
rect 189800 32960 189960 33120
rect 189800 33120 189960 33280
rect 189800 33280 189960 33440
rect 189800 33440 189960 33600
rect 189800 33600 189960 33760
rect 189800 33760 189960 33920
rect 189800 33920 189960 34080
rect 189800 34080 189960 34240
rect 189800 34240 189960 34400
rect 189800 34400 189960 34560
rect 189800 34560 189960 34720
rect 189800 34720 189960 34880
rect 189800 34880 189960 35040
rect 189800 35040 189960 35200
rect 189800 35200 189960 35360
rect 189800 35360 189960 35520
rect 189800 35520 189960 35680
rect 189800 35680 189960 35840
rect 189800 35840 189960 36000
rect 189800 36000 189960 36160
rect 189800 36160 189960 36320
rect 189800 36320 189960 36480
rect 189800 36480 189960 36640
rect 189960 26080 190120 26240
rect 189960 26240 190120 26400
rect 189960 26400 190120 26560
rect 189960 26560 190120 26720
rect 189960 26720 190120 26880
rect 189960 26880 190120 27040
rect 189960 27040 190120 27200
rect 189960 27200 190120 27360
rect 189960 27360 190120 27520
rect 189960 27520 190120 27680
rect 189960 27680 190120 27840
rect 189960 27840 190120 28000
rect 189960 28000 190120 28160
rect 189960 28160 190120 28320
rect 189960 28320 190120 28480
rect 189960 28480 190120 28640
rect 189960 28640 190120 28800
rect 189960 28800 190120 28960
rect 189960 28960 190120 29120
rect 189960 29120 190120 29280
rect 189960 29280 190120 29440
rect 189960 29440 190120 29600
rect 189960 29600 190120 29760
rect 189960 29760 190120 29920
rect 189960 29920 190120 30080
rect 189960 30080 190120 30240
rect 189960 30240 190120 30400
rect 189960 30400 190120 30560
rect 189960 30560 190120 30720
rect 189960 30720 190120 30880
rect 189960 30880 190120 31040
rect 189960 31040 190120 31200
rect 189960 31200 190120 31360
rect 189960 31360 190120 31520
rect 189960 31520 190120 31680
rect 189960 31680 190120 31840
rect 189960 31840 190120 32000
rect 189960 32000 190120 32160
rect 189960 32160 190120 32320
rect 189960 32320 190120 32480
rect 189960 32480 190120 32640
rect 189960 32640 190120 32800
rect 189960 32800 190120 32960
rect 189960 32960 190120 33120
rect 189960 33120 190120 33280
rect 189960 33280 190120 33440
rect 189960 33440 190120 33600
rect 189960 33600 190120 33760
rect 189960 33760 190120 33920
rect 189960 33920 190120 34080
rect 189960 34080 190120 34240
rect 189960 34240 190120 34400
rect 189960 34400 190120 34560
rect 189960 34560 190120 34720
rect 189960 34720 190120 34880
rect 189960 34880 190120 35040
rect 189960 35040 190120 35200
rect 189960 35200 190120 35360
rect 189960 35360 190120 35520
rect 189960 35520 190120 35680
rect 189960 35680 190120 35840
rect 190120 26080 190280 26240
rect 190120 26240 190280 26400
rect 190120 26400 190280 26560
rect 190120 26560 190280 26720
rect 190120 26720 190280 26880
rect 190120 26880 190280 27040
rect 190120 27040 190280 27200
rect 190120 27200 190280 27360
rect 190120 27360 190280 27520
rect 190120 27520 190280 27680
rect 190120 27680 190280 27840
rect 190120 27840 190280 28000
rect 190120 28000 190280 28160
rect 190120 28160 190280 28320
rect 190120 28320 190280 28480
rect 190120 28480 190280 28640
rect 190120 28640 190280 28800
rect 190120 28800 190280 28960
rect 190120 28960 190280 29120
rect 190120 29120 190280 29280
rect 190120 29280 190280 29440
rect 190120 29440 190280 29600
rect 190120 29600 190280 29760
rect 190120 29760 190280 29920
rect 190120 29920 190280 30080
rect 190120 30080 190280 30240
rect 190120 30240 190280 30400
rect 190120 30400 190280 30560
rect 190120 30560 190280 30720
rect 190120 30720 190280 30880
rect 190120 30880 190280 31040
rect 190120 31040 190280 31200
rect 190120 31200 190280 31360
rect 190120 31360 190280 31520
rect 190120 31520 190280 31680
rect 190120 31680 190280 31840
rect 190120 31840 190280 32000
rect 190120 32000 190280 32160
rect 190120 32160 190280 32320
rect 190120 32320 190280 32480
rect 190120 32480 190280 32640
rect 190120 32640 190280 32800
rect 190120 32800 190280 32960
rect 190120 32960 190280 33120
rect 190120 33120 190280 33280
rect 190120 33280 190280 33440
rect 190120 33440 190280 33600
rect 190120 33600 190280 33760
rect 190120 33760 190280 33920
rect 190120 33920 190280 34080
rect 190120 34080 190280 34240
rect 190120 34240 190280 34400
rect 190120 34400 190280 34560
rect 190120 34560 190280 34720
rect 190120 34720 190280 34880
rect 190120 34880 190280 35040
rect 190120 35040 190280 35200
rect 190280 26080 190440 26240
rect 190280 26240 190440 26400
rect 190280 26400 190440 26560
rect 190280 26560 190440 26720
rect 190280 26720 190440 26880
rect 190280 26880 190440 27040
rect 190280 27040 190440 27200
rect 190280 27200 190440 27360
rect 190280 27360 190440 27520
rect 190280 27520 190440 27680
rect 190280 27680 190440 27840
rect 190280 27840 190440 28000
rect 190280 28000 190440 28160
rect 190280 28160 190440 28320
rect 190280 28320 190440 28480
rect 190280 28480 190440 28640
rect 190280 28640 190440 28800
rect 190280 28800 190440 28960
rect 190280 28960 190440 29120
rect 190280 29120 190440 29280
rect 190280 29280 190440 29440
rect 190280 29440 190440 29600
rect 190280 29600 190440 29760
rect 190280 29760 190440 29920
rect 190280 29920 190440 30080
rect 190280 30080 190440 30240
rect 190280 30240 190440 30400
rect 190280 30400 190440 30560
rect 190280 30560 190440 30720
rect 190280 30720 190440 30880
rect 190280 30880 190440 31040
rect 190280 31040 190440 31200
rect 190280 31200 190440 31360
rect 190280 31360 190440 31520
rect 190280 31520 190440 31680
rect 190280 31680 190440 31840
rect 190280 31840 190440 32000
rect 190280 32000 190440 32160
rect 190280 32160 190440 32320
rect 190280 32320 190440 32480
rect 190280 32480 190440 32640
rect 190280 32640 190440 32800
rect 190280 32800 190440 32960
rect 190280 32960 190440 33120
rect 190280 33120 190440 33280
rect 190280 33280 190440 33440
rect 190280 33440 190440 33600
rect 190280 33600 190440 33760
rect 190280 33760 190440 33920
rect 190280 33920 190440 34080
rect 190280 34080 190440 34240
rect 190280 34240 190440 34400
rect 190440 26080 190600 26240
rect 190440 26240 190600 26400
rect 190440 26400 190600 26560
rect 190440 26560 190600 26720
rect 190440 26720 190600 26880
rect 190440 26880 190600 27040
rect 190440 27040 190600 27200
rect 190440 27200 190600 27360
rect 190440 27360 190600 27520
rect 190440 27520 190600 27680
rect 190440 27680 190600 27840
rect 190440 27840 190600 28000
rect 190440 28000 190600 28160
rect 190440 28160 190600 28320
rect 190440 28320 190600 28480
rect 190440 28480 190600 28640
rect 190440 28640 190600 28800
rect 190440 28800 190600 28960
rect 190440 28960 190600 29120
rect 190440 29120 190600 29280
rect 190440 29280 190600 29440
rect 190440 29440 190600 29600
rect 190440 29600 190600 29760
rect 190440 29760 190600 29920
rect 190440 29920 190600 30080
rect 190440 30080 190600 30240
rect 190440 30240 190600 30400
rect 190440 30400 190600 30560
rect 190440 30560 190600 30720
rect 190440 30720 190600 30880
rect 190440 30880 190600 31040
rect 190440 31040 190600 31200
rect 190440 31200 190600 31360
rect 190440 31360 190600 31520
rect 190440 31520 190600 31680
rect 190440 31680 190600 31840
rect 190440 31840 190600 32000
rect 190440 32000 190600 32160
rect 190440 32160 190600 32320
rect 190440 32320 190600 32480
rect 190440 32480 190600 32640
rect 190440 32640 190600 32800
rect 190440 32800 190600 32960
rect 190440 32960 190600 33120
rect 190440 33120 190600 33280
rect 190440 33280 190600 33440
rect 190440 33440 190600 33600
rect 190440 33600 190600 33760
rect 190600 26080 190760 26240
rect 190600 26240 190760 26400
rect 190600 26400 190760 26560
rect 190600 26560 190760 26720
rect 190600 26720 190760 26880
rect 190600 26880 190760 27040
rect 190600 27040 190760 27200
rect 190600 27200 190760 27360
rect 190600 27360 190760 27520
rect 190600 27520 190760 27680
rect 190600 27680 190760 27840
rect 190600 27840 190760 28000
rect 190600 28000 190760 28160
rect 190600 28160 190760 28320
rect 190600 28320 190760 28480
rect 190600 28480 190760 28640
rect 190600 28640 190760 28800
rect 190600 28800 190760 28960
rect 190600 28960 190760 29120
rect 190600 29120 190760 29280
rect 190600 29280 190760 29440
rect 190600 29440 190760 29600
rect 190600 29600 190760 29760
rect 190600 29760 190760 29920
rect 190600 29920 190760 30080
rect 190600 30080 190760 30240
rect 190600 30240 190760 30400
rect 190600 30400 190760 30560
rect 190600 30560 190760 30720
rect 190600 30720 190760 30880
rect 190600 30880 190760 31040
rect 190600 31040 190760 31200
rect 190600 31200 190760 31360
rect 190600 31360 190760 31520
rect 190600 31520 190760 31680
rect 190600 31680 190760 31840
rect 190600 31840 190760 32000
rect 190600 32000 190760 32160
rect 190600 32160 190760 32320
rect 190600 32320 190760 32480
rect 190600 32480 190760 32640
rect 190600 32640 190760 32800
rect 190600 32800 190760 32960
rect 190760 26080 190920 26240
rect 190760 26240 190920 26400
rect 190760 26400 190920 26560
rect 190760 26560 190920 26720
rect 190760 26720 190920 26880
rect 190760 26880 190920 27040
rect 190760 27040 190920 27200
rect 190760 27200 190920 27360
rect 190760 27360 190920 27520
rect 190760 27520 190920 27680
rect 190760 27680 190920 27840
rect 190760 27840 190920 28000
rect 190760 28000 190920 28160
rect 190760 28160 190920 28320
rect 190760 28320 190920 28480
rect 190760 28480 190920 28640
rect 190760 28640 190920 28800
rect 190760 28800 190920 28960
rect 190760 28960 190920 29120
rect 190760 29120 190920 29280
rect 190760 29280 190920 29440
rect 190760 29440 190920 29600
rect 190760 29600 190920 29760
rect 190760 29760 190920 29920
rect 190760 29920 190920 30080
rect 190760 30080 190920 30240
rect 190760 30240 190920 30400
rect 190760 30400 190920 30560
rect 190760 30560 190920 30720
rect 190760 30720 190920 30880
rect 190760 30880 190920 31040
rect 190760 31040 190920 31200
rect 190760 31200 190920 31360
rect 190760 31360 190920 31520
rect 190760 31520 190920 31680
rect 190760 31680 190920 31840
rect 190760 31840 190920 32000
rect 190760 32000 190920 32160
rect 190920 26080 191080 26240
rect 190920 26240 191080 26400
rect 190920 26400 191080 26560
rect 190920 26560 191080 26720
rect 190920 26720 191080 26880
rect 190920 26880 191080 27040
rect 190920 27040 191080 27200
rect 190920 27200 191080 27360
rect 190920 27360 191080 27520
rect 190920 27520 191080 27680
rect 190920 27680 191080 27840
rect 190920 27840 191080 28000
rect 190920 28000 191080 28160
rect 190920 28160 191080 28320
rect 190920 28320 191080 28480
rect 190920 28480 191080 28640
rect 190920 28640 191080 28800
rect 190920 28800 191080 28960
rect 190920 28960 191080 29120
rect 190920 29120 191080 29280
rect 190920 29280 191080 29440
rect 190920 29440 191080 29600
rect 190920 29600 191080 29760
rect 190920 29760 191080 29920
rect 190920 29920 191080 30080
rect 190920 30080 191080 30240
rect 190920 30240 191080 30400
rect 190920 30400 191080 30560
rect 190920 30560 191080 30720
rect 190920 30720 191080 30880
rect 190920 30880 191080 31040
rect 190920 31040 191080 31200
rect 190920 31200 191080 31360
rect 190920 31360 191080 31520
rect 190920 31520 191080 31680
rect 191080 26080 191240 26240
rect 191080 26240 191240 26400
rect 191080 26400 191240 26560
rect 191080 26560 191240 26720
rect 191080 26720 191240 26880
rect 191080 26880 191240 27040
rect 191080 27040 191240 27200
rect 191080 27200 191240 27360
rect 191080 27360 191240 27520
rect 191080 27520 191240 27680
rect 191080 27680 191240 27840
rect 191080 27840 191240 28000
rect 191080 28000 191240 28160
rect 191080 28160 191240 28320
rect 191080 28320 191240 28480
rect 191080 28480 191240 28640
rect 191080 28640 191240 28800
rect 191080 28800 191240 28960
rect 191080 28960 191240 29120
rect 191080 29120 191240 29280
rect 191080 29280 191240 29440
rect 191080 29440 191240 29600
rect 191080 29600 191240 29760
rect 191080 29760 191240 29920
rect 191080 29920 191240 30080
rect 191080 30080 191240 30240
rect 191080 30240 191240 30400
rect 191080 30400 191240 30560
rect 191080 30560 191240 30720
rect 191080 30720 191240 30880
rect 191080 30880 191240 31040
rect 191080 31040 191240 31200
rect 191080 31200 191240 31360
rect 191080 31360 191240 31520
rect 191080 31520 191240 31680
rect 191080 31680 191240 31840
rect 191080 31840 191240 32000
rect 191240 26240 191400 26400
rect 191240 26400 191400 26560
rect 191240 26560 191400 26720
rect 191240 26720 191400 26880
rect 191240 26880 191400 27040
rect 191240 27040 191400 27200
rect 191240 27200 191400 27360
rect 191240 27360 191400 27520
rect 191240 27520 191400 27680
rect 191240 27680 191400 27840
rect 191240 27840 191400 28000
rect 191240 28000 191400 28160
rect 191240 28160 191400 28320
rect 191240 28320 191400 28480
rect 191240 28480 191400 28640
rect 191240 28640 191400 28800
rect 191240 28800 191400 28960
rect 191240 28960 191400 29120
rect 191240 29120 191400 29280
rect 191240 29280 191400 29440
rect 191240 29440 191400 29600
rect 191240 29600 191400 29760
rect 191240 29760 191400 29920
rect 191240 29920 191400 30080
rect 191240 30080 191400 30240
rect 191240 30240 191400 30400
rect 191240 30400 191400 30560
rect 191240 30560 191400 30720
rect 191240 30720 191400 30880
rect 191240 30880 191400 31040
rect 191240 31040 191400 31200
rect 191240 31200 191400 31360
rect 191240 31360 191400 31520
rect 191240 31520 191400 31680
rect 191240 31680 191400 31840
rect 191240 31840 191400 32000
rect 191240 32000 191400 32160
rect 191240 32160 191400 32320
rect 191400 26240 191560 26400
rect 191400 26400 191560 26560
rect 191400 26560 191560 26720
rect 191400 26720 191560 26880
rect 191400 26880 191560 27040
rect 191400 27040 191560 27200
rect 191400 27200 191560 27360
rect 191400 27360 191560 27520
rect 191400 27520 191560 27680
rect 191400 27680 191560 27840
rect 191400 27840 191560 28000
rect 191400 28000 191560 28160
rect 191400 28160 191560 28320
rect 191400 28320 191560 28480
rect 191400 28480 191560 28640
rect 191400 28640 191560 28800
rect 191400 28800 191560 28960
rect 191400 28960 191560 29120
rect 191400 29120 191560 29280
rect 191400 29280 191560 29440
rect 191400 29440 191560 29600
rect 191400 29600 191560 29760
rect 191400 29760 191560 29920
rect 191400 29920 191560 30080
rect 191400 30080 191560 30240
rect 191400 30240 191560 30400
rect 191400 30400 191560 30560
rect 191400 30560 191560 30720
rect 191400 30720 191560 30880
rect 191400 30880 191560 31040
rect 191400 31040 191560 31200
rect 191400 31200 191560 31360
rect 191400 31360 191560 31520
rect 191400 31520 191560 31680
rect 191400 31680 191560 31840
rect 191400 31840 191560 32000
rect 191400 32000 191560 32160
rect 191400 32160 191560 32320
rect 191400 32320 191560 32480
rect 191400 32480 191560 32640
rect 191560 26240 191720 26400
rect 191560 26400 191720 26560
rect 191560 26560 191720 26720
rect 191560 26720 191720 26880
rect 191560 26880 191720 27040
rect 191560 27040 191720 27200
rect 191560 27200 191720 27360
rect 191560 27360 191720 27520
rect 191560 27520 191720 27680
rect 191560 27680 191720 27840
rect 191560 27840 191720 28000
rect 191560 28000 191720 28160
rect 191560 28160 191720 28320
rect 191560 28320 191720 28480
rect 191560 28480 191720 28640
rect 191560 28640 191720 28800
rect 191560 28800 191720 28960
rect 191560 28960 191720 29120
rect 191560 29120 191720 29280
rect 191560 29280 191720 29440
rect 191560 29440 191720 29600
rect 191560 29600 191720 29760
rect 191560 29760 191720 29920
rect 191560 29920 191720 30080
rect 191560 30080 191720 30240
rect 191560 30240 191720 30400
rect 191560 30400 191720 30560
rect 191560 30560 191720 30720
rect 191560 30720 191720 30880
rect 191560 30880 191720 31040
rect 191560 31040 191720 31200
rect 191560 31200 191720 31360
rect 191560 31360 191720 31520
rect 191560 31520 191720 31680
rect 191560 31680 191720 31840
rect 191560 31840 191720 32000
rect 191560 32000 191720 32160
rect 191560 32160 191720 32320
rect 191560 32320 191720 32480
rect 191560 32480 191720 32640
rect 191560 32640 191720 32800
rect 191560 32800 191720 32960
rect 191560 32960 191720 33120
rect 191720 26400 191880 26560
rect 191720 26560 191880 26720
rect 191720 26720 191880 26880
rect 191720 26880 191880 27040
rect 191720 27040 191880 27200
rect 191720 27200 191880 27360
rect 191720 27360 191880 27520
rect 191720 27520 191880 27680
rect 191720 27680 191880 27840
rect 191720 27840 191880 28000
rect 191720 28000 191880 28160
rect 191720 28160 191880 28320
rect 191720 28320 191880 28480
rect 191720 28480 191880 28640
rect 191720 28640 191880 28800
rect 191720 28800 191880 28960
rect 191720 28960 191880 29120
rect 191720 29120 191880 29280
rect 191720 29280 191880 29440
rect 191720 29440 191880 29600
rect 191720 29600 191880 29760
rect 191720 29760 191880 29920
rect 191720 29920 191880 30080
rect 191720 30080 191880 30240
rect 191720 30240 191880 30400
rect 191720 30400 191880 30560
rect 191720 30560 191880 30720
rect 191720 30720 191880 30880
rect 191720 30880 191880 31040
rect 191720 31040 191880 31200
rect 191720 31200 191880 31360
rect 191720 31360 191880 31520
rect 191720 31520 191880 31680
rect 191720 31680 191880 31840
rect 191720 31840 191880 32000
rect 191720 32000 191880 32160
rect 191720 32160 191880 32320
rect 191720 32320 191880 32480
rect 191720 32480 191880 32640
rect 191720 32640 191880 32800
rect 191720 32800 191880 32960
rect 191720 32960 191880 33120
rect 191720 33120 191880 33280
rect 191720 33280 191880 33440
rect 191880 26560 192040 26720
rect 191880 26720 192040 26880
rect 191880 26880 192040 27040
rect 191880 27040 192040 27200
rect 191880 27200 192040 27360
rect 191880 27360 192040 27520
rect 191880 27520 192040 27680
rect 191880 27680 192040 27840
rect 191880 27840 192040 28000
rect 191880 28000 192040 28160
rect 191880 28160 192040 28320
rect 191880 28320 192040 28480
rect 191880 28480 192040 28640
rect 191880 28640 192040 28800
rect 191880 28800 192040 28960
rect 191880 28960 192040 29120
rect 191880 29120 192040 29280
rect 191880 29280 192040 29440
rect 191880 29440 192040 29600
rect 191880 29600 192040 29760
rect 191880 29760 192040 29920
rect 191880 29920 192040 30080
rect 191880 30080 192040 30240
rect 191880 30240 192040 30400
rect 191880 30400 192040 30560
rect 191880 30560 192040 30720
rect 191880 30720 192040 30880
rect 191880 30880 192040 31040
rect 191880 31040 192040 31200
rect 191880 31200 192040 31360
rect 191880 31360 192040 31520
rect 191880 31520 192040 31680
rect 191880 31680 192040 31840
rect 191880 31840 192040 32000
rect 191880 32000 192040 32160
rect 191880 32160 192040 32320
rect 191880 32320 192040 32480
rect 191880 32480 192040 32640
rect 191880 32640 192040 32800
rect 191880 32800 192040 32960
rect 191880 32960 192040 33120
rect 191880 33120 192040 33280
rect 191880 33280 192040 33440
rect 191880 33440 192040 33600
rect 191880 33600 192040 33760
rect 191880 33760 192040 33920
rect 192040 26720 192200 26880
rect 192040 26880 192200 27040
rect 192040 27040 192200 27200
rect 192040 27200 192200 27360
rect 192040 27360 192200 27520
rect 192040 27520 192200 27680
rect 192040 27680 192200 27840
rect 192040 27840 192200 28000
rect 192040 28000 192200 28160
rect 192040 28160 192200 28320
rect 192040 28320 192200 28480
rect 192040 28480 192200 28640
rect 192040 28640 192200 28800
rect 192040 28800 192200 28960
rect 192040 28960 192200 29120
rect 192040 29120 192200 29280
rect 192040 29280 192200 29440
rect 192040 29440 192200 29600
rect 192040 29600 192200 29760
rect 192040 29760 192200 29920
rect 192040 29920 192200 30080
rect 192040 30080 192200 30240
rect 192040 30240 192200 30400
rect 192040 30400 192200 30560
rect 192040 30560 192200 30720
rect 192040 30720 192200 30880
rect 192040 30880 192200 31040
rect 192040 31040 192200 31200
rect 192040 31200 192200 31360
rect 192040 31360 192200 31520
rect 192040 31520 192200 31680
rect 192040 31680 192200 31840
rect 192040 31840 192200 32000
rect 192040 32000 192200 32160
rect 192040 32160 192200 32320
rect 192040 32320 192200 32480
rect 192040 32480 192200 32640
rect 192040 32640 192200 32800
rect 192040 32800 192200 32960
rect 192040 32960 192200 33120
rect 192040 33120 192200 33280
rect 192040 33280 192200 33440
rect 192040 33440 192200 33600
rect 192040 33600 192200 33760
rect 192040 33760 192200 33920
rect 192040 33920 192200 34080
rect 192040 34080 192200 34240
rect 192200 26880 192360 27040
rect 192200 27040 192360 27200
rect 192200 27200 192360 27360
rect 192200 27360 192360 27520
rect 192200 27520 192360 27680
rect 192200 27680 192360 27840
rect 192200 27840 192360 28000
rect 192200 28000 192360 28160
rect 192200 28160 192360 28320
rect 192200 28320 192360 28480
rect 192200 28480 192360 28640
rect 192200 28640 192360 28800
rect 192200 28800 192360 28960
rect 192200 28960 192360 29120
rect 192200 29120 192360 29280
rect 192200 29280 192360 29440
rect 192200 29440 192360 29600
rect 192200 29600 192360 29760
rect 192200 29760 192360 29920
rect 192200 29920 192360 30080
rect 192200 30080 192360 30240
rect 192200 30240 192360 30400
rect 192200 30400 192360 30560
rect 192200 30560 192360 30720
rect 192200 30720 192360 30880
rect 192200 30880 192360 31040
rect 192200 31040 192360 31200
rect 192200 31200 192360 31360
rect 192200 31360 192360 31520
rect 192200 31520 192360 31680
rect 192200 31680 192360 31840
rect 192200 31840 192360 32000
rect 192200 32000 192360 32160
rect 192200 32160 192360 32320
rect 192200 32320 192360 32480
rect 192200 32480 192360 32640
rect 192200 32640 192360 32800
rect 192200 32800 192360 32960
rect 192200 32960 192360 33120
rect 192200 33120 192360 33280
rect 192200 33280 192360 33440
rect 192200 33440 192360 33600
rect 192200 33600 192360 33760
rect 192200 33760 192360 33920
rect 192200 33920 192360 34080
rect 192200 34080 192360 34240
rect 192200 34240 192360 34400
rect 192200 34400 192360 34560
rect 192200 34560 192360 34720
rect 192360 27200 192520 27360
rect 192360 27360 192520 27520
rect 192360 27520 192520 27680
rect 192360 27680 192520 27840
rect 192360 27840 192520 28000
rect 192360 28000 192520 28160
rect 192360 28160 192520 28320
rect 192360 28320 192520 28480
rect 192360 28480 192520 28640
rect 192360 28640 192520 28800
rect 192360 28800 192520 28960
rect 192360 28960 192520 29120
rect 192360 29120 192520 29280
rect 192360 29280 192520 29440
rect 192360 29440 192520 29600
rect 192360 29600 192520 29760
rect 192360 29760 192520 29920
rect 192360 29920 192520 30080
rect 192360 30080 192520 30240
rect 192360 30240 192520 30400
rect 192360 30400 192520 30560
rect 192360 30560 192520 30720
rect 192360 30720 192520 30880
rect 192360 30880 192520 31040
rect 192360 31040 192520 31200
rect 192360 31200 192520 31360
rect 192360 31360 192520 31520
rect 192360 31520 192520 31680
rect 192360 31680 192520 31840
rect 192360 31840 192520 32000
rect 192360 32000 192520 32160
rect 192360 32160 192520 32320
rect 192360 32320 192520 32480
rect 192360 32480 192520 32640
rect 192360 32640 192520 32800
rect 192360 32800 192520 32960
rect 192360 32960 192520 33120
rect 192360 33120 192520 33280
rect 192360 33280 192520 33440
rect 192360 33440 192520 33600
rect 192360 33600 192520 33760
rect 192360 33760 192520 33920
rect 192360 33920 192520 34080
rect 192360 34080 192520 34240
rect 192360 34240 192520 34400
rect 192360 34400 192520 34560
rect 192360 34560 192520 34720
rect 192360 34720 192520 34880
rect 192360 34880 192520 35040
rect 192520 27520 192680 27680
rect 192520 27680 192680 27840
rect 192520 27840 192680 28000
rect 192520 28000 192680 28160
rect 192520 28160 192680 28320
rect 192520 28320 192680 28480
rect 192520 28480 192680 28640
rect 192520 28640 192680 28800
rect 192520 28800 192680 28960
rect 192520 28960 192680 29120
rect 192520 29120 192680 29280
rect 192520 29280 192680 29440
rect 192520 29440 192680 29600
rect 192520 29600 192680 29760
rect 192520 29760 192680 29920
rect 192520 29920 192680 30080
rect 192520 30080 192680 30240
rect 192520 30240 192680 30400
rect 192520 30400 192680 30560
rect 192520 30560 192680 30720
rect 192520 30720 192680 30880
rect 192520 30880 192680 31040
rect 192520 31040 192680 31200
rect 192520 31200 192680 31360
rect 192520 31360 192680 31520
rect 192520 31520 192680 31680
rect 192520 31680 192680 31840
rect 192520 31840 192680 32000
rect 192520 32000 192680 32160
rect 192520 32160 192680 32320
rect 192520 32320 192680 32480
rect 192520 32480 192680 32640
rect 192520 32640 192680 32800
rect 192520 32800 192680 32960
rect 192520 32960 192680 33120
rect 192520 33120 192680 33280
rect 192520 33280 192680 33440
rect 192520 33440 192680 33600
rect 192520 33600 192680 33760
rect 192520 33760 192680 33920
rect 192520 33920 192680 34080
rect 192520 34080 192680 34240
rect 192520 34240 192680 34400
rect 192520 34400 192680 34560
rect 192520 34560 192680 34720
rect 192520 34720 192680 34880
rect 192520 34880 192680 35040
rect 192520 35040 192680 35200
rect 192520 35200 192680 35360
rect 192520 35360 192680 35520
rect 192680 27840 192840 28000
rect 192680 28000 192840 28160
rect 192680 28160 192840 28320
rect 192680 28320 192840 28480
rect 192680 28480 192840 28640
rect 192680 28640 192840 28800
rect 192680 28800 192840 28960
rect 192680 28960 192840 29120
rect 192680 29120 192840 29280
rect 192680 29280 192840 29440
rect 192680 29440 192840 29600
rect 192680 29600 192840 29760
rect 192680 29760 192840 29920
rect 192680 29920 192840 30080
rect 192680 30080 192840 30240
rect 192680 30240 192840 30400
rect 192680 30400 192840 30560
rect 192680 30560 192840 30720
rect 192680 30720 192840 30880
rect 192680 30880 192840 31040
rect 192680 31040 192840 31200
rect 192680 31200 192840 31360
rect 192680 31360 192840 31520
rect 192680 31520 192840 31680
rect 192680 31680 192840 31840
rect 192680 31840 192840 32000
rect 192680 32000 192840 32160
rect 192680 32160 192840 32320
rect 192680 32320 192840 32480
rect 192680 32480 192840 32640
rect 192680 32640 192840 32800
rect 192680 32800 192840 32960
rect 192680 32960 192840 33120
rect 192680 33120 192840 33280
rect 192680 33280 192840 33440
rect 192680 33440 192840 33600
rect 192680 33600 192840 33760
rect 192680 33760 192840 33920
rect 192680 33920 192840 34080
rect 192680 34080 192840 34240
rect 192680 34240 192840 34400
rect 192680 34400 192840 34560
rect 192680 34560 192840 34720
rect 192680 34720 192840 34880
rect 192680 34880 192840 35040
rect 192680 35040 192840 35200
rect 192680 35200 192840 35360
rect 192680 35360 192840 35520
rect 192680 35520 192840 35680
rect 192680 35680 192840 35840
rect 192680 35840 192840 36000
rect 192840 28320 193000 28480
rect 192840 28480 193000 28640
rect 192840 28640 193000 28800
rect 192840 28800 193000 28960
rect 192840 28960 193000 29120
rect 192840 29120 193000 29280
rect 192840 29280 193000 29440
rect 192840 29440 193000 29600
rect 192840 29600 193000 29760
rect 192840 29760 193000 29920
rect 192840 29920 193000 30080
rect 192840 30080 193000 30240
rect 192840 30240 193000 30400
rect 192840 30400 193000 30560
rect 192840 30560 193000 30720
rect 192840 30720 193000 30880
rect 192840 30880 193000 31040
rect 192840 31040 193000 31200
rect 192840 31200 193000 31360
rect 192840 31360 193000 31520
rect 192840 31520 193000 31680
rect 192840 31680 193000 31840
rect 192840 31840 193000 32000
rect 192840 32000 193000 32160
rect 192840 32160 193000 32320
rect 192840 32320 193000 32480
rect 192840 32480 193000 32640
rect 192840 32640 193000 32800
rect 192840 32800 193000 32960
rect 192840 32960 193000 33120
rect 192840 33120 193000 33280
rect 192840 33280 193000 33440
rect 192840 33440 193000 33600
rect 192840 33600 193000 33760
rect 192840 33760 193000 33920
rect 192840 33920 193000 34080
rect 192840 34080 193000 34240
rect 192840 34240 193000 34400
rect 192840 34400 193000 34560
rect 192840 34560 193000 34720
rect 192840 34720 193000 34880
rect 192840 34880 193000 35040
rect 192840 35040 193000 35200
rect 192840 35200 193000 35360
rect 192840 35360 193000 35520
rect 192840 35520 193000 35680
rect 192840 35680 193000 35840
rect 192840 35840 193000 36000
rect 192840 36000 193000 36160
rect 192840 36160 193000 36320
rect 193000 28640 193160 28800
rect 193000 28800 193160 28960
rect 193000 28960 193160 29120
rect 193000 29120 193160 29280
rect 193000 29280 193160 29440
rect 193000 29440 193160 29600
rect 193000 29600 193160 29760
rect 193000 29760 193160 29920
rect 193000 29920 193160 30080
rect 193000 30080 193160 30240
rect 193000 30240 193160 30400
rect 193000 30400 193160 30560
rect 193000 30560 193160 30720
rect 193000 30720 193160 30880
rect 193000 30880 193160 31040
rect 193000 31040 193160 31200
rect 193000 31200 193160 31360
rect 193000 31360 193160 31520
rect 193000 31520 193160 31680
rect 193000 31680 193160 31840
rect 193000 31840 193160 32000
rect 193000 32000 193160 32160
rect 193000 32160 193160 32320
rect 193000 32320 193160 32480
rect 193000 32480 193160 32640
rect 193000 32640 193160 32800
rect 193000 32800 193160 32960
rect 193000 32960 193160 33120
rect 193000 33120 193160 33280
rect 193000 33280 193160 33440
rect 193000 33440 193160 33600
rect 193000 33600 193160 33760
rect 193000 33760 193160 33920
rect 193000 33920 193160 34080
rect 193000 34080 193160 34240
rect 193000 34240 193160 34400
rect 193000 34400 193160 34560
rect 193000 34560 193160 34720
rect 193000 34720 193160 34880
rect 193000 34880 193160 35040
rect 193000 35040 193160 35200
rect 193000 35200 193160 35360
rect 193000 35360 193160 35520
rect 193000 35520 193160 35680
rect 193000 35680 193160 35840
rect 193000 35840 193160 36000
rect 193000 36000 193160 36160
rect 193000 36160 193160 36320
rect 193000 36320 193160 36480
rect 193000 36480 193160 36640
rect 193000 36640 193160 36800
rect 193160 28960 193320 29120
rect 193160 29120 193320 29280
rect 193160 29280 193320 29440
rect 193160 29440 193320 29600
rect 193160 29600 193320 29760
rect 193160 29760 193320 29920
rect 193160 29920 193320 30080
rect 193160 30080 193320 30240
rect 193160 30240 193320 30400
rect 193160 30400 193320 30560
rect 193160 30560 193320 30720
rect 193160 30720 193320 30880
rect 193160 30880 193320 31040
rect 193160 31040 193320 31200
rect 193160 31200 193320 31360
rect 193160 31360 193320 31520
rect 193160 31520 193320 31680
rect 193160 31680 193320 31840
rect 193160 31840 193320 32000
rect 193160 32000 193320 32160
rect 193160 32160 193320 32320
rect 193160 32320 193320 32480
rect 193160 32480 193320 32640
rect 193160 32640 193320 32800
rect 193160 32800 193320 32960
rect 193160 32960 193320 33120
rect 193160 33120 193320 33280
rect 193160 33280 193320 33440
rect 193160 33440 193320 33600
rect 193160 33600 193320 33760
rect 193160 33760 193320 33920
rect 193160 33920 193320 34080
rect 193160 34080 193320 34240
rect 193160 34240 193320 34400
rect 193160 34400 193320 34560
rect 193160 34560 193320 34720
rect 193160 34720 193320 34880
rect 193160 34880 193320 35040
rect 193160 35040 193320 35200
rect 193160 35200 193320 35360
rect 193160 35360 193320 35520
rect 193160 35520 193320 35680
rect 193160 35680 193320 35840
rect 193160 35840 193320 36000
rect 193160 36000 193320 36160
rect 193160 36160 193320 36320
rect 193160 36320 193320 36480
rect 193160 36480 193320 36640
rect 193160 36640 193320 36800
rect 193160 36800 193320 36960
rect 193160 36960 193320 37120
rect 193320 29440 193480 29600
rect 193320 29600 193480 29760
rect 193320 29760 193480 29920
rect 193320 29920 193480 30080
rect 193320 30080 193480 30240
rect 193320 30240 193480 30400
rect 193320 30400 193480 30560
rect 193320 30560 193480 30720
rect 193320 30720 193480 30880
rect 193320 30880 193480 31040
rect 193320 31040 193480 31200
rect 193320 31200 193480 31360
rect 193320 31360 193480 31520
rect 193320 31520 193480 31680
rect 193320 31680 193480 31840
rect 193320 31840 193480 32000
rect 193320 32000 193480 32160
rect 193320 32160 193480 32320
rect 193320 32320 193480 32480
rect 193320 32480 193480 32640
rect 193320 32640 193480 32800
rect 193320 32800 193480 32960
rect 193320 32960 193480 33120
rect 193320 33120 193480 33280
rect 193320 33280 193480 33440
rect 193320 33440 193480 33600
rect 193320 33600 193480 33760
rect 193320 33760 193480 33920
rect 193320 33920 193480 34080
rect 193320 34080 193480 34240
rect 193320 34240 193480 34400
rect 193320 34400 193480 34560
rect 193320 34560 193480 34720
rect 193320 34720 193480 34880
rect 193320 34880 193480 35040
rect 193320 35040 193480 35200
rect 193320 35200 193480 35360
rect 193320 35360 193480 35520
rect 193320 35520 193480 35680
rect 193320 35680 193480 35840
rect 193320 35840 193480 36000
rect 193320 36000 193480 36160
rect 193320 36160 193480 36320
rect 193320 36320 193480 36480
rect 193320 36480 193480 36640
rect 193320 36640 193480 36800
rect 193320 36800 193480 36960
rect 193320 36960 193480 37120
rect 193320 37120 193480 37280
rect 193320 37280 193480 37440
rect 193320 37440 193480 37600
rect 193480 29760 193640 29920
rect 193480 29920 193640 30080
rect 193480 30080 193640 30240
rect 193480 30240 193640 30400
rect 193480 30400 193640 30560
rect 193480 30560 193640 30720
rect 193480 30720 193640 30880
rect 193480 30880 193640 31040
rect 193480 31040 193640 31200
rect 193480 31200 193640 31360
rect 193480 31360 193640 31520
rect 193480 31520 193640 31680
rect 193480 31680 193640 31840
rect 193480 31840 193640 32000
rect 193480 32000 193640 32160
rect 193480 32160 193640 32320
rect 193480 32320 193640 32480
rect 193480 32480 193640 32640
rect 193480 32640 193640 32800
rect 193480 32800 193640 32960
rect 193480 32960 193640 33120
rect 193480 33120 193640 33280
rect 193480 33280 193640 33440
rect 193480 33440 193640 33600
rect 193480 33600 193640 33760
rect 193480 33760 193640 33920
rect 193480 33920 193640 34080
rect 193480 34080 193640 34240
rect 193480 34240 193640 34400
rect 193480 34400 193640 34560
rect 193480 34560 193640 34720
rect 193480 34720 193640 34880
rect 193480 34880 193640 35040
rect 193480 35040 193640 35200
rect 193480 35200 193640 35360
rect 193480 35360 193640 35520
rect 193480 35520 193640 35680
rect 193480 35680 193640 35840
rect 193480 35840 193640 36000
rect 193480 36000 193640 36160
rect 193480 36160 193640 36320
rect 193480 36320 193640 36480
rect 193480 36480 193640 36640
rect 193480 36640 193640 36800
rect 193480 36800 193640 36960
rect 193480 36960 193640 37120
rect 193480 37120 193640 37280
rect 193480 37280 193640 37440
rect 193480 37440 193640 37600
rect 193480 37600 193640 37760
rect 193480 37760 193640 37920
rect 193640 30240 193800 30400
rect 193640 30400 193800 30560
rect 193640 30560 193800 30720
rect 193640 30720 193800 30880
rect 193640 30880 193800 31040
rect 193640 31040 193800 31200
rect 193640 31200 193800 31360
rect 193640 31360 193800 31520
rect 193640 31520 193800 31680
rect 193640 31680 193800 31840
rect 193640 31840 193800 32000
rect 193640 32000 193800 32160
rect 193640 32160 193800 32320
rect 193640 32320 193800 32480
rect 193640 32480 193800 32640
rect 193640 32640 193800 32800
rect 193640 32800 193800 32960
rect 193640 32960 193800 33120
rect 193640 33120 193800 33280
rect 193640 33280 193800 33440
rect 193640 33440 193800 33600
rect 193640 33600 193800 33760
rect 193640 33760 193800 33920
rect 193640 33920 193800 34080
rect 193640 34080 193800 34240
rect 193640 34240 193800 34400
rect 193640 34400 193800 34560
rect 193640 34560 193800 34720
rect 193640 34720 193800 34880
rect 193640 34880 193800 35040
rect 193640 35040 193800 35200
rect 193640 35200 193800 35360
rect 193640 35360 193800 35520
rect 193640 35520 193800 35680
rect 193640 35680 193800 35840
rect 193640 35840 193800 36000
rect 193640 36000 193800 36160
rect 193640 36160 193800 36320
rect 193640 36320 193800 36480
rect 193640 36480 193800 36640
rect 193640 36640 193800 36800
rect 193640 36800 193800 36960
rect 193640 36960 193800 37120
rect 193640 37120 193800 37280
rect 193640 37280 193800 37440
rect 193640 37440 193800 37600
rect 193640 37600 193800 37760
rect 193640 37760 193800 37920
rect 193640 37920 193800 38080
rect 193640 38080 193800 38240
rect 193640 38240 193800 38400
rect 193800 30560 193960 30720
rect 193800 30720 193960 30880
rect 193800 30880 193960 31040
rect 193800 31040 193960 31200
rect 193800 31200 193960 31360
rect 193800 31360 193960 31520
rect 193800 31520 193960 31680
rect 193800 31680 193960 31840
rect 193800 31840 193960 32000
rect 193800 32000 193960 32160
rect 193800 32160 193960 32320
rect 193800 32320 193960 32480
rect 193800 32480 193960 32640
rect 193800 32640 193960 32800
rect 193800 32800 193960 32960
rect 193800 32960 193960 33120
rect 193800 33120 193960 33280
rect 193800 33280 193960 33440
rect 193800 33440 193960 33600
rect 193800 33600 193960 33760
rect 193800 33760 193960 33920
rect 193800 33920 193960 34080
rect 193800 34080 193960 34240
rect 193800 34240 193960 34400
rect 193800 34400 193960 34560
rect 193800 34560 193960 34720
rect 193800 34720 193960 34880
rect 193800 34880 193960 35040
rect 193800 35040 193960 35200
rect 193800 35200 193960 35360
rect 193800 35360 193960 35520
rect 193800 35520 193960 35680
rect 193800 35680 193960 35840
rect 193800 35840 193960 36000
rect 193800 36000 193960 36160
rect 193800 36160 193960 36320
rect 193800 36320 193960 36480
rect 193800 36480 193960 36640
rect 193800 36640 193960 36800
rect 193800 36800 193960 36960
rect 193800 36960 193960 37120
rect 193800 37120 193960 37280
rect 193800 37280 193960 37440
rect 193800 37440 193960 37600
rect 193800 37600 193960 37760
rect 193800 37760 193960 37920
rect 193800 37920 193960 38080
rect 193800 38080 193960 38240
rect 193800 38240 193960 38400
rect 193800 38400 193960 38560
rect 193800 38560 193960 38720
rect 193800 38720 193960 38880
rect 193960 30880 194120 31040
rect 193960 31040 194120 31200
rect 193960 31200 194120 31360
rect 193960 31360 194120 31520
rect 193960 31520 194120 31680
rect 193960 31680 194120 31840
rect 193960 31840 194120 32000
rect 193960 32000 194120 32160
rect 193960 32160 194120 32320
rect 193960 32320 194120 32480
rect 193960 32480 194120 32640
rect 193960 32640 194120 32800
rect 193960 32800 194120 32960
rect 193960 32960 194120 33120
rect 193960 33120 194120 33280
rect 193960 33280 194120 33440
rect 193960 33440 194120 33600
rect 193960 33600 194120 33760
rect 193960 33760 194120 33920
rect 193960 33920 194120 34080
rect 193960 34080 194120 34240
rect 193960 34240 194120 34400
rect 193960 34400 194120 34560
rect 193960 34560 194120 34720
rect 193960 34720 194120 34880
rect 193960 34880 194120 35040
rect 193960 35040 194120 35200
rect 193960 35200 194120 35360
rect 193960 35360 194120 35520
rect 193960 35520 194120 35680
rect 193960 35680 194120 35840
rect 193960 35840 194120 36000
rect 193960 36000 194120 36160
rect 193960 36160 194120 36320
rect 193960 36320 194120 36480
rect 193960 36480 194120 36640
rect 193960 36640 194120 36800
rect 193960 36800 194120 36960
rect 193960 36960 194120 37120
rect 193960 37120 194120 37280
rect 193960 37280 194120 37440
rect 193960 37440 194120 37600
rect 193960 37600 194120 37760
rect 193960 37760 194120 37920
rect 193960 37920 194120 38080
rect 193960 38080 194120 38240
rect 193960 38240 194120 38400
rect 193960 38400 194120 38560
rect 193960 38560 194120 38720
rect 193960 38720 194120 38880
rect 193960 38880 194120 39040
rect 193960 39040 194120 39200
rect 194120 31360 194280 31520
rect 194120 31520 194280 31680
rect 194120 31680 194280 31840
rect 194120 31840 194280 32000
rect 194120 32000 194280 32160
rect 194120 32160 194280 32320
rect 194120 32320 194280 32480
rect 194120 32480 194280 32640
rect 194120 32640 194280 32800
rect 194120 32800 194280 32960
rect 194120 32960 194280 33120
rect 194120 33120 194280 33280
rect 194120 33280 194280 33440
rect 194120 33440 194280 33600
rect 194120 33600 194280 33760
rect 194120 33760 194280 33920
rect 194120 33920 194280 34080
rect 194120 34080 194280 34240
rect 194120 34240 194280 34400
rect 194120 34400 194280 34560
rect 194120 34560 194280 34720
rect 194120 34720 194280 34880
rect 194120 34880 194280 35040
rect 194120 35040 194280 35200
rect 194120 35200 194280 35360
rect 194120 35360 194280 35520
rect 194120 35520 194280 35680
rect 194120 35680 194280 35840
rect 194120 35840 194280 36000
rect 194120 36000 194280 36160
rect 194120 36160 194280 36320
rect 194120 36320 194280 36480
rect 194120 36480 194280 36640
rect 194120 36640 194280 36800
rect 194120 36800 194280 36960
rect 194120 36960 194280 37120
rect 194120 37120 194280 37280
rect 194120 37280 194280 37440
rect 194120 37440 194280 37600
rect 194120 37600 194280 37760
rect 194120 37760 194280 37920
rect 194120 37920 194280 38080
rect 194120 38080 194280 38240
rect 194120 38240 194280 38400
rect 194120 38400 194280 38560
rect 194120 38560 194280 38720
rect 194120 38720 194280 38880
rect 194120 38880 194280 39040
rect 194120 39040 194280 39200
rect 194120 39200 194280 39360
rect 194120 39360 194280 39520
rect 194120 39520 194280 39680
rect 194280 31840 194440 32000
rect 194280 32000 194440 32160
rect 194280 32160 194440 32320
rect 194280 32320 194440 32480
rect 194280 32480 194440 32640
rect 194280 32640 194440 32800
rect 194280 32800 194440 32960
rect 194280 32960 194440 33120
rect 194280 33120 194440 33280
rect 194280 33280 194440 33440
rect 194280 33440 194440 33600
rect 194280 33600 194440 33760
rect 194280 33760 194440 33920
rect 194280 33920 194440 34080
rect 194280 34080 194440 34240
rect 194280 34240 194440 34400
rect 194280 34400 194440 34560
rect 194280 34560 194440 34720
rect 194280 34720 194440 34880
rect 194280 34880 194440 35040
rect 194280 35040 194440 35200
rect 194280 35200 194440 35360
rect 194280 35360 194440 35520
rect 194280 35520 194440 35680
rect 194280 35680 194440 35840
rect 194280 35840 194440 36000
rect 194280 36000 194440 36160
rect 194280 36160 194440 36320
rect 194280 36320 194440 36480
rect 194280 36480 194440 36640
rect 194280 36640 194440 36800
rect 194280 36800 194440 36960
rect 194280 36960 194440 37120
rect 194280 37120 194440 37280
rect 194280 37280 194440 37440
rect 194280 37440 194440 37600
rect 194280 37600 194440 37760
rect 194280 37760 194440 37920
rect 194280 37920 194440 38080
rect 194280 38080 194440 38240
rect 194280 38240 194440 38400
rect 194280 38400 194440 38560
rect 194280 38560 194440 38720
rect 194280 38720 194440 38880
rect 194280 38880 194440 39040
rect 194280 39040 194440 39200
rect 194280 39200 194440 39360
rect 194280 39360 194440 39520
rect 194280 39520 194440 39680
rect 194280 39680 194440 39840
rect 194280 39840 194440 40000
rect 194280 40000 194440 40160
rect 194440 32160 194600 32320
rect 194440 32320 194600 32480
rect 194440 32480 194600 32640
rect 194440 32640 194600 32800
rect 194440 32800 194600 32960
rect 194440 32960 194600 33120
rect 194440 33120 194600 33280
rect 194440 33280 194600 33440
rect 194440 33440 194600 33600
rect 194440 33600 194600 33760
rect 194440 33760 194600 33920
rect 194440 33920 194600 34080
rect 194440 34080 194600 34240
rect 194440 34240 194600 34400
rect 194440 34400 194600 34560
rect 194440 34560 194600 34720
rect 194440 34720 194600 34880
rect 194440 34880 194600 35040
rect 194440 35040 194600 35200
rect 194440 35200 194600 35360
rect 194440 35360 194600 35520
rect 194440 35520 194600 35680
rect 194440 35680 194600 35840
rect 194440 35840 194600 36000
rect 194440 36000 194600 36160
rect 194440 36160 194600 36320
rect 194440 36320 194600 36480
rect 194440 36480 194600 36640
rect 194440 36640 194600 36800
rect 194440 36800 194600 36960
rect 194440 36960 194600 37120
rect 194440 37120 194600 37280
rect 194440 37280 194600 37440
rect 194440 37440 194600 37600
rect 194440 37600 194600 37760
rect 194440 37760 194600 37920
rect 194440 37920 194600 38080
rect 194440 38080 194600 38240
rect 194440 38240 194600 38400
rect 194440 38400 194600 38560
rect 194440 38560 194600 38720
rect 194440 38720 194600 38880
rect 194440 38880 194600 39040
rect 194440 39040 194600 39200
rect 194440 39200 194600 39360
rect 194440 39360 194600 39520
rect 194440 39520 194600 39680
rect 194440 39680 194600 39840
rect 194440 39840 194600 40000
rect 194440 40000 194600 40160
rect 194440 40160 194600 40320
rect 194440 40320 194600 40480
rect 194600 32640 194760 32800
rect 194600 32800 194760 32960
rect 194600 32960 194760 33120
rect 194600 33120 194760 33280
rect 194600 33280 194760 33440
rect 194600 33440 194760 33600
rect 194600 33600 194760 33760
rect 194600 33760 194760 33920
rect 194600 33920 194760 34080
rect 194600 34080 194760 34240
rect 194600 34240 194760 34400
rect 194600 34400 194760 34560
rect 194600 34560 194760 34720
rect 194600 34720 194760 34880
rect 194600 34880 194760 35040
rect 194600 35040 194760 35200
rect 194600 35200 194760 35360
rect 194600 35360 194760 35520
rect 194600 35520 194760 35680
rect 194600 35680 194760 35840
rect 194600 35840 194760 36000
rect 194600 36000 194760 36160
rect 194600 36160 194760 36320
rect 194600 36320 194760 36480
rect 194600 36480 194760 36640
rect 194600 36640 194760 36800
rect 194600 36800 194760 36960
rect 194600 36960 194760 37120
rect 194600 37120 194760 37280
rect 194600 37280 194760 37440
rect 194600 37440 194760 37600
rect 194600 37600 194760 37760
rect 194600 37760 194760 37920
rect 194600 37920 194760 38080
rect 194600 38080 194760 38240
rect 194600 38240 194760 38400
rect 194600 38400 194760 38560
rect 194600 38560 194760 38720
rect 194600 38720 194760 38880
rect 194600 38880 194760 39040
rect 194600 39040 194760 39200
rect 194600 39200 194760 39360
rect 194600 39360 194760 39520
rect 194600 39520 194760 39680
rect 194600 39680 194760 39840
rect 194600 39840 194760 40000
rect 194600 40000 194760 40160
rect 194600 40160 194760 40320
rect 194600 40320 194760 40480
rect 194600 40480 194760 40640
rect 194600 40640 194760 40800
rect 194600 40800 194760 40960
rect 194760 33120 194920 33280
rect 194760 33280 194920 33440
rect 194760 33440 194920 33600
rect 194760 33600 194920 33760
rect 194760 33760 194920 33920
rect 194760 33920 194920 34080
rect 194760 34080 194920 34240
rect 194760 34240 194920 34400
rect 194760 34400 194920 34560
rect 194760 34560 194920 34720
rect 194760 34720 194920 34880
rect 194760 34880 194920 35040
rect 194760 35040 194920 35200
rect 194760 35200 194920 35360
rect 194760 35360 194920 35520
rect 194760 35520 194920 35680
rect 194760 35680 194920 35840
rect 194760 35840 194920 36000
rect 194760 36000 194920 36160
rect 194760 36160 194920 36320
rect 194760 36320 194920 36480
rect 194760 36480 194920 36640
rect 194760 36640 194920 36800
rect 194760 36800 194920 36960
rect 194760 36960 194920 37120
rect 194760 37120 194920 37280
rect 194760 37280 194920 37440
rect 194760 37440 194920 37600
rect 194760 37600 194920 37760
rect 194760 37760 194920 37920
rect 194760 37920 194920 38080
rect 194760 38080 194920 38240
rect 194760 38240 194920 38400
rect 194760 38400 194920 38560
rect 194760 38560 194920 38720
rect 194760 38720 194920 38880
rect 194760 38880 194920 39040
rect 194760 39040 194920 39200
rect 194760 39200 194920 39360
rect 194760 39360 194920 39520
rect 194760 39520 194920 39680
rect 194760 39680 194920 39840
rect 194760 39840 194920 40000
rect 194760 40000 194920 40160
rect 194760 40160 194920 40320
rect 194760 40320 194920 40480
rect 194760 40480 194920 40640
rect 194760 40640 194920 40800
rect 194760 40800 194920 40960
rect 194760 40960 194920 41120
rect 194760 41120 194920 41280
rect 194920 33440 195080 33600
rect 194920 33600 195080 33760
rect 194920 33760 195080 33920
rect 194920 33920 195080 34080
rect 194920 34080 195080 34240
rect 194920 34240 195080 34400
rect 194920 34400 195080 34560
rect 194920 34560 195080 34720
rect 194920 34720 195080 34880
rect 194920 34880 195080 35040
rect 194920 35040 195080 35200
rect 194920 35200 195080 35360
rect 194920 35360 195080 35520
rect 194920 35520 195080 35680
rect 194920 35680 195080 35840
rect 194920 35840 195080 36000
rect 194920 36000 195080 36160
rect 194920 36160 195080 36320
rect 194920 36320 195080 36480
rect 194920 36480 195080 36640
rect 194920 36640 195080 36800
rect 194920 36800 195080 36960
rect 194920 36960 195080 37120
rect 194920 37120 195080 37280
rect 194920 37280 195080 37440
rect 194920 37440 195080 37600
rect 194920 37600 195080 37760
rect 194920 37760 195080 37920
rect 194920 37920 195080 38080
rect 194920 38080 195080 38240
rect 194920 38240 195080 38400
rect 194920 38400 195080 38560
rect 194920 38560 195080 38720
rect 194920 38720 195080 38880
rect 194920 38880 195080 39040
rect 194920 39040 195080 39200
rect 194920 39200 195080 39360
rect 194920 39360 195080 39520
rect 194920 39520 195080 39680
rect 194920 39680 195080 39840
rect 194920 39840 195080 40000
rect 194920 40000 195080 40160
rect 194920 40160 195080 40320
rect 194920 40320 195080 40480
rect 194920 40480 195080 40640
rect 194920 40640 195080 40800
rect 194920 40800 195080 40960
rect 194920 40960 195080 41120
rect 194920 41120 195080 41280
rect 194920 41280 195080 41440
rect 194920 41440 195080 41600
rect 194920 41600 195080 41760
rect 195080 33760 195240 33920
rect 195080 33920 195240 34080
rect 195080 34080 195240 34240
rect 195080 34240 195240 34400
rect 195080 34400 195240 34560
rect 195080 34560 195240 34720
rect 195080 34720 195240 34880
rect 195080 34880 195240 35040
rect 195080 35040 195240 35200
rect 195080 35200 195240 35360
rect 195080 35360 195240 35520
rect 195080 35520 195240 35680
rect 195080 35680 195240 35840
rect 195080 35840 195240 36000
rect 195080 36000 195240 36160
rect 195080 36160 195240 36320
rect 195080 36320 195240 36480
rect 195080 36480 195240 36640
rect 195080 36640 195240 36800
rect 195080 36800 195240 36960
rect 195080 36960 195240 37120
rect 195080 37120 195240 37280
rect 195080 37280 195240 37440
rect 195080 37440 195240 37600
rect 195080 37600 195240 37760
rect 195080 37760 195240 37920
rect 195080 37920 195240 38080
rect 195080 38080 195240 38240
rect 195080 38240 195240 38400
rect 195080 38400 195240 38560
rect 195080 38560 195240 38720
rect 195080 38720 195240 38880
rect 195080 38880 195240 39040
rect 195080 39040 195240 39200
rect 195080 39200 195240 39360
rect 195080 39360 195240 39520
rect 195080 39520 195240 39680
rect 195080 39680 195240 39840
rect 195080 39840 195240 40000
rect 195080 40000 195240 40160
rect 195080 40160 195240 40320
rect 195080 40320 195240 40480
rect 195080 40480 195240 40640
rect 195080 40640 195240 40800
rect 195080 40800 195240 40960
rect 195080 40960 195240 41120
rect 195080 41120 195240 41280
rect 195080 41280 195240 41440
rect 195080 41440 195240 41600
rect 195080 41600 195240 41760
rect 195080 41760 195240 41920
rect 195080 41920 195240 42080
rect 195080 42080 195240 42240
rect 195240 34240 195400 34400
rect 195240 34400 195400 34560
rect 195240 34560 195400 34720
rect 195240 34720 195400 34880
rect 195240 34880 195400 35040
rect 195240 35040 195400 35200
rect 195240 35200 195400 35360
rect 195240 35360 195400 35520
rect 195240 35520 195400 35680
rect 195240 35680 195400 35840
rect 195240 35840 195400 36000
rect 195240 36000 195400 36160
rect 195240 36160 195400 36320
rect 195240 36320 195400 36480
rect 195240 36480 195400 36640
rect 195240 36640 195400 36800
rect 195240 36800 195400 36960
rect 195240 36960 195400 37120
rect 195240 37120 195400 37280
rect 195240 37280 195400 37440
rect 195240 37440 195400 37600
rect 195240 37600 195400 37760
rect 195240 37760 195400 37920
rect 195240 37920 195400 38080
rect 195240 38080 195400 38240
rect 195240 38240 195400 38400
rect 195240 38400 195400 38560
rect 195240 38560 195400 38720
rect 195240 38720 195400 38880
rect 195240 38880 195400 39040
rect 195240 39040 195400 39200
rect 195240 39200 195400 39360
rect 195240 39360 195400 39520
rect 195240 39520 195400 39680
rect 195240 39680 195400 39840
rect 195240 39840 195400 40000
rect 195240 40000 195400 40160
rect 195240 40160 195400 40320
rect 195240 40320 195400 40480
rect 195240 40480 195400 40640
rect 195240 40640 195400 40800
rect 195240 40800 195400 40960
rect 195240 40960 195400 41120
rect 195240 41120 195400 41280
rect 195240 41280 195400 41440
rect 195240 41440 195400 41600
rect 195240 41600 195400 41760
rect 195240 41760 195400 41920
rect 195240 41920 195400 42080
rect 195240 42080 195400 42240
rect 195240 42240 195400 42400
rect 195240 42400 195400 42560
rect 195400 34560 195560 34720
rect 195400 34720 195560 34880
rect 195400 34880 195560 35040
rect 195400 35040 195560 35200
rect 195400 35200 195560 35360
rect 195400 35360 195560 35520
rect 195400 35520 195560 35680
rect 195400 35680 195560 35840
rect 195400 35840 195560 36000
rect 195400 36000 195560 36160
rect 195400 36160 195560 36320
rect 195400 36320 195560 36480
rect 195400 36480 195560 36640
rect 195400 36640 195560 36800
rect 195400 36800 195560 36960
rect 195400 36960 195560 37120
rect 195400 37120 195560 37280
rect 195400 37280 195560 37440
rect 195400 37440 195560 37600
rect 195400 37600 195560 37760
rect 195400 37760 195560 37920
rect 195400 37920 195560 38080
rect 195400 38080 195560 38240
rect 195400 38240 195560 38400
rect 195400 38400 195560 38560
rect 195400 38560 195560 38720
rect 195400 38720 195560 38880
rect 195400 38880 195560 39040
rect 195400 39040 195560 39200
rect 195400 39200 195560 39360
rect 195400 39360 195560 39520
rect 195400 39520 195560 39680
rect 195400 39680 195560 39840
rect 195400 39840 195560 40000
rect 195400 40000 195560 40160
rect 195400 40160 195560 40320
rect 195400 40320 195560 40480
rect 195400 40480 195560 40640
rect 195400 40640 195560 40800
rect 195400 40800 195560 40960
rect 195400 40960 195560 41120
rect 195400 41120 195560 41280
rect 195400 41280 195560 41440
rect 195400 41440 195560 41600
rect 195400 41600 195560 41760
rect 195400 41760 195560 41920
rect 195400 41920 195560 42080
rect 195400 42080 195560 42240
rect 195400 42240 195560 42400
rect 195400 42400 195560 42560
rect 195400 42560 195560 42720
rect 195400 42720 195560 42880
rect 195400 42880 195560 43040
rect 195560 35040 195720 35200
rect 195560 35200 195720 35360
rect 195560 35360 195720 35520
rect 195560 35520 195720 35680
rect 195560 35680 195720 35840
rect 195560 35840 195720 36000
rect 195560 36000 195720 36160
rect 195560 36160 195720 36320
rect 195560 36320 195720 36480
rect 195560 36480 195720 36640
rect 195560 36640 195720 36800
rect 195560 36800 195720 36960
rect 195560 36960 195720 37120
rect 195560 37120 195720 37280
rect 195560 37280 195720 37440
rect 195560 37440 195720 37600
rect 195560 37600 195720 37760
rect 195560 37760 195720 37920
rect 195560 37920 195720 38080
rect 195560 38080 195720 38240
rect 195560 38240 195720 38400
rect 195560 38400 195720 38560
rect 195560 38560 195720 38720
rect 195560 38720 195720 38880
rect 195560 38880 195720 39040
rect 195560 39040 195720 39200
rect 195560 39200 195720 39360
rect 195560 39360 195720 39520
rect 195560 39520 195720 39680
rect 195560 39680 195720 39840
rect 195560 39840 195720 40000
rect 195560 40000 195720 40160
rect 195560 40160 195720 40320
rect 195560 40320 195720 40480
rect 195560 40480 195720 40640
rect 195560 40640 195720 40800
rect 195560 40800 195720 40960
rect 195560 40960 195720 41120
rect 195560 41120 195720 41280
rect 195560 41280 195720 41440
rect 195560 41440 195720 41600
rect 195560 41600 195720 41760
rect 195560 41760 195720 41920
rect 195560 41920 195720 42080
rect 195560 42080 195720 42240
rect 195560 42240 195720 42400
rect 195560 42400 195720 42560
rect 195560 42560 195720 42720
rect 195560 42720 195720 42880
rect 195560 42880 195720 43040
rect 195560 43040 195720 43200
rect 195560 43200 195720 43360
rect 195560 43360 195720 43520
rect 195720 35360 195880 35520
rect 195720 35520 195880 35680
rect 195720 35680 195880 35840
rect 195720 35840 195880 36000
rect 195720 36000 195880 36160
rect 195720 36160 195880 36320
rect 195720 36320 195880 36480
rect 195720 36480 195880 36640
rect 195720 36640 195880 36800
rect 195720 36800 195880 36960
rect 195720 36960 195880 37120
rect 195720 37120 195880 37280
rect 195720 37280 195880 37440
rect 195720 37440 195880 37600
rect 195720 37600 195880 37760
rect 195720 37760 195880 37920
rect 195720 37920 195880 38080
rect 195720 38080 195880 38240
rect 195720 38240 195880 38400
rect 195720 38400 195880 38560
rect 195720 38560 195880 38720
rect 195720 38720 195880 38880
rect 195720 38880 195880 39040
rect 195720 39040 195880 39200
rect 195720 39200 195880 39360
rect 195720 39360 195880 39520
rect 195720 39520 195880 39680
rect 195720 39680 195880 39840
rect 195720 39840 195880 40000
rect 195720 40000 195880 40160
rect 195720 40160 195880 40320
rect 195720 40320 195880 40480
rect 195720 40480 195880 40640
rect 195720 40640 195880 40800
rect 195720 40800 195880 40960
rect 195720 40960 195880 41120
rect 195720 41120 195880 41280
rect 195720 41280 195880 41440
rect 195720 41440 195880 41600
rect 195720 41600 195880 41760
rect 195720 41760 195880 41920
rect 195720 41920 195880 42080
rect 195720 42080 195880 42240
rect 195720 42240 195880 42400
rect 195720 42400 195880 42560
rect 195720 42560 195880 42720
rect 195720 42720 195880 42880
rect 195720 42880 195880 43040
rect 195720 43040 195880 43200
rect 195720 43200 195880 43360
rect 195720 43360 195880 43520
rect 195720 43520 195880 43680
rect 195720 43680 195880 43840
rect 195720 43840 195880 44000
rect 195880 35840 196040 36000
rect 195880 36000 196040 36160
rect 195880 36160 196040 36320
rect 195880 36320 196040 36480
rect 195880 36480 196040 36640
rect 195880 36640 196040 36800
rect 195880 36800 196040 36960
rect 195880 36960 196040 37120
rect 195880 37120 196040 37280
rect 195880 37280 196040 37440
rect 195880 37440 196040 37600
rect 195880 37600 196040 37760
rect 195880 37760 196040 37920
rect 195880 37920 196040 38080
rect 195880 38080 196040 38240
rect 195880 38240 196040 38400
rect 195880 38400 196040 38560
rect 195880 38560 196040 38720
rect 195880 38720 196040 38880
rect 195880 38880 196040 39040
rect 195880 39040 196040 39200
rect 195880 39200 196040 39360
rect 195880 39360 196040 39520
rect 195880 39520 196040 39680
rect 195880 39680 196040 39840
rect 195880 39840 196040 40000
rect 195880 40000 196040 40160
rect 195880 40160 196040 40320
rect 195880 40320 196040 40480
rect 195880 40480 196040 40640
rect 195880 40640 196040 40800
rect 195880 40800 196040 40960
rect 195880 40960 196040 41120
rect 195880 41120 196040 41280
rect 195880 41280 196040 41440
rect 195880 41440 196040 41600
rect 195880 41600 196040 41760
rect 195880 41760 196040 41920
rect 195880 41920 196040 42080
rect 195880 42080 196040 42240
rect 195880 42240 196040 42400
rect 195880 42400 196040 42560
rect 195880 42560 196040 42720
rect 195880 42720 196040 42880
rect 195880 42880 196040 43040
rect 195880 43040 196040 43200
rect 195880 43200 196040 43360
rect 195880 43360 196040 43520
rect 195880 43520 196040 43680
rect 195880 43680 196040 43840
rect 195880 43840 196040 44000
rect 195880 44000 196040 44160
rect 195880 44160 196040 44320
rect 196040 36160 196200 36320
rect 196040 36320 196200 36480
rect 196040 36480 196200 36640
rect 196040 36640 196200 36800
rect 196040 36800 196200 36960
rect 196040 36960 196200 37120
rect 196040 37120 196200 37280
rect 196040 37280 196200 37440
rect 196040 37440 196200 37600
rect 196040 37600 196200 37760
rect 196040 37760 196200 37920
rect 196040 37920 196200 38080
rect 196040 38080 196200 38240
rect 196040 38240 196200 38400
rect 196040 38400 196200 38560
rect 196040 38560 196200 38720
rect 196040 38720 196200 38880
rect 196040 38880 196200 39040
rect 196040 39040 196200 39200
rect 196040 39200 196200 39360
rect 196040 39360 196200 39520
rect 196040 39520 196200 39680
rect 196040 39680 196200 39840
rect 196040 39840 196200 40000
rect 196040 40000 196200 40160
rect 196040 40160 196200 40320
rect 196040 40320 196200 40480
rect 196040 40480 196200 40640
rect 196040 40640 196200 40800
rect 196040 40800 196200 40960
rect 196040 40960 196200 41120
rect 196040 41120 196200 41280
rect 196040 41280 196200 41440
rect 196040 41440 196200 41600
rect 196040 41600 196200 41760
rect 196040 41760 196200 41920
rect 196040 41920 196200 42080
rect 196040 42080 196200 42240
rect 196040 42240 196200 42400
rect 196040 42400 196200 42560
rect 196040 42560 196200 42720
rect 196040 42720 196200 42880
rect 196040 42880 196200 43040
rect 196040 43040 196200 43200
rect 196040 43200 196200 43360
rect 196040 43360 196200 43520
rect 196040 43520 196200 43680
rect 196040 43680 196200 43840
rect 196040 43840 196200 44000
rect 196040 44000 196200 44160
rect 196040 44160 196200 44320
rect 196040 44320 196200 44480
rect 196040 44480 196200 44640
rect 196040 44640 196200 44800
rect 196200 36640 196360 36800
rect 196200 36800 196360 36960
rect 196200 36960 196360 37120
rect 196200 37120 196360 37280
rect 196200 37280 196360 37440
rect 196200 37440 196360 37600
rect 196200 37600 196360 37760
rect 196200 37760 196360 37920
rect 196200 37920 196360 38080
rect 196200 38080 196360 38240
rect 196200 38240 196360 38400
rect 196200 38400 196360 38560
rect 196200 38560 196360 38720
rect 196200 38720 196360 38880
rect 196200 38880 196360 39040
rect 196200 39040 196360 39200
rect 196200 39200 196360 39360
rect 196200 39360 196360 39520
rect 196200 39520 196360 39680
rect 196200 39680 196360 39840
rect 196200 39840 196360 40000
rect 196200 40000 196360 40160
rect 196200 40160 196360 40320
rect 196200 40320 196360 40480
rect 196200 40480 196360 40640
rect 196200 40640 196360 40800
rect 196200 40800 196360 40960
rect 196200 40960 196360 41120
rect 196200 41120 196360 41280
rect 196200 41280 196360 41440
rect 196200 41440 196360 41600
rect 196200 41600 196360 41760
rect 196200 41760 196360 41920
rect 196200 41920 196360 42080
rect 196200 42080 196360 42240
rect 196200 42240 196360 42400
rect 196200 42400 196360 42560
rect 196200 42560 196360 42720
rect 196200 42720 196360 42880
rect 196200 42880 196360 43040
rect 196200 43040 196360 43200
rect 196200 43200 196360 43360
rect 196200 43360 196360 43520
rect 196200 43520 196360 43680
rect 196200 43680 196360 43840
rect 196200 43840 196360 44000
rect 196200 44000 196360 44160
rect 196200 44160 196360 44320
rect 196200 44320 196360 44480
rect 196200 44480 196360 44640
rect 196200 44640 196360 44800
rect 196200 44800 196360 44960
rect 196200 44960 196360 45120
rect 196200 45120 196360 45280
rect 196360 36960 196520 37120
rect 196360 37120 196520 37280
rect 196360 37280 196520 37440
rect 196360 37440 196520 37600
rect 196360 37600 196520 37760
rect 196360 37760 196520 37920
rect 196360 37920 196520 38080
rect 196360 38080 196520 38240
rect 196360 38240 196520 38400
rect 196360 38400 196520 38560
rect 196360 38560 196520 38720
rect 196360 38720 196520 38880
rect 196360 38880 196520 39040
rect 196360 39040 196520 39200
rect 196360 39200 196520 39360
rect 196360 39360 196520 39520
rect 196360 39520 196520 39680
rect 196360 39680 196520 39840
rect 196360 39840 196520 40000
rect 196360 40000 196520 40160
rect 196360 40160 196520 40320
rect 196360 40320 196520 40480
rect 196360 40480 196520 40640
rect 196360 40640 196520 40800
rect 196360 40800 196520 40960
rect 196360 40960 196520 41120
rect 196360 41120 196520 41280
rect 196360 41280 196520 41440
rect 196360 41440 196520 41600
rect 196360 41600 196520 41760
rect 196360 41760 196520 41920
rect 196360 41920 196520 42080
rect 196360 42080 196520 42240
rect 196360 42240 196520 42400
rect 196360 42400 196520 42560
rect 196360 42560 196520 42720
rect 196360 42720 196520 42880
rect 196360 42880 196520 43040
rect 196360 43040 196520 43200
rect 196360 43200 196520 43360
rect 196360 43360 196520 43520
rect 196360 43520 196520 43680
rect 196360 43680 196520 43840
rect 196360 43840 196520 44000
rect 196360 44000 196520 44160
rect 196360 44160 196520 44320
rect 196360 44320 196520 44480
rect 196360 44480 196520 44640
rect 196360 44640 196520 44800
rect 196360 44800 196520 44960
rect 196360 44960 196520 45120
rect 196360 45120 196520 45280
rect 196360 45280 196520 45440
rect 196360 45440 196520 45600
rect 196520 37280 196680 37440
rect 196520 37440 196680 37600
rect 196520 37600 196680 37760
rect 196520 37760 196680 37920
rect 196520 37920 196680 38080
rect 196520 38080 196680 38240
rect 196520 38240 196680 38400
rect 196520 38400 196680 38560
rect 196520 38560 196680 38720
rect 196520 38720 196680 38880
rect 196520 38880 196680 39040
rect 196520 39040 196680 39200
rect 196520 39200 196680 39360
rect 196520 39360 196680 39520
rect 196520 39520 196680 39680
rect 196520 39680 196680 39840
rect 196520 39840 196680 40000
rect 196520 40000 196680 40160
rect 196520 40160 196680 40320
rect 196520 40320 196680 40480
rect 196520 40480 196680 40640
rect 196520 40640 196680 40800
rect 196520 40800 196680 40960
rect 196520 40960 196680 41120
rect 196520 41120 196680 41280
rect 196520 41280 196680 41440
rect 196520 41440 196680 41600
rect 196520 41600 196680 41760
rect 196520 41760 196680 41920
rect 196520 41920 196680 42080
rect 196520 42080 196680 42240
rect 196520 42240 196680 42400
rect 196520 42400 196680 42560
rect 196520 42560 196680 42720
rect 196520 42720 196680 42880
rect 196520 42880 196680 43040
rect 196520 43040 196680 43200
rect 196520 43200 196680 43360
rect 196520 43360 196680 43520
rect 196520 43520 196680 43680
rect 196520 43680 196680 43840
rect 196520 43840 196680 44000
rect 196520 44000 196680 44160
rect 196520 44160 196680 44320
rect 196520 44320 196680 44480
rect 196520 44480 196680 44640
rect 196520 44640 196680 44800
rect 196520 44800 196680 44960
rect 196520 44960 196680 45120
rect 196520 45120 196680 45280
rect 196520 45280 196680 45440
rect 196520 45440 196680 45600
rect 196520 45600 196680 45760
rect 196520 45760 196680 45920
rect 196520 45920 196680 46080
rect 196680 37760 196840 37920
rect 196680 37920 196840 38080
rect 196680 38080 196840 38240
rect 196680 38240 196840 38400
rect 196680 38400 196840 38560
rect 196680 38560 196840 38720
rect 196680 38720 196840 38880
rect 196680 38880 196840 39040
rect 196680 39040 196840 39200
rect 196680 39200 196840 39360
rect 196680 39360 196840 39520
rect 196680 39520 196840 39680
rect 196680 39680 196840 39840
rect 196680 39840 196840 40000
rect 196680 40000 196840 40160
rect 196680 40160 196840 40320
rect 196680 40320 196840 40480
rect 196680 40480 196840 40640
rect 196680 40640 196840 40800
rect 196680 40800 196840 40960
rect 196680 40960 196840 41120
rect 196680 41120 196840 41280
rect 196680 41280 196840 41440
rect 196680 41440 196840 41600
rect 196680 41600 196840 41760
rect 196680 41760 196840 41920
rect 196680 41920 196840 42080
rect 196680 42080 196840 42240
rect 196680 42240 196840 42400
rect 196680 42400 196840 42560
rect 196680 42560 196840 42720
rect 196680 42720 196840 42880
rect 196680 42880 196840 43040
rect 196680 43040 196840 43200
rect 196680 43200 196840 43360
rect 196680 43360 196840 43520
rect 196680 43520 196840 43680
rect 196680 43680 196840 43840
rect 196680 43840 196840 44000
rect 196680 44000 196840 44160
rect 196680 44160 196840 44320
rect 196680 44320 196840 44480
rect 196680 44480 196840 44640
rect 196680 44640 196840 44800
rect 196680 44800 196840 44960
rect 196680 44960 196840 45120
rect 196680 45120 196840 45280
rect 196680 45280 196840 45440
rect 196680 45440 196840 45600
rect 196680 45600 196840 45760
rect 196680 45760 196840 45920
rect 196680 45920 196840 46080
rect 196680 46080 196840 46240
rect 196680 46240 196840 46400
rect 196680 46400 196840 46560
rect 196680 46560 196840 46720
rect 196840 38080 197000 38240
rect 196840 38240 197000 38400
rect 196840 38400 197000 38560
rect 196840 38560 197000 38720
rect 196840 38720 197000 38880
rect 196840 38880 197000 39040
rect 196840 39040 197000 39200
rect 196840 39200 197000 39360
rect 196840 39360 197000 39520
rect 196840 39520 197000 39680
rect 196840 39680 197000 39840
rect 196840 39840 197000 40000
rect 196840 40000 197000 40160
rect 196840 40160 197000 40320
rect 196840 40320 197000 40480
rect 196840 40480 197000 40640
rect 196840 40640 197000 40800
rect 196840 40800 197000 40960
rect 196840 40960 197000 41120
rect 196840 41120 197000 41280
rect 196840 41280 197000 41440
rect 196840 41440 197000 41600
rect 196840 41600 197000 41760
rect 196840 41760 197000 41920
rect 196840 41920 197000 42080
rect 196840 42080 197000 42240
rect 196840 42240 197000 42400
rect 196840 42400 197000 42560
rect 196840 42560 197000 42720
rect 196840 42720 197000 42880
rect 196840 42880 197000 43040
rect 196840 43040 197000 43200
rect 196840 43200 197000 43360
rect 196840 43360 197000 43520
rect 196840 43520 197000 43680
rect 196840 43680 197000 43840
rect 196840 43840 197000 44000
rect 196840 44000 197000 44160
rect 196840 44160 197000 44320
rect 196840 44320 197000 44480
rect 196840 44480 197000 44640
rect 196840 44640 197000 44800
rect 196840 44800 197000 44960
rect 196840 44960 197000 45120
rect 196840 45120 197000 45280
rect 196840 45280 197000 45440
rect 196840 45440 197000 45600
rect 196840 45600 197000 45760
rect 196840 45760 197000 45920
rect 196840 45920 197000 46080
rect 196840 46080 197000 46240
rect 196840 46240 197000 46400
rect 196840 46400 197000 46560
rect 196840 46560 197000 46720
rect 196840 46720 197000 46880
rect 196840 46880 197000 47040
rect 196840 47040 197000 47200
rect 197000 38560 197160 38720
rect 197000 38720 197160 38880
rect 197000 38880 197160 39040
rect 197000 39040 197160 39200
rect 197000 39200 197160 39360
rect 197000 39360 197160 39520
rect 197000 39520 197160 39680
rect 197000 39680 197160 39840
rect 197000 39840 197160 40000
rect 197000 40000 197160 40160
rect 197000 40160 197160 40320
rect 197000 40320 197160 40480
rect 197000 40480 197160 40640
rect 197000 40640 197160 40800
rect 197000 40800 197160 40960
rect 197000 40960 197160 41120
rect 197000 41120 197160 41280
rect 197000 41280 197160 41440
rect 197000 41440 197160 41600
rect 197000 41600 197160 41760
rect 197000 41760 197160 41920
rect 197000 41920 197160 42080
rect 197000 42080 197160 42240
rect 197000 42240 197160 42400
rect 197000 42400 197160 42560
rect 197000 42560 197160 42720
rect 197000 42720 197160 42880
rect 197000 42880 197160 43040
rect 197000 43040 197160 43200
rect 197000 43200 197160 43360
rect 197000 43360 197160 43520
rect 197000 43520 197160 43680
rect 197000 43680 197160 43840
rect 197000 43840 197160 44000
rect 197000 44000 197160 44160
rect 197000 44160 197160 44320
rect 197000 44320 197160 44480
rect 197000 44480 197160 44640
rect 197000 44640 197160 44800
rect 197000 44800 197160 44960
rect 197000 44960 197160 45120
rect 197000 45120 197160 45280
rect 197000 45280 197160 45440
rect 197000 45440 197160 45600
rect 197000 45600 197160 45760
rect 197000 45760 197160 45920
rect 197000 45920 197160 46080
rect 197000 46080 197160 46240
rect 197000 46240 197160 46400
rect 197000 46400 197160 46560
rect 197000 46560 197160 46720
rect 197000 46720 197160 46880
rect 197000 46880 197160 47040
rect 197000 47040 197160 47200
rect 197000 47200 197160 47360
rect 197000 47360 197160 47520
rect 197000 47520 197160 47680
rect 197000 47680 197160 47840
rect 197160 38880 197320 39040
rect 197160 39040 197320 39200
rect 197160 39200 197320 39360
rect 197160 39360 197320 39520
rect 197160 39520 197320 39680
rect 197160 39680 197320 39840
rect 197160 39840 197320 40000
rect 197160 40000 197320 40160
rect 197160 40160 197320 40320
rect 197160 40320 197320 40480
rect 197160 40480 197320 40640
rect 197160 40640 197320 40800
rect 197160 40800 197320 40960
rect 197160 40960 197320 41120
rect 197160 41120 197320 41280
rect 197160 41280 197320 41440
rect 197160 41440 197320 41600
rect 197160 41600 197320 41760
rect 197160 41760 197320 41920
rect 197160 41920 197320 42080
rect 197160 42080 197320 42240
rect 197160 42240 197320 42400
rect 197160 42400 197320 42560
rect 197160 42560 197320 42720
rect 197160 42720 197320 42880
rect 197160 42880 197320 43040
rect 197160 43040 197320 43200
rect 197160 43200 197320 43360
rect 197160 43360 197320 43520
rect 197160 43520 197320 43680
rect 197160 43680 197320 43840
rect 197160 43840 197320 44000
rect 197160 44000 197320 44160
rect 197160 44160 197320 44320
rect 197160 44320 197320 44480
rect 197160 44480 197320 44640
rect 197160 44640 197320 44800
rect 197160 44800 197320 44960
rect 197160 44960 197320 45120
rect 197160 45120 197320 45280
rect 197160 45280 197320 45440
rect 197160 45440 197320 45600
rect 197160 45600 197320 45760
rect 197160 45760 197320 45920
rect 197160 45920 197320 46080
rect 197160 46080 197320 46240
rect 197160 46240 197320 46400
rect 197160 46400 197320 46560
rect 197160 46560 197320 46720
rect 197160 46720 197320 46880
rect 197160 46880 197320 47040
rect 197160 47040 197320 47200
rect 197160 47200 197320 47360
rect 197160 47360 197320 47520
rect 197160 47520 197320 47680
rect 197160 47680 197320 47840
rect 197160 47840 197320 48000
rect 197160 48000 197320 48160
rect 197160 48160 197320 48320
rect 197160 48320 197320 48480
rect 197320 39360 197480 39520
rect 197320 39520 197480 39680
rect 197320 39680 197480 39840
rect 197320 39840 197480 40000
rect 197320 40000 197480 40160
rect 197320 40160 197480 40320
rect 197320 40320 197480 40480
rect 197320 40480 197480 40640
rect 197320 40640 197480 40800
rect 197320 40800 197480 40960
rect 197320 40960 197480 41120
rect 197320 41120 197480 41280
rect 197320 41280 197480 41440
rect 197320 41440 197480 41600
rect 197320 41600 197480 41760
rect 197320 41760 197480 41920
rect 197320 41920 197480 42080
rect 197320 42080 197480 42240
rect 197320 42240 197480 42400
rect 197320 42400 197480 42560
rect 197320 42560 197480 42720
rect 197320 42720 197480 42880
rect 197320 42880 197480 43040
rect 197320 43040 197480 43200
rect 197320 43200 197480 43360
rect 197320 43360 197480 43520
rect 197320 43520 197480 43680
rect 197320 43680 197480 43840
rect 197320 43840 197480 44000
rect 197320 44000 197480 44160
rect 197320 44160 197480 44320
rect 197320 44320 197480 44480
rect 197320 44480 197480 44640
rect 197320 44640 197480 44800
rect 197320 44800 197480 44960
rect 197320 44960 197480 45120
rect 197320 45120 197480 45280
rect 197320 45280 197480 45440
rect 197320 45440 197480 45600
rect 197320 45600 197480 45760
rect 197320 45760 197480 45920
rect 197320 45920 197480 46080
rect 197320 46080 197480 46240
rect 197320 46240 197480 46400
rect 197320 46400 197480 46560
rect 197320 46560 197480 46720
rect 197320 46720 197480 46880
rect 197320 46880 197480 47040
rect 197320 47040 197480 47200
rect 197320 47200 197480 47360
rect 197320 47360 197480 47520
rect 197320 47520 197480 47680
rect 197320 47680 197480 47840
rect 197320 47840 197480 48000
rect 197320 48000 197480 48160
rect 197320 48160 197480 48320
rect 197320 48320 197480 48480
rect 197320 48480 197480 48640
rect 197320 48640 197480 48800
rect 197320 48800 197480 48960
rect 197320 48960 197480 49120
rect 197480 39680 197640 39840
rect 197480 39840 197640 40000
rect 197480 40000 197640 40160
rect 197480 40160 197640 40320
rect 197480 40320 197640 40480
rect 197480 40480 197640 40640
rect 197480 40640 197640 40800
rect 197480 40800 197640 40960
rect 197480 40960 197640 41120
rect 197480 41120 197640 41280
rect 197480 41280 197640 41440
rect 197480 41440 197640 41600
rect 197480 41600 197640 41760
rect 197480 41760 197640 41920
rect 197480 41920 197640 42080
rect 197480 42080 197640 42240
rect 197480 42240 197640 42400
rect 197480 42400 197640 42560
rect 197480 42560 197640 42720
rect 197480 42720 197640 42880
rect 197480 42880 197640 43040
rect 197480 43040 197640 43200
rect 197480 43200 197640 43360
rect 197480 43360 197640 43520
rect 197480 43520 197640 43680
rect 197480 43680 197640 43840
rect 197480 43840 197640 44000
rect 197480 44000 197640 44160
rect 197480 44160 197640 44320
rect 197480 44320 197640 44480
rect 197480 44480 197640 44640
rect 197480 44640 197640 44800
rect 197480 44800 197640 44960
rect 197480 44960 197640 45120
rect 197480 45120 197640 45280
rect 197480 45280 197640 45440
rect 197480 45440 197640 45600
rect 197480 45600 197640 45760
rect 197480 45760 197640 45920
rect 197480 45920 197640 46080
rect 197480 46080 197640 46240
rect 197480 46240 197640 46400
rect 197480 46400 197640 46560
rect 197480 46560 197640 46720
rect 197480 46720 197640 46880
rect 197480 46880 197640 47040
rect 197480 47040 197640 47200
rect 197480 47200 197640 47360
rect 197480 47360 197640 47520
rect 197480 47520 197640 47680
rect 197480 47680 197640 47840
rect 197480 47840 197640 48000
rect 197480 48000 197640 48160
rect 197480 48160 197640 48320
rect 197480 48320 197640 48480
rect 197480 48480 197640 48640
rect 197480 48640 197640 48800
rect 197480 48800 197640 48960
rect 197480 48960 197640 49120
rect 197480 49120 197640 49280
rect 197480 49280 197640 49440
rect 197480 49440 197640 49600
rect 197480 49600 197640 49760
rect 197640 40000 197800 40160
rect 197640 40160 197800 40320
rect 197640 40320 197800 40480
rect 197640 40480 197800 40640
rect 197640 40640 197800 40800
rect 197640 40800 197800 40960
rect 197640 40960 197800 41120
rect 197640 41120 197800 41280
rect 197640 41280 197800 41440
rect 197640 41440 197800 41600
rect 197640 41600 197800 41760
rect 197640 41760 197800 41920
rect 197640 41920 197800 42080
rect 197640 42080 197800 42240
rect 197640 42240 197800 42400
rect 197640 42400 197800 42560
rect 197640 42560 197800 42720
rect 197640 42720 197800 42880
rect 197640 42880 197800 43040
rect 197640 43040 197800 43200
rect 197640 43200 197800 43360
rect 197640 43360 197800 43520
rect 197640 43520 197800 43680
rect 197640 43680 197800 43840
rect 197640 43840 197800 44000
rect 197640 44000 197800 44160
rect 197640 44160 197800 44320
rect 197640 44320 197800 44480
rect 197640 44480 197800 44640
rect 197640 44640 197800 44800
rect 197640 44800 197800 44960
rect 197640 44960 197800 45120
rect 197640 45120 197800 45280
rect 197640 45280 197800 45440
rect 197640 45440 197800 45600
rect 197640 45600 197800 45760
rect 197640 45760 197800 45920
rect 197640 45920 197800 46080
rect 197640 46080 197800 46240
rect 197640 46240 197800 46400
rect 197640 46400 197800 46560
rect 197640 46560 197800 46720
rect 197640 46720 197800 46880
rect 197640 46880 197800 47040
rect 197640 47040 197800 47200
rect 197640 47200 197800 47360
rect 197640 47360 197800 47520
rect 197640 47520 197800 47680
rect 197640 47680 197800 47840
rect 197640 47840 197800 48000
rect 197640 48000 197800 48160
rect 197640 48160 197800 48320
rect 197640 48320 197800 48480
rect 197640 48480 197800 48640
rect 197640 48640 197800 48800
rect 197640 48800 197800 48960
rect 197640 48960 197800 49120
rect 197640 49120 197800 49280
rect 197640 49280 197800 49440
rect 197640 49440 197800 49600
rect 197640 49600 197800 49760
rect 197640 49760 197800 49920
rect 197640 49920 197800 50080
rect 197640 50080 197800 50240
rect 197800 40480 197960 40640
rect 197800 40640 197960 40800
rect 197800 40800 197960 40960
rect 197800 40960 197960 41120
rect 197800 41120 197960 41280
rect 197800 41280 197960 41440
rect 197800 41440 197960 41600
rect 197800 41600 197960 41760
rect 197800 41760 197960 41920
rect 197800 41920 197960 42080
rect 197800 42080 197960 42240
rect 197800 42240 197960 42400
rect 197800 42400 197960 42560
rect 197800 42560 197960 42720
rect 197800 42720 197960 42880
rect 197800 42880 197960 43040
rect 197800 43040 197960 43200
rect 197800 43200 197960 43360
rect 197800 43360 197960 43520
rect 197800 43520 197960 43680
rect 197800 43680 197960 43840
rect 197800 43840 197960 44000
rect 197800 44000 197960 44160
rect 197800 44160 197960 44320
rect 197800 44320 197960 44480
rect 197800 44480 197960 44640
rect 197800 44640 197960 44800
rect 197800 44800 197960 44960
rect 197800 44960 197960 45120
rect 197800 45120 197960 45280
rect 197800 45280 197960 45440
rect 197800 45440 197960 45600
rect 197800 45600 197960 45760
rect 197800 45760 197960 45920
rect 197800 45920 197960 46080
rect 197800 46080 197960 46240
rect 197800 46240 197960 46400
rect 197800 46400 197960 46560
rect 197800 46560 197960 46720
rect 197800 46720 197960 46880
rect 197800 46880 197960 47040
rect 197800 47040 197960 47200
rect 197800 47200 197960 47360
rect 197800 47360 197960 47520
rect 197800 47520 197960 47680
rect 197800 47680 197960 47840
rect 197800 47840 197960 48000
rect 197800 48000 197960 48160
rect 197800 48160 197960 48320
rect 197800 48320 197960 48480
rect 197800 48480 197960 48640
rect 197800 48640 197960 48800
rect 197800 48800 197960 48960
rect 197800 48960 197960 49120
rect 197800 49120 197960 49280
rect 197800 49280 197960 49440
rect 197800 49440 197960 49600
rect 197800 49600 197960 49760
rect 197800 49760 197960 49920
rect 197800 49920 197960 50080
rect 197800 50080 197960 50240
rect 197800 50240 197960 50400
rect 197800 50400 197960 50560
rect 197800 50560 197960 50720
rect 197960 40800 198120 40960
rect 197960 40960 198120 41120
rect 197960 41120 198120 41280
rect 197960 41280 198120 41440
rect 197960 41440 198120 41600
rect 197960 41600 198120 41760
rect 197960 41760 198120 41920
rect 197960 41920 198120 42080
rect 197960 42080 198120 42240
rect 197960 42240 198120 42400
rect 197960 42400 198120 42560
rect 197960 42560 198120 42720
rect 197960 42720 198120 42880
rect 197960 42880 198120 43040
rect 197960 43040 198120 43200
rect 197960 43200 198120 43360
rect 197960 43360 198120 43520
rect 197960 43520 198120 43680
rect 197960 43680 198120 43840
rect 197960 43840 198120 44000
rect 197960 44000 198120 44160
rect 197960 44160 198120 44320
rect 197960 44320 198120 44480
rect 197960 44480 198120 44640
rect 197960 44640 198120 44800
rect 197960 44800 198120 44960
rect 197960 44960 198120 45120
rect 197960 45120 198120 45280
rect 197960 45280 198120 45440
rect 197960 45440 198120 45600
rect 197960 45600 198120 45760
rect 197960 45760 198120 45920
rect 197960 45920 198120 46080
rect 197960 46080 198120 46240
rect 197960 46240 198120 46400
rect 197960 46400 198120 46560
rect 197960 46560 198120 46720
rect 197960 46720 198120 46880
rect 197960 46880 198120 47040
rect 197960 47040 198120 47200
rect 197960 47200 198120 47360
rect 197960 47360 198120 47520
rect 197960 47520 198120 47680
rect 197960 47680 198120 47840
rect 197960 47840 198120 48000
rect 197960 48000 198120 48160
rect 197960 48160 198120 48320
rect 197960 48320 198120 48480
rect 197960 48480 198120 48640
rect 197960 48640 198120 48800
rect 197960 48800 198120 48960
rect 197960 48960 198120 49120
rect 197960 49120 198120 49280
rect 197960 49280 198120 49440
rect 197960 49440 198120 49600
rect 197960 49600 198120 49760
rect 197960 49760 198120 49920
rect 197960 49920 198120 50080
rect 197960 50080 198120 50240
rect 197960 50240 198120 50400
rect 197960 50400 198120 50560
rect 197960 50560 198120 50720
rect 197960 50720 198120 50880
rect 197960 50880 198120 51040
rect 197960 51040 198120 51200
rect 198120 41280 198280 41440
rect 198120 41440 198280 41600
rect 198120 41600 198280 41760
rect 198120 41760 198280 41920
rect 198120 41920 198280 42080
rect 198120 42080 198280 42240
rect 198120 42240 198280 42400
rect 198120 42400 198280 42560
rect 198120 42560 198280 42720
rect 198120 42720 198280 42880
rect 198120 42880 198280 43040
rect 198120 43040 198280 43200
rect 198120 43200 198280 43360
rect 198120 43360 198280 43520
rect 198120 43520 198280 43680
rect 198120 43680 198280 43840
rect 198120 43840 198280 44000
rect 198120 44000 198280 44160
rect 198120 44160 198280 44320
rect 198120 44320 198280 44480
rect 198120 44480 198280 44640
rect 198120 44640 198280 44800
rect 198120 44800 198280 44960
rect 198120 44960 198280 45120
rect 198120 45120 198280 45280
rect 198120 45280 198280 45440
rect 198120 45440 198280 45600
rect 198120 45600 198280 45760
rect 198120 45760 198280 45920
rect 198120 45920 198280 46080
rect 198120 46080 198280 46240
rect 198120 46240 198280 46400
rect 198120 46400 198280 46560
rect 198120 46560 198280 46720
rect 198120 46720 198280 46880
rect 198120 46880 198280 47040
rect 198120 47040 198280 47200
rect 198120 47200 198280 47360
rect 198120 47360 198280 47520
rect 198120 47520 198280 47680
rect 198120 47680 198280 47840
rect 198120 47840 198280 48000
rect 198120 48000 198280 48160
rect 198120 48160 198280 48320
rect 198120 48320 198280 48480
rect 198120 48480 198280 48640
rect 198120 48640 198280 48800
rect 198120 48800 198280 48960
rect 198120 48960 198280 49120
rect 198120 49120 198280 49280
rect 198120 49280 198280 49440
rect 198120 49440 198280 49600
rect 198120 49600 198280 49760
rect 198120 49760 198280 49920
rect 198120 49920 198280 50080
rect 198120 50080 198280 50240
rect 198120 50240 198280 50400
rect 198120 50400 198280 50560
rect 198120 50560 198280 50720
rect 198120 50720 198280 50880
rect 198120 50880 198280 51040
rect 198120 51040 198280 51200
rect 198120 51200 198280 51360
rect 198120 51360 198280 51520
rect 198280 41600 198440 41760
rect 198280 41760 198440 41920
rect 198280 41920 198440 42080
rect 198280 42080 198440 42240
rect 198280 42240 198440 42400
rect 198280 42400 198440 42560
rect 198280 42560 198440 42720
rect 198280 42720 198440 42880
rect 198280 42880 198440 43040
rect 198280 43040 198440 43200
rect 198280 43200 198440 43360
rect 198280 43360 198440 43520
rect 198280 43520 198440 43680
rect 198280 43680 198440 43840
rect 198280 43840 198440 44000
rect 198280 44000 198440 44160
rect 198280 44160 198440 44320
rect 198280 44320 198440 44480
rect 198280 44480 198440 44640
rect 198280 44640 198440 44800
rect 198280 44800 198440 44960
rect 198280 44960 198440 45120
rect 198280 45120 198440 45280
rect 198280 45280 198440 45440
rect 198280 45440 198440 45600
rect 198280 45600 198440 45760
rect 198280 45760 198440 45920
rect 198280 45920 198440 46080
rect 198280 46080 198440 46240
rect 198280 46240 198440 46400
rect 198280 46400 198440 46560
rect 198280 46560 198440 46720
rect 198280 46720 198440 46880
rect 198280 46880 198440 47040
rect 198280 47040 198440 47200
rect 198280 47200 198440 47360
rect 198280 47360 198440 47520
rect 198280 47520 198440 47680
rect 198280 47680 198440 47840
rect 198280 47840 198440 48000
rect 198280 48000 198440 48160
rect 198280 48160 198440 48320
rect 198280 48320 198440 48480
rect 198280 48480 198440 48640
rect 198280 48640 198440 48800
rect 198280 48800 198440 48960
rect 198280 48960 198440 49120
rect 198280 49120 198440 49280
rect 198280 49280 198440 49440
rect 198280 49440 198440 49600
rect 198280 49600 198440 49760
rect 198280 49760 198440 49920
rect 198280 49920 198440 50080
rect 198280 50080 198440 50240
rect 198280 50240 198440 50400
rect 198280 50400 198440 50560
rect 198280 50560 198440 50720
rect 198280 50720 198440 50880
rect 198280 50880 198440 51040
rect 198280 51040 198440 51200
rect 198280 51200 198440 51360
rect 198280 51360 198440 51520
rect 198280 51520 198440 51680
rect 198280 51680 198440 51840
rect 198440 42080 198600 42240
rect 198440 42240 198600 42400
rect 198440 42400 198600 42560
rect 198440 42560 198600 42720
rect 198440 42720 198600 42880
rect 198440 42880 198600 43040
rect 198440 43040 198600 43200
rect 198440 43200 198600 43360
rect 198440 43360 198600 43520
rect 198440 43520 198600 43680
rect 198440 43680 198600 43840
rect 198440 43840 198600 44000
rect 198440 44000 198600 44160
rect 198440 44160 198600 44320
rect 198440 44320 198600 44480
rect 198440 44480 198600 44640
rect 198440 44640 198600 44800
rect 198440 44800 198600 44960
rect 198440 44960 198600 45120
rect 198440 45120 198600 45280
rect 198440 45280 198600 45440
rect 198440 45440 198600 45600
rect 198440 45600 198600 45760
rect 198440 45760 198600 45920
rect 198440 45920 198600 46080
rect 198440 46080 198600 46240
rect 198440 46240 198600 46400
rect 198440 46400 198600 46560
rect 198440 46560 198600 46720
rect 198440 46720 198600 46880
rect 198440 46880 198600 47040
rect 198440 47040 198600 47200
rect 198440 47200 198600 47360
rect 198440 47360 198600 47520
rect 198440 47520 198600 47680
rect 198440 47680 198600 47840
rect 198440 47840 198600 48000
rect 198440 48000 198600 48160
rect 198440 48160 198600 48320
rect 198440 48320 198600 48480
rect 198440 48480 198600 48640
rect 198440 48640 198600 48800
rect 198440 48800 198600 48960
rect 198440 48960 198600 49120
rect 198440 49120 198600 49280
rect 198440 49280 198600 49440
rect 198440 49440 198600 49600
rect 198440 49600 198600 49760
rect 198440 49760 198600 49920
rect 198440 49920 198600 50080
rect 198440 50080 198600 50240
rect 198440 50240 198600 50400
rect 198440 50400 198600 50560
rect 198440 50560 198600 50720
rect 198440 50720 198600 50880
rect 198440 50880 198600 51040
rect 198440 51040 198600 51200
rect 198440 51200 198600 51360
rect 198440 51360 198600 51520
rect 198440 51520 198600 51680
rect 198440 51680 198600 51840
rect 198440 51840 198600 52000
rect 198440 52000 198600 52160
rect 198600 42400 198760 42560
rect 198600 42560 198760 42720
rect 198600 42720 198760 42880
rect 198600 42880 198760 43040
rect 198600 43040 198760 43200
rect 198600 43200 198760 43360
rect 198600 43360 198760 43520
rect 198600 43520 198760 43680
rect 198600 43680 198760 43840
rect 198600 43840 198760 44000
rect 198600 44000 198760 44160
rect 198600 44160 198760 44320
rect 198600 44320 198760 44480
rect 198600 44480 198760 44640
rect 198600 44640 198760 44800
rect 198600 44800 198760 44960
rect 198600 44960 198760 45120
rect 198600 45120 198760 45280
rect 198600 45280 198760 45440
rect 198600 45440 198760 45600
rect 198600 45600 198760 45760
rect 198600 45760 198760 45920
rect 198600 45920 198760 46080
rect 198600 46080 198760 46240
rect 198600 46240 198760 46400
rect 198600 46400 198760 46560
rect 198600 46560 198760 46720
rect 198600 46720 198760 46880
rect 198600 46880 198760 47040
rect 198600 47040 198760 47200
rect 198600 47200 198760 47360
rect 198600 47360 198760 47520
rect 198600 47520 198760 47680
rect 198600 47680 198760 47840
rect 198600 47840 198760 48000
rect 198600 48000 198760 48160
rect 198600 48160 198760 48320
rect 198600 48320 198760 48480
rect 198600 48480 198760 48640
rect 198600 48640 198760 48800
rect 198600 48800 198760 48960
rect 198600 48960 198760 49120
rect 198600 49120 198760 49280
rect 198600 49280 198760 49440
rect 198600 49440 198760 49600
rect 198600 49600 198760 49760
rect 198600 49760 198760 49920
rect 198600 49920 198760 50080
rect 198600 50080 198760 50240
rect 198600 50240 198760 50400
rect 198600 50400 198760 50560
rect 198600 50560 198760 50720
rect 198600 50720 198760 50880
rect 198600 50880 198760 51040
rect 198600 51040 198760 51200
rect 198600 51200 198760 51360
rect 198600 51360 198760 51520
rect 198600 51520 198760 51680
rect 198600 51680 198760 51840
rect 198600 51840 198760 52000
rect 198600 52000 198760 52160
rect 198600 52160 198760 52320
rect 198760 42720 198920 42880
rect 198760 42880 198920 43040
rect 198760 43040 198920 43200
rect 198760 43200 198920 43360
rect 198760 43360 198920 43520
rect 198760 43520 198920 43680
rect 198760 43680 198920 43840
rect 198760 43840 198920 44000
rect 198760 44000 198920 44160
rect 198760 44160 198920 44320
rect 198760 44320 198920 44480
rect 198760 44480 198920 44640
rect 198760 44640 198920 44800
rect 198760 44800 198920 44960
rect 198760 44960 198920 45120
rect 198760 45120 198920 45280
rect 198760 45280 198920 45440
rect 198760 45440 198920 45600
rect 198760 45600 198920 45760
rect 198760 45760 198920 45920
rect 198760 45920 198920 46080
rect 198760 46080 198920 46240
rect 198760 46240 198920 46400
rect 198760 46400 198920 46560
rect 198760 46560 198920 46720
rect 198760 46720 198920 46880
rect 198760 46880 198920 47040
rect 198760 47040 198920 47200
rect 198760 47200 198920 47360
rect 198760 47360 198920 47520
rect 198760 47520 198920 47680
rect 198760 47680 198920 47840
rect 198760 47840 198920 48000
rect 198760 48000 198920 48160
rect 198760 48160 198920 48320
rect 198760 48320 198920 48480
rect 198760 48480 198920 48640
rect 198760 48640 198920 48800
rect 198760 48800 198920 48960
rect 198760 48960 198920 49120
rect 198760 49120 198920 49280
rect 198760 49280 198920 49440
rect 198760 49440 198920 49600
rect 198760 49600 198920 49760
rect 198760 49760 198920 49920
rect 198760 49920 198920 50080
rect 198760 50080 198920 50240
rect 198760 50240 198920 50400
rect 198760 50400 198920 50560
rect 198760 50560 198920 50720
rect 198760 50720 198920 50880
rect 198760 50880 198920 51040
rect 198760 51040 198920 51200
rect 198760 51200 198920 51360
rect 198760 51360 198920 51520
rect 198760 51520 198920 51680
rect 198760 51680 198920 51840
rect 198760 51840 198920 52000
rect 198760 52000 198920 52160
rect 198760 52160 198920 52320
rect 198760 52320 198920 52480
rect 198760 52480 198920 52640
rect 198920 43200 199080 43360
rect 198920 43360 199080 43520
rect 198920 43520 199080 43680
rect 198920 43680 199080 43840
rect 198920 43840 199080 44000
rect 198920 44000 199080 44160
rect 198920 44160 199080 44320
rect 198920 44320 199080 44480
rect 198920 44480 199080 44640
rect 198920 44640 199080 44800
rect 198920 44800 199080 44960
rect 198920 44960 199080 45120
rect 198920 45120 199080 45280
rect 198920 45280 199080 45440
rect 198920 45440 199080 45600
rect 198920 45600 199080 45760
rect 198920 45760 199080 45920
rect 198920 45920 199080 46080
rect 198920 46080 199080 46240
rect 198920 46240 199080 46400
rect 198920 46400 199080 46560
rect 198920 46560 199080 46720
rect 198920 46720 199080 46880
rect 198920 46880 199080 47040
rect 198920 47040 199080 47200
rect 198920 47200 199080 47360
rect 198920 47360 199080 47520
rect 198920 47520 199080 47680
rect 198920 47680 199080 47840
rect 198920 47840 199080 48000
rect 198920 48000 199080 48160
rect 198920 48160 199080 48320
rect 198920 48320 199080 48480
rect 198920 48480 199080 48640
rect 198920 48640 199080 48800
rect 198920 48800 199080 48960
rect 198920 48960 199080 49120
rect 198920 49120 199080 49280
rect 198920 49280 199080 49440
rect 198920 49440 199080 49600
rect 198920 49600 199080 49760
rect 198920 49760 199080 49920
rect 198920 49920 199080 50080
rect 198920 50080 199080 50240
rect 198920 50240 199080 50400
rect 198920 50400 199080 50560
rect 198920 50560 199080 50720
rect 198920 50720 199080 50880
rect 198920 50880 199080 51040
rect 198920 51040 199080 51200
rect 198920 51200 199080 51360
rect 198920 51360 199080 51520
rect 198920 51520 199080 51680
rect 198920 51680 199080 51840
rect 198920 51840 199080 52000
rect 198920 52000 199080 52160
rect 198920 52160 199080 52320
rect 198920 52320 199080 52480
rect 198920 52480 199080 52640
rect 198920 52640 199080 52800
rect 199080 43520 199240 43680
rect 199080 43680 199240 43840
rect 199080 43840 199240 44000
rect 199080 44000 199240 44160
rect 199080 44160 199240 44320
rect 199080 44320 199240 44480
rect 199080 44480 199240 44640
rect 199080 44640 199240 44800
rect 199080 44800 199240 44960
rect 199080 44960 199240 45120
rect 199080 45120 199240 45280
rect 199080 45280 199240 45440
rect 199080 45440 199240 45600
rect 199080 45600 199240 45760
rect 199080 45760 199240 45920
rect 199080 45920 199240 46080
rect 199080 46080 199240 46240
rect 199080 46240 199240 46400
rect 199080 46400 199240 46560
rect 199080 46560 199240 46720
rect 199080 46720 199240 46880
rect 199080 46880 199240 47040
rect 199080 47040 199240 47200
rect 199080 47200 199240 47360
rect 199080 47360 199240 47520
rect 199080 47520 199240 47680
rect 199080 47680 199240 47840
rect 199080 47840 199240 48000
rect 199080 48000 199240 48160
rect 199080 48160 199240 48320
rect 199080 48320 199240 48480
rect 199080 48480 199240 48640
rect 199080 48640 199240 48800
rect 199080 48800 199240 48960
rect 199080 48960 199240 49120
rect 199080 49120 199240 49280
rect 199080 49280 199240 49440
rect 199080 49440 199240 49600
rect 199080 49600 199240 49760
rect 199080 49760 199240 49920
rect 199080 49920 199240 50080
rect 199080 50080 199240 50240
rect 199080 50240 199240 50400
rect 199080 50400 199240 50560
rect 199080 50560 199240 50720
rect 199080 50720 199240 50880
rect 199080 50880 199240 51040
rect 199080 51040 199240 51200
rect 199080 51200 199240 51360
rect 199080 51360 199240 51520
rect 199080 51520 199240 51680
rect 199080 51680 199240 51840
rect 199080 51840 199240 52000
rect 199080 52000 199240 52160
rect 199080 52160 199240 52320
rect 199080 52320 199240 52480
rect 199080 52480 199240 52640
rect 199080 52640 199240 52800
rect 199080 52800 199240 52960
rect 199240 44000 199400 44160
rect 199240 44160 199400 44320
rect 199240 44320 199400 44480
rect 199240 44480 199400 44640
rect 199240 44640 199400 44800
rect 199240 44800 199400 44960
rect 199240 44960 199400 45120
rect 199240 45120 199400 45280
rect 199240 45280 199400 45440
rect 199240 45440 199400 45600
rect 199240 45600 199400 45760
rect 199240 45760 199400 45920
rect 199240 45920 199400 46080
rect 199240 46080 199400 46240
rect 199240 46240 199400 46400
rect 199240 46400 199400 46560
rect 199240 46560 199400 46720
rect 199240 46720 199400 46880
rect 199240 46880 199400 47040
rect 199240 47040 199400 47200
rect 199240 47200 199400 47360
rect 199240 47360 199400 47520
rect 199240 47520 199400 47680
rect 199240 47680 199400 47840
rect 199240 47840 199400 48000
rect 199240 48000 199400 48160
rect 199240 48160 199400 48320
rect 199240 48320 199400 48480
rect 199240 48480 199400 48640
rect 199240 48640 199400 48800
rect 199240 48800 199400 48960
rect 199240 48960 199400 49120
rect 199240 49120 199400 49280
rect 199240 49280 199400 49440
rect 199240 49440 199400 49600
rect 199240 49600 199400 49760
rect 199240 49760 199400 49920
rect 199240 49920 199400 50080
rect 199240 50080 199400 50240
rect 199240 50240 199400 50400
rect 199240 50400 199400 50560
rect 199240 50560 199400 50720
rect 199240 50720 199400 50880
rect 199240 50880 199400 51040
rect 199240 51040 199400 51200
rect 199240 51200 199400 51360
rect 199240 51360 199400 51520
rect 199240 51520 199400 51680
rect 199240 51680 199400 51840
rect 199240 51840 199400 52000
rect 199240 52000 199400 52160
rect 199240 52160 199400 52320
rect 199240 52320 199400 52480
rect 199240 52480 199400 52640
rect 199240 52640 199400 52800
rect 199240 52800 199400 52960
rect 199400 44320 199560 44480
rect 199400 44480 199560 44640
rect 199400 44640 199560 44800
rect 199400 44800 199560 44960
rect 199400 44960 199560 45120
rect 199400 45120 199560 45280
rect 199400 45280 199560 45440
rect 199400 45440 199560 45600
rect 199400 45600 199560 45760
rect 199400 45760 199560 45920
rect 199400 45920 199560 46080
rect 199400 46080 199560 46240
rect 199400 46240 199560 46400
rect 199400 46400 199560 46560
rect 199400 46560 199560 46720
rect 199400 46720 199560 46880
rect 199400 46880 199560 47040
rect 199400 47040 199560 47200
rect 199400 47200 199560 47360
rect 199400 47360 199560 47520
rect 199400 47520 199560 47680
rect 199400 47680 199560 47840
rect 199400 47840 199560 48000
rect 199400 48000 199560 48160
rect 199400 48160 199560 48320
rect 199400 48320 199560 48480
rect 199400 48480 199560 48640
rect 199400 48640 199560 48800
rect 199400 48800 199560 48960
rect 199400 48960 199560 49120
rect 199400 49120 199560 49280
rect 199400 49280 199560 49440
rect 199400 49440 199560 49600
rect 199400 49600 199560 49760
rect 199400 49760 199560 49920
rect 199400 49920 199560 50080
rect 199400 50080 199560 50240
rect 199400 50240 199560 50400
rect 199400 50400 199560 50560
rect 199400 50560 199560 50720
rect 199400 50720 199560 50880
rect 199400 50880 199560 51040
rect 199400 51040 199560 51200
rect 199400 51200 199560 51360
rect 199400 51360 199560 51520
rect 199400 51520 199560 51680
rect 199400 51680 199560 51840
rect 199400 51840 199560 52000
rect 199400 52000 199560 52160
rect 199400 52160 199560 52320
rect 199400 52320 199560 52480
rect 199400 52480 199560 52640
rect 199400 52640 199560 52800
rect 199400 52800 199560 52960
rect 199400 52960 199560 53120
rect 199560 44800 199720 44960
rect 199560 44960 199720 45120
rect 199560 45120 199720 45280
rect 199560 45280 199720 45440
rect 199560 45440 199720 45600
rect 199560 45600 199720 45760
rect 199560 45760 199720 45920
rect 199560 45920 199720 46080
rect 199560 46080 199720 46240
rect 199560 46240 199720 46400
rect 199560 46400 199720 46560
rect 199560 46560 199720 46720
rect 199560 46720 199720 46880
rect 199560 46880 199720 47040
rect 199560 47040 199720 47200
rect 199560 47200 199720 47360
rect 199560 47360 199720 47520
rect 199560 47520 199720 47680
rect 199560 47680 199720 47840
rect 199560 47840 199720 48000
rect 199560 48000 199720 48160
rect 199560 48160 199720 48320
rect 199560 48320 199720 48480
rect 199560 48480 199720 48640
rect 199560 48640 199720 48800
rect 199560 48800 199720 48960
rect 199560 48960 199720 49120
rect 199560 49120 199720 49280
rect 199560 49280 199720 49440
rect 199560 49440 199720 49600
rect 199560 49600 199720 49760
rect 199560 49760 199720 49920
rect 199560 49920 199720 50080
rect 199560 50080 199720 50240
rect 199560 50240 199720 50400
rect 199560 50400 199720 50560
rect 199560 50560 199720 50720
rect 199560 50720 199720 50880
rect 199560 50880 199720 51040
rect 199560 51040 199720 51200
rect 199560 51200 199720 51360
rect 199560 51360 199720 51520
rect 199560 51520 199720 51680
rect 199560 51680 199720 51840
rect 199560 51840 199720 52000
rect 199560 52000 199720 52160
rect 199560 52160 199720 52320
rect 199560 52320 199720 52480
rect 199560 52480 199720 52640
rect 199560 52640 199720 52800
rect 199560 52800 199720 52960
rect 199560 52960 199720 53120
rect 199720 45120 199880 45280
rect 199720 45280 199880 45440
rect 199720 45440 199880 45600
rect 199720 45600 199880 45760
rect 199720 45760 199880 45920
rect 199720 45920 199880 46080
rect 199720 46080 199880 46240
rect 199720 46240 199880 46400
rect 199720 46400 199880 46560
rect 199720 46560 199880 46720
rect 199720 46720 199880 46880
rect 199720 46880 199880 47040
rect 199720 47040 199880 47200
rect 199720 47200 199880 47360
rect 199720 47360 199880 47520
rect 199720 47520 199880 47680
rect 199720 47680 199880 47840
rect 199720 47840 199880 48000
rect 199720 48000 199880 48160
rect 199720 48160 199880 48320
rect 199720 48320 199880 48480
rect 199720 48480 199880 48640
rect 199720 48640 199880 48800
rect 199720 48800 199880 48960
rect 199720 48960 199880 49120
rect 199720 49120 199880 49280
rect 199720 49280 199880 49440
rect 199720 49440 199880 49600
rect 199720 49600 199880 49760
rect 199720 49760 199880 49920
rect 199720 49920 199880 50080
rect 199720 50080 199880 50240
rect 199720 50240 199880 50400
rect 199720 50400 199880 50560
rect 199720 50560 199880 50720
rect 199720 50720 199880 50880
rect 199720 50880 199880 51040
rect 199720 51040 199880 51200
rect 199720 51200 199880 51360
rect 199720 51360 199880 51520
rect 199720 51520 199880 51680
rect 199720 51680 199880 51840
rect 199720 51840 199880 52000
rect 199720 52000 199880 52160
rect 199720 52160 199880 52320
rect 199720 52320 199880 52480
rect 199720 52480 199880 52640
rect 199720 52640 199880 52800
rect 199720 52800 199880 52960
rect 199720 52960 199880 53120
rect 199720 53120 199880 53280
rect 199880 45600 200040 45760
rect 199880 45760 200040 45920
rect 199880 45920 200040 46080
rect 199880 46080 200040 46240
rect 199880 46240 200040 46400
rect 199880 46400 200040 46560
rect 199880 46560 200040 46720
rect 199880 46720 200040 46880
rect 199880 46880 200040 47040
rect 199880 47040 200040 47200
rect 199880 47200 200040 47360
rect 199880 47360 200040 47520
rect 199880 47520 200040 47680
rect 199880 47680 200040 47840
rect 199880 47840 200040 48000
rect 199880 48000 200040 48160
rect 199880 48160 200040 48320
rect 199880 48320 200040 48480
rect 199880 48480 200040 48640
rect 199880 48640 200040 48800
rect 199880 48800 200040 48960
rect 199880 48960 200040 49120
rect 199880 49120 200040 49280
rect 199880 49280 200040 49440
rect 199880 49440 200040 49600
rect 199880 49600 200040 49760
rect 199880 49760 200040 49920
rect 199880 49920 200040 50080
rect 199880 50080 200040 50240
rect 199880 50240 200040 50400
rect 199880 50400 200040 50560
rect 199880 50560 200040 50720
rect 199880 50720 200040 50880
rect 199880 50880 200040 51040
rect 199880 51040 200040 51200
rect 199880 51200 200040 51360
rect 199880 51360 200040 51520
rect 199880 51520 200040 51680
rect 199880 51680 200040 51840
rect 199880 51840 200040 52000
rect 199880 52000 200040 52160
rect 199880 52160 200040 52320
rect 199880 52320 200040 52480
rect 199880 52480 200040 52640
rect 199880 52640 200040 52800
rect 199880 52800 200040 52960
rect 199880 52960 200040 53120
rect 199880 53120 200040 53280
rect 200040 46080 200200 46240
rect 200040 46240 200200 46400
rect 200040 46400 200200 46560
rect 200040 46560 200200 46720
rect 200040 46720 200200 46880
rect 200040 46880 200200 47040
rect 200040 47040 200200 47200
rect 200040 47200 200200 47360
rect 200040 47360 200200 47520
rect 200040 47520 200200 47680
rect 200040 47680 200200 47840
rect 200040 47840 200200 48000
rect 200040 48000 200200 48160
rect 200040 48160 200200 48320
rect 200040 48320 200200 48480
rect 200040 48480 200200 48640
rect 200040 48640 200200 48800
rect 200040 48800 200200 48960
rect 200040 48960 200200 49120
rect 200040 49120 200200 49280
rect 200040 49280 200200 49440
rect 200040 49440 200200 49600
rect 200040 49600 200200 49760
rect 200040 49760 200200 49920
rect 200040 49920 200200 50080
rect 200040 50080 200200 50240
rect 200040 50240 200200 50400
rect 200040 50400 200200 50560
rect 200040 50560 200200 50720
rect 200040 50720 200200 50880
rect 200040 50880 200200 51040
rect 200040 51040 200200 51200
rect 200040 51200 200200 51360
rect 200040 51360 200200 51520
rect 200040 51520 200200 51680
rect 200040 51680 200200 51840
rect 200040 51840 200200 52000
rect 200040 52000 200200 52160
rect 200040 52160 200200 52320
rect 200040 52320 200200 52480
rect 200040 52480 200200 52640
rect 200040 52640 200200 52800
rect 200040 52800 200200 52960
rect 200040 52960 200200 53120
rect 200040 53120 200200 53280
rect 200200 46720 200360 46880
rect 200200 46880 200360 47040
rect 200200 47040 200360 47200
rect 200200 47200 200360 47360
rect 200200 47360 200360 47520
rect 200200 47520 200360 47680
rect 200200 47680 200360 47840
rect 200200 47840 200360 48000
rect 200200 48000 200360 48160
rect 200200 48160 200360 48320
rect 200200 48320 200360 48480
rect 200200 48480 200360 48640
rect 200200 48640 200360 48800
rect 200200 48800 200360 48960
rect 200200 48960 200360 49120
rect 200200 49120 200360 49280
rect 200200 49280 200360 49440
rect 200200 49440 200360 49600
rect 200200 49600 200360 49760
rect 200200 49760 200360 49920
rect 200200 49920 200360 50080
rect 200200 50080 200360 50240
rect 200200 50240 200360 50400
rect 200200 50400 200360 50560
rect 200200 50560 200360 50720
rect 200200 50720 200360 50880
rect 200200 50880 200360 51040
rect 200200 51040 200360 51200
rect 200200 51200 200360 51360
rect 200200 51360 200360 51520
rect 200200 51520 200360 51680
rect 200200 51680 200360 51840
rect 200200 51840 200360 52000
rect 200200 52000 200360 52160
rect 200200 52160 200360 52320
rect 200200 52320 200360 52480
rect 200200 52480 200360 52640
rect 200200 52640 200360 52800
rect 200200 52800 200360 52960
rect 200200 52960 200360 53120
rect 200200 53120 200360 53280
rect 200360 47200 200520 47360
rect 200360 47360 200520 47520
rect 200360 47520 200520 47680
rect 200360 47680 200520 47840
rect 200360 47840 200520 48000
rect 200360 48000 200520 48160
rect 200360 48160 200520 48320
rect 200360 48320 200520 48480
rect 200360 48480 200520 48640
rect 200360 48640 200520 48800
rect 200360 48800 200520 48960
rect 200360 48960 200520 49120
rect 200360 49120 200520 49280
rect 200360 49280 200520 49440
rect 200360 49440 200520 49600
rect 200360 49600 200520 49760
rect 200360 49760 200520 49920
rect 200360 49920 200520 50080
rect 200360 50080 200520 50240
rect 200360 50240 200520 50400
rect 200360 50400 200520 50560
rect 200360 50560 200520 50720
rect 200360 50720 200520 50880
rect 200360 50880 200520 51040
rect 200360 51040 200520 51200
rect 200360 51200 200520 51360
rect 200360 51360 200520 51520
rect 200360 51520 200520 51680
rect 200360 51680 200520 51840
rect 200360 51840 200520 52000
rect 200360 52000 200520 52160
rect 200360 52160 200520 52320
rect 200360 52320 200520 52480
rect 200360 52480 200520 52640
rect 200360 52640 200520 52800
rect 200360 52800 200520 52960
rect 200360 52960 200520 53120
rect 200360 53120 200520 53280
rect 200520 47680 200680 47840
rect 200520 47840 200680 48000
rect 200520 48000 200680 48160
rect 200520 48160 200680 48320
rect 200520 48320 200680 48480
rect 200520 48480 200680 48640
rect 200520 48640 200680 48800
rect 200520 48800 200680 48960
rect 200520 48960 200680 49120
rect 200520 49120 200680 49280
rect 200520 49280 200680 49440
rect 200520 49440 200680 49600
rect 200520 49600 200680 49760
rect 200520 49760 200680 49920
rect 200520 49920 200680 50080
rect 200520 50080 200680 50240
rect 200520 50240 200680 50400
rect 200520 50400 200680 50560
rect 200520 50560 200680 50720
rect 200520 50720 200680 50880
rect 200520 50880 200680 51040
rect 200520 51040 200680 51200
rect 200520 51200 200680 51360
rect 200520 51360 200680 51520
rect 200520 51520 200680 51680
rect 200520 51680 200680 51840
rect 200520 51840 200680 52000
rect 200520 52000 200680 52160
rect 200520 52160 200680 52320
rect 200520 52320 200680 52480
rect 200520 52480 200680 52640
rect 200520 52640 200680 52800
rect 200520 52800 200680 52960
rect 200520 52960 200680 53120
rect 200520 53120 200680 53280
rect 200680 48160 200840 48320
rect 200680 48320 200840 48480
rect 200680 48480 200840 48640
rect 200680 48640 200840 48800
rect 200680 48800 200840 48960
rect 200680 48960 200840 49120
rect 200680 49120 200840 49280
rect 200680 49280 200840 49440
rect 200680 49440 200840 49600
rect 200680 49600 200840 49760
rect 200680 49760 200840 49920
rect 200680 49920 200840 50080
rect 200680 50080 200840 50240
rect 200680 50240 200840 50400
rect 200680 50400 200840 50560
rect 200680 50560 200840 50720
rect 200680 50720 200840 50880
rect 200680 50880 200840 51040
rect 200680 51040 200840 51200
rect 200680 51200 200840 51360
rect 200680 51360 200840 51520
rect 200680 51520 200840 51680
rect 200680 51680 200840 51840
rect 200680 51840 200840 52000
rect 200680 52000 200840 52160
rect 200680 52160 200840 52320
rect 200680 52320 200840 52480
rect 200680 52480 200840 52640
rect 200680 52640 200840 52800
rect 200680 52800 200840 52960
rect 200680 52960 200840 53120
rect 200680 53120 200840 53280
rect 200840 48640 201000 48800
rect 200840 48800 201000 48960
rect 200840 48960 201000 49120
rect 200840 49120 201000 49280
rect 200840 49280 201000 49440
rect 200840 49440 201000 49600
rect 200840 49600 201000 49760
rect 200840 49760 201000 49920
rect 200840 49920 201000 50080
rect 200840 50080 201000 50240
rect 200840 50240 201000 50400
rect 200840 50400 201000 50560
rect 200840 50560 201000 50720
rect 200840 50720 201000 50880
rect 200840 50880 201000 51040
rect 200840 51040 201000 51200
rect 200840 51200 201000 51360
rect 200840 51360 201000 51520
rect 200840 51520 201000 51680
rect 200840 51680 201000 51840
rect 200840 51840 201000 52000
rect 200840 52000 201000 52160
rect 200840 52160 201000 52320
rect 200840 52320 201000 52480
rect 200840 52480 201000 52640
rect 200840 52640 201000 52800
rect 200840 52800 201000 52960
rect 200840 52960 201000 53120
rect 201000 49120 201160 49280
rect 201000 49280 201160 49440
rect 201000 49440 201160 49600
rect 201000 49600 201160 49760
rect 201000 49760 201160 49920
rect 201000 49920 201160 50080
rect 201000 50080 201160 50240
rect 201000 50240 201160 50400
rect 201000 50400 201160 50560
rect 201000 50560 201160 50720
rect 201000 50720 201160 50880
rect 201000 50880 201160 51040
rect 201000 51040 201160 51200
rect 201000 51200 201160 51360
rect 201000 51360 201160 51520
rect 201000 51520 201160 51680
rect 201000 51680 201160 51840
rect 201000 51840 201160 52000
rect 201000 52000 201160 52160
rect 201000 52160 201160 52320
rect 201000 52320 201160 52480
rect 201000 52480 201160 52640
rect 201000 52640 201160 52800
rect 201000 52800 201160 52960
rect 201000 52960 201160 53120
rect 201160 49440 201320 49600
rect 201160 49600 201320 49760
rect 201160 49760 201320 49920
rect 201160 49920 201320 50080
rect 201160 50080 201320 50240
rect 201160 50240 201320 50400
rect 201160 50400 201320 50560
rect 201160 50560 201320 50720
rect 201160 50720 201320 50880
rect 201160 50880 201320 51040
rect 201160 51040 201320 51200
rect 201160 51200 201320 51360
rect 201160 51360 201320 51520
rect 201160 51520 201320 51680
rect 201160 51680 201320 51840
rect 201160 51840 201320 52000
rect 201160 52000 201320 52160
rect 201160 52160 201320 52320
rect 201160 52320 201320 52480
rect 201160 52480 201320 52640
rect 201160 52640 201320 52800
rect 201160 52800 201320 52960
rect 201160 52960 201320 53120
rect 201320 49920 201480 50080
rect 201320 50080 201480 50240
rect 201320 50240 201480 50400
rect 201320 50400 201480 50560
rect 201320 50560 201480 50720
rect 201320 50720 201480 50880
rect 201320 50880 201480 51040
rect 201320 51040 201480 51200
rect 201320 51200 201480 51360
rect 201320 51360 201480 51520
rect 201320 51520 201480 51680
rect 201320 51680 201480 51840
rect 201320 51840 201480 52000
rect 201320 52000 201480 52160
rect 201320 52160 201480 52320
rect 201320 52320 201480 52480
rect 201320 52480 201480 52640
rect 201320 52640 201480 52800
rect 201320 52800 201480 52960
rect 201320 52960 201480 53120
rect 201480 50240 201640 50400
rect 201480 50400 201640 50560
rect 201480 50560 201640 50720
rect 201480 50720 201640 50880
rect 201480 50880 201640 51040
rect 201480 51040 201640 51200
rect 201480 51200 201640 51360
rect 201480 51360 201640 51520
rect 201480 51520 201640 51680
rect 201480 51680 201640 51840
rect 201480 51840 201640 52000
rect 201480 52000 201640 52160
rect 201480 52160 201640 52320
rect 201480 52320 201640 52480
rect 201480 52480 201640 52640
rect 201480 52640 201640 52800
rect 201480 52800 201640 52960
rect 201640 50400 201800 50560
rect 201640 50560 201800 50720
rect 201640 50720 201800 50880
rect 201640 50880 201800 51040
rect 201640 51040 201800 51200
rect 201640 51200 201800 51360
rect 201640 51360 201800 51520
rect 201640 51520 201800 51680
rect 201640 51680 201800 51840
rect 201640 51840 201800 52000
rect 201640 52000 201800 52160
rect 201640 52160 201800 52320
rect 201640 52320 201800 52480
rect 201640 52480 201800 52640
rect 201640 52640 201800 52800
rect 201640 52800 201800 52960
rect 201800 50560 201960 50720
rect 201800 50720 201960 50880
rect 201800 50880 201960 51040
rect 201800 51040 201960 51200
rect 201800 51200 201960 51360
rect 201800 51360 201960 51520
rect 201800 51520 201960 51680
rect 201800 51680 201960 51840
rect 201800 51840 201960 52000
rect 201800 52000 201960 52160
rect 201800 52160 201960 52320
rect 201800 52320 201960 52480
rect 201800 52480 201960 52640
rect 201800 52640 201960 52800
rect 201960 50720 202120 50880
rect 201960 50880 202120 51040
rect 201960 51040 202120 51200
rect 201960 51200 202120 51360
rect 201960 51360 202120 51520
rect 201960 51520 202120 51680
rect 201960 51680 202120 51840
rect 201960 51840 202120 52000
rect 201960 52000 202120 52160
rect 201960 52160 202120 52320
rect 201960 52320 202120 52480
rect 201960 52480 202120 52640
rect 201960 52640 202120 52800
rect 202120 50720 202280 50880
rect 202120 50880 202280 51040
rect 202120 51040 202280 51200
rect 202120 51200 202280 51360
rect 202120 51360 202280 51520
rect 202120 51520 202280 51680
rect 202120 51680 202280 51840
rect 202120 51840 202280 52000
rect 202120 52000 202280 52160
rect 202120 52160 202280 52320
rect 202120 52320 202280 52480
rect 202120 52480 202280 52640
rect 202280 50880 202440 51040
rect 202280 51040 202440 51200
rect 202280 51200 202440 51360
rect 202280 51360 202440 51520
rect 202280 51520 202440 51680
rect 202280 51680 202440 51840
rect 202280 51840 202440 52000
rect 202280 52000 202440 52160
rect 202280 52160 202440 52320
rect 202280 52320 202440 52480
rect 202280 52480 202440 52640
rect 202440 50880 202600 51040
rect 202440 51040 202600 51200
rect 202440 51200 202600 51360
rect 202440 51360 202600 51520
rect 202440 51520 202600 51680
rect 202440 51680 202600 51840
rect 202440 51840 202600 52000
rect 202440 52000 202600 52160
rect 202440 52160 202600 52320
rect 202440 52320 202600 52480
rect 202600 51040 202760 51200
rect 202600 51200 202760 51360
rect 202600 51360 202760 51520
rect 202600 51520 202760 51680
rect 202600 51680 202760 51840
rect 202600 51840 202760 52000
rect 202600 52000 202760 52160
rect 202600 52160 202760 52320
rect 202760 51040 202920 51200
rect 202760 51200 202920 51360
rect 202760 51360 202920 51520
rect 202760 51520 202920 51680
rect 202760 51680 202920 51840
rect 202760 51840 202920 52000
rect 202760 52000 202920 52160
rect 202920 51200 203080 51360
rect 202920 51360 203080 51520
rect 202920 51520 203080 51680
rect 202920 51680 203080 51840
rect 202920 51840 203080 52000
rect 203080 51360 203240 51520
rect 203080 51520 203240 51680
rect 205480 27040 205640 27200
rect 205480 27200 205640 27360
rect 205480 27360 205640 27520
rect 205480 27520 205640 27680
rect 205480 27680 205640 27840
rect 205480 27840 205640 28000
rect 205480 28000 205640 28160
rect 205480 28160 205640 28320
rect 205480 28320 205640 28480
rect 205480 28480 205640 28640
rect 205480 28640 205640 28800
rect 205480 28800 205640 28960
rect 205480 28960 205640 29120
rect 205640 26720 205800 26880
rect 205640 26880 205800 27040
rect 205640 27040 205800 27200
rect 205640 27200 205800 27360
rect 205640 27360 205800 27520
rect 205640 27520 205800 27680
rect 205640 27680 205800 27840
rect 205640 27840 205800 28000
rect 205640 28000 205800 28160
rect 205640 28160 205800 28320
rect 205640 28320 205800 28480
rect 205640 28480 205800 28640
rect 205640 28640 205800 28800
rect 205640 28800 205800 28960
rect 205640 28960 205800 29120
rect 205640 29120 205800 29280
rect 205640 29280 205800 29440
rect 205640 29440 205800 29600
rect 205640 29600 205800 29760
rect 205640 29760 205800 29920
rect 205640 29920 205800 30080
rect 205640 30080 205800 30240
rect 205640 30240 205800 30400
rect 205640 30400 205800 30560
rect 205640 30560 205800 30720
rect 205640 30720 205800 30880
rect 205640 30880 205800 31040
rect 205640 31040 205800 31200
rect 205640 31200 205800 31360
rect 205640 31520 205800 31680
rect 205640 31840 205800 32000
rect 205640 32160 205800 32320
rect 205640 32480 205800 32640
rect 205640 32800 205800 32960
rect 205640 33280 205800 33440
rect 205800 26560 205960 26720
rect 205800 26720 205960 26880
rect 205800 26880 205960 27040
rect 205800 27040 205960 27200
rect 205800 27200 205960 27360
rect 205800 27360 205960 27520
rect 205800 27520 205960 27680
rect 205800 27680 205960 27840
rect 205800 27840 205960 28000
rect 205800 28000 205960 28160
rect 205800 28160 205960 28320
rect 205800 28320 205960 28480
rect 205800 28480 205960 28640
rect 205800 28640 205960 28800
rect 205800 28800 205960 28960
rect 205800 28960 205960 29120
rect 205800 29120 205960 29280
rect 205800 29280 205960 29440
rect 205800 29440 205960 29600
rect 205800 29600 205960 29760
rect 205800 29760 205960 29920
rect 205800 29920 205960 30080
rect 205800 30080 205960 30240
rect 205800 30240 205960 30400
rect 205800 30400 205960 30560
rect 205800 30560 205960 30720
rect 205800 30720 205960 30880
rect 205800 30880 205960 31040
rect 205800 31040 205960 31200
rect 205800 31200 205960 31360
rect 205800 31360 205960 31520
rect 205800 31520 205960 31680
rect 205800 31680 205960 31840
rect 205800 31840 205960 32000
rect 205800 32000 205960 32160
rect 205800 32160 205960 32320
rect 205800 32320 205960 32480
rect 205800 32480 205960 32640
rect 205800 32640 205960 32800
rect 205800 32800 205960 32960
rect 205800 32960 205960 33120
rect 205800 33120 205960 33280
rect 205800 33280 205960 33440
rect 205800 33440 205960 33600
rect 205800 33600 205960 33760
rect 205800 33760 205960 33920
rect 205800 33920 205960 34080
rect 205800 34080 205960 34240
rect 205800 34240 205960 34400
rect 205800 34400 205960 34560
rect 205800 34560 205960 34720
rect 205800 34720 205960 34880
rect 205800 34880 205960 35040
rect 205800 35040 205960 35200
rect 205800 35200 205960 35360
rect 205800 35360 205960 35520
rect 205800 35520 205960 35680
rect 205800 35680 205960 35840
rect 205800 35840 205960 36000
rect 205800 36000 205960 36160
rect 205800 36160 205960 36320
rect 205800 36320 205960 36480
rect 205800 36480 205960 36640
rect 205800 36640 205960 36800
rect 205800 36800 205960 36960
rect 205800 36960 205960 37120
rect 205800 37120 205960 37280
rect 205800 37280 205960 37440
rect 205800 37440 205960 37600
rect 205800 37600 205960 37760
rect 205800 37920 205960 38080
rect 205800 49600 205960 49760
rect 205800 49760 205960 49920
rect 205800 49920 205960 50080
rect 205800 50080 205960 50240
rect 205800 50240 205960 50400
rect 205800 50400 205960 50560
rect 205800 50560 205960 50720
rect 205800 50720 205960 50880
rect 205800 50880 205960 51040
rect 205800 51040 205960 51200
rect 205960 26400 206120 26560
rect 205960 26560 206120 26720
rect 205960 26720 206120 26880
rect 205960 26880 206120 27040
rect 205960 27040 206120 27200
rect 205960 27200 206120 27360
rect 205960 27360 206120 27520
rect 205960 27520 206120 27680
rect 205960 27680 206120 27840
rect 205960 27840 206120 28000
rect 205960 28000 206120 28160
rect 205960 28160 206120 28320
rect 205960 28320 206120 28480
rect 205960 28480 206120 28640
rect 205960 28640 206120 28800
rect 205960 28800 206120 28960
rect 205960 28960 206120 29120
rect 205960 29120 206120 29280
rect 205960 29280 206120 29440
rect 205960 29440 206120 29600
rect 205960 29600 206120 29760
rect 205960 29760 206120 29920
rect 205960 29920 206120 30080
rect 205960 30080 206120 30240
rect 205960 30240 206120 30400
rect 205960 30400 206120 30560
rect 205960 30560 206120 30720
rect 205960 30720 206120 30880
rect 205960 30880 206120 31040
rect 205960 31040 206120 31200
rect 205960 31200 206120 31360
rect 205960 31360 206120 31520
rect 205960 31520 206120 31680
rect 205960 31680 206120 31840
rect 205960 31840 206120 32000
rect 205960 32000 206120 32160
rect 205960 32160 206120 32320
rect 205960 32320 206120 32480
rect 205960 32480 206120 32640
rect 205960 32640 206120 32800
rect 205960 32800 206120 32960
rect 205960 32960 206120 33120
rect 205960 33120 206120 33280
rect 205960 33280 206120 33440
rect 205960 33440 206120 33600
rect 205960 33600 206120 33760
rect 205960 33760 206120 33920
rect 205960 33920 206120 34080
rect 205960 34080 206120 34240
rect 205960 34240 206120 34400
rect 205960 34400 206120 34560
rect 205960 34560 206120 34720
rect 205960 34720 206120 34880
rect 205960 34880 206120 35040
rect 205960 35040 206120 35200
rect 205960 35200 206120 35360
rect 205960 35360 206120 35520
rect 205960 35520 206120 35680
rect 205960 35680 206120 35840
rect 205960 35840 206120 36000
rect 205960 36000 206120 36160
rect 205960 36160 206120 36320
rect 205960 36320 206120 36480
rect 205960 36480 206120 36640
rect 205960 36640 206120 36800
rect 205960 36800 206120 36960
rect 205960 36960 206120 37120
rect 205960 37120 206120 37280
rect 205960 37280 206120 37440
rect 205960 37440 206120 37600
rect 205960 37600 206120 37760
rect 205960 37760 206120 37920
rect 205960 37920 206120 38080
rect 205960 38080 206120 38240
rect 205960 38240 206120 38400
rect 205960 38400 206120 38560
rect 205960 38560 206120 38720
rect 205960 38720 206120 38880
rect 205960 38880 206120 39040
rect 205960 39040 206120 39200
rect 205960 39200 206120 39360
rect 205960 39360 206120 39520
rect 205960 39520 206120 39680
rect 205960 39680 206120 39840
rect 205960 39840 206120 40000
rect 205960 40000 206120 40160
rect 205960 40160 206120 40320
rect 205960 40480 206120 40640
rect 205960 49280 206120 49440
rect 205960 49440 206120 49600
rect 205960 49600 206120 49760
rect 205960 49760 206120 49920
rect 205960 49920 206120 50080
rect 205960 50080 206120 50240
rect 205960 50240 206120 50400
rect 205960 50400 206120 50560
rect 205960 50560 206120 50720
rect 205960 50720 206120 50880
rect 205960 50880 206120 51040
rect 205960 51040 206120 51200
rect 205960 51200 206120 51360
rect 205960 51360 206120 51520
rect 205960 51520 206120 51680
rect 205960 51680 206120 51840
rect 206120 26240 206280 26400
rect 206120 26400 206280 26560
rect 206120 26560 206280 26720
rect 206120 26720 206280 26880
rect 206120 26880 206280 27040
rect 206120 27040 206280 27200
rect 206120 27200 206280 27360
rect 206120 27360 206280 27520
rect 206120 27520 206280 27680
rect 206120 27680 206280 27840
rect 206120 27840 206280 28000
rect 206120 28000 206280 28160
rect 206120 28160 206280 28320
rect 206120 28320 206280 28480
rect 206120 28480 206280 28640
rect 206120 28640 206280 28800
rect 206120 28800 206280 28960
rect 206120 28960 206280 29120
rect 206120 29120 206280 29280
rect 206120 29280 206280 29440
rect 206120 29440 206280 29600
rect 206120 29600 206280 29760
rect 206120 29760 206280 29920
rect 206120 29920 206280 30080
rect 206120 30080 206280 30240
rect 206120 30240 206280 30400
rect 206120 30400 206280 30560
rect 206120 30560 206280 30720
rect 206120 30720 206280 30880
rect 206120 30880 206280 31040
rect 206120 31040 206280 31200
rect 206120 31200 206280 31360
rect 206120 31360 206280 31520
rect 206120 31520 206280 31680
rect 206120 31680 206280 31840
rect 206120 31840 206280 32000
rect 206120 32000 206280 32160
rect 206120 32160 206280 32320
rect 206120 32320 206280 32480
rect 206120 32480 206280 32640
rect 206120 32640 206280 32800
rect 206120 32800 206280 32960
rect 206120 32960 206280 33120
rect 206120 33120 206280 33280
rect 206120 33280 206280 33440
rect 206120 33440 206280 33600
rect 206120 33600 206280 33760
rect 206120 33760 206280 33920
rect 206120 33920 206280 34080
rect 206120 34080 206280 34240
rect 206120 34240 206280 34400
rect 206120 34400 206280 34560
rect 206120 34560 206280 34720
rect 206120 34720 206280 34880
rect 206120 34880 206280 35040
rect 206120 35040 206280 35200
rect 206120 35200 206280 35360
rect 206120 35360 206280 35520
rect 206120 35520 206280 35680
rect 206120 35680 206280 35840
rect 206120 35840 206280 36000
rect 206120 36000 206280 36160
rect 206120 36160 206280 36320
rect 206120 36320 206280 36480
rect 206120 36480 206280 36640
rect 206120 36640 206280 36800
rect 206120 36800 206280 36960
rect 206120 36960 206280 37120
rect 206120 37120 206280 37280
rect 206120 37280 206280 37440
rect 206120 37440 206280 37600
rect 206120 37600 206280 37760
rect 206120 37760 206280 37920
rect 206120 37920 206280 38080
rect 206120 38080 206280 38240
rect 206120 38240 206280 38400
rect 206120 38400 206280 38560
rect 206120 38560 206280 38720
rect 206120 38720 206280 38880
rect 206120 38880 206280 39040
rect 206120 39040 206280 39200
rect 206120 39200 206280 39360
rect 206120 39360 206280 39520
rect 206120 39520 206280 39680
rect 206120 39680 206280 39840
rect 206120 39840 206280 40000
rect 206120 40000 206280 40160
rect 206120 40160 206280 40320
rect 206120 40320 206280 40480
rect 206120 40480 206280 40640
rect 206120 40640 206280 40800
rect 206120 40800 206280 40960
rect 206120 40960 206280 41120
rect 206120 41120 206280 41280
rect 206120 41280 206280 41440
rect 206120 41440 206280 41600
rect 206120 41600 206280 41760
rect 206120 41760 206280 41920
rect 206120 41920 206280 42080
rect 206120 42080 206280 42240
rect 206120 42240 206280 42400
rect 206120 48960 206280 49120
rect 206120 49120 206280 49280
rect 206120 49280 206280 49440
rect 206120 49440 206280 49600
rect 206120 49600 206280 49760
rect 206120 49760 206280 49920
rect 206120 49920 206280 50080
rect 206120 50080 206280 50240
rect 206120 50240 206280 50400
rect 206120 50400 206280 50560
rect 206120 50560 206280 50720
rect 206120 50720 206280 50880
rect 206120 50880 206280 51040
rect 206120 51040 206280 51200
rect 206120 51200 206280 51360
rect 206120 51360 206280 51520
rect 206120 51520 206280 51680
rect 206120 51680 206280 51840
rect 206120 51840 206280 52000
rect 206120 52000 206280 52160
rect 206280 26240 206440 26400
rect 206280 26400 206440 26560
rect 206280 26560 206440 26720
rect 206280 26720 206440 26880
rect 206280 26880 206440 27040
rect 206280 27040 206440 27200
rect 206280 27200 206440 27360
rect 206280 27360 206440 27520
rect 206280 27520 206440 27680
rect 206280 27680 206440 27840
rect 206280 27840 206440 28000
rect 206280 28000 206440 28160
rect 206280 28160 206440 28320
rect 206280 28320 206440 28480
rect 206280 28480 206440 28640
rect 206280 28640 206440 28800
rect 206280 28800 206440 28960
rect 206280 28960 206440 29120
rect 206280 29120 206440 29280
rect 206280 29280 206440 29440
rect 206280 29440 206440 29600
rect 206280 29600 206440 29760
rect 206280 29760 206440 29920
rect 206280 29920 206440 30080
rect 206280 30080 206440 30240
rect 206280 30240 206440 30400
rect 206280 30400 206440 30560
rect 206280 30560 206440 30720
rect 206280 30720 206440 30880
rect 206280 30880 206440 31040
rect 206280 31040 206440 31200
rect 206280 31200 206440 31360
rect 206280 31360 206440 31520
rect 206280 31520 206440 31680
rect 206280 31680 206440 31840
rect 206280 31840 206440 32000
rect 206280 32000 206440 32160
rect 206280 32160 206440 32320
rect 206280 32320 206440 32480
rect 206280 32480 206440 32640
rect 206280 32640 206440 32800
rect 206280 32800 206440 32960
rect 206280 32960 206440 33120
rect 206280 33120 206440 33280
rect 206280 33280 206440 33440
rect 206280 33440 206440 33600
rect 206280 33600 206440 33760
rect 206280 33760 206440 33920
rect 206280 33920 206440 34080
rect 206280 34080 206440 34240
rect 206280 34240 206440 34400
rect 206280 34400 206440 34560
rect 206280 34560 206440 34720
rect 206280 34720 206440 34880
rect 206280 34880 206440 35040
rect 206280 35040 206440 35200
rect 206280 35200 206440 35360
rect 206280 35360 206440 35520
rect 206280 35520 206440 35680
rect 206280 35680 206440 35840
rect 206280 35840 206440 36000
rect 206280 36000 206440 36160
rect 206280 36160 206440 36320
rect 206280 36320 206440 36480
rect 206280 36480 206440 36640
rect 206280 36640 206440 36800
rect 206280 36800 206440 36960
rect 206280 36960 206440 37120
rect 206280 37120 206440 37280
rect 206280 37280 206440 37440
rect 206280 37440 206440 37600
rect 206280 37600 206440 37760
rect 206280 37760 206440 37920
rect 206280 37920 206440 38080
rect 206280 38080 206440 38240
rect 206280 38240 206440 38400
rect 206280 38400 206440 38560
rect 206280 38560 206440 38720
rect 206280 38720 206440 38880
rect 206280 38880 206440 39040
rect 206280 39040 206440 39200
rect 206280 39200 206440 39360
rect 206280 39360 206440 39520
rect 206280 39520 206440 39680
rect 206280 39680 206440 39840
rect 206280 39840 206440 40000
rect 206280 40000 206440 40160
rect 206280 40160 206440 40320
rect 206280 40320 206440 40480
rect 206280 40480 206440 40640
rect 206280 40640 206440 40800
rect 206280 40800 206440 40960
rect 206280 40960 206440 41120
rect 206280 41120 206440 41280
rect 206280 41280 206440 41440
rect 206280 41440 206440 41600
rect 206280 41600 206440 41760
rect 206280 41760 206440 41920
rect 206280 41920 206440 42080
rect 206280 42080 206440 42240
rect 206280 42240 206440 42400
rect 206280 42400 206440 42560
rect 206280 42560 206440 42720
rect 206280 42720 206440 42880
rect 206280 48640 206440 48800
rect 206280 48800 206440 48960
rect 206280 48960 206440 49120
rect 206280 49120 206440 49280
rect 206280 49280 206440 49440
rect 206280 49440 206440 49600
rect 206280 49600 206440 49760
rect 206280 49760 206440 49920
rect 206280 49920 206440 50080
rect 206280 50080 206440 50240
rect 206280 50240 206440 50400
rect 206280 50400 206440 50560
rect 206280 50560 206440 50720
rect 206280 50720 206440 50880
rect 206280 50880 206440 51040
rect 206280 51040 206440 51200
rect 206280 51200 206440 51360
rect 206280 51360 206440 51520
rect 206280 51520 206440 51680
rect 206280 51680 206440 51840
rect 206280 51840 206440 52000
rect 206280 52000 206440 52160
rect 206280 52160 206440 52320
rect 206280 52320 206440 52480
rect 206440 26080 206600 26240
rect 206440 26240 206600 26400
rect 206440 26400 206600 26560
rect 206440 26560 206600 26720
rect 206440 26720 206600 26880
rect 206440 26880 206600 27040
rect 206440 27040 206600 27200
rect 206440 27200 206600 27360
rect 206440 27360 206600 27520
rect 206440 27520 206600 27680
rect 206440 27680 206600 27840
rect 206440 27840 206600 28000
rect 206440 28000 206600 28160
rect 206440 28160 206600 28320
rect 206440 28320 206600 28480
rect 206440 28480 206600 28640
rect 206440 28640 206600 28800
rect 206440 28800 206600 28960
rect 206440 28960 206600 29120
rect 206440 29120 206600 29280
rect 206440 29280 206600 29440
rect 206440 29440 206600 29600
rect 206440 29600 206600 29760
rect 206440 29760 206600 29920
rect 206440 29920 206600 30080
rect 206440 30080 206600 30240
rect 206440 30240 206600 30400
rect 206440 30400 206600 30560
rect 206440 30560 206600 30720
rect 206440 30720 206600 30880
rect 206440 30880 206600 31040
rect 206440 31040 206600 31200
rect 206440 31200 206600 31360
rect 206440 31360 206600 31520
rect 206440 31520 206600 31680
rect 206440 31680 206600 31840
rect 206440 31840 206600 32000
rect 206440 32000 206600 32160
rect 206440 32160 206600 32320
rect 206440 32320 206600 32480
rect 206440 32480 206600 32640
rect 206440 32640 206600 32800
rect 206440 32800 206600 32960
rect 206440 32960 206600 33120
rect 206440 33120 206600 33280
rect 206440 33280 206600 33440
rect 206440 33440 206600 33600
rect 206440 33600 206600 33760
rect 206440 33760 206600 33920
rect 206440 33920 206600 34080
rect 206440 34080 206600 34240
rect 206440 34240 206600 34400
rect 206440 34400 206600 34560
rect 206440 34560 206600 34720
rect 206440 34720 206600 34880
rect 206440 34880 206600 35040
rect 206440 35040 206600 35200
rect 206440 35200 206600 35360
rect 206440 35360 206600 35520
rect 206440 35520 206600 35680
rect 206440 35680 206600 35840
rect 206440 35840 206600 36000
rect 206440 36000 206600 36160
rect 206440 36160 206600 36320
rect 206440 36320 206600 36480
rect 206440 36480 206600 36640
rect 206440 36640 206600 36800
rect 206440 36800 206600 36960
rect 206440 36960 206600 37120
rect 206440 37120 206600 37280
rect 206440 37280 206600 37440
rect 206440 37440 206600 37600
rect 206440 37600 206600 37760
rect 206440 37760 206600 37920
rect 206440 37920 206600 38080
rect 206440 38080 206600 38240
rect 206440 38240 206600 38400
rect 206440 38400 206600 38560
rect 206440 38560 206600 38720
rect 206440 38720 206600 38880
rect 206440 38880 206600 39040
rect 206440 39040 206600 39200
rect 206440 39200 206600 39360
rect 206440 39360 206600 39520
rect 206440 39520 206600 39680
rect 206440 39680 206600 39840
rect 206440 39840 206600 40000
rect 206440 40000 206600 40160
rect 206440 40160 206600 40320
rect 206440 40320 206600 40480
rect 206440 40480 206600 40640
rect 206440 40640 206600 40800
rect 206440 40800 206600 40960
rect 206440 40960 206600 41120
rect 206440 41120 206600 41280
rect 206440 41280 206600 41440
rect 206440 41440 206600 41600
rect 206440 41600 206600 41760
rect 206440 41760 206600 41920
rect 206440 41920 206600 42080
rect 206440 42080 206600 42240
rect 206440 42240 206600 42400
rect 206440 42400 206600 42560
rect 206440 42560 206600 42720
rect 206440 42720 206600 42880
rect 206440 42880 206600 43040
rect 206440 43040 206600 43200
rect 206440 48480 206600 48640
rect 206440 48640 206600 48800
rect 206440 48800 206600 48960
rect 206440 48960 206600 49120
rect 206440 49120 206600 49280
rect 206440 49280 206600 49440
rect 206440 49440 206600 49600
rect 206440 49600 206600 49760
rect 206440 49760 206600 49920
rect 206440 49920 206600 50080
rect 206440 50080 206600 50240
rect 206440 50240 206600 50400
rect 206440 50400 206600 50560
rect 206440 50560 206600 50720
rect 206440 50720 206600 50880
rect 206440 50880 206600 51040
rect 206440 51040 206600 51200
rect 206440 51200 206600 51360
rect 206440 51360 206600 51520
rect 206440 51520 206600 51680
rect 206440 51680 206600 51840
rect 206440 51840 206600 52000
rect 206440 52000 206600 52160
rect 206440 52160 206600 52320
rect 206440 52320 206600 52480
rect 206440 52480 206600 52640
rect 206440 52640 206600 52800
rect 206600 26080 206760 26240
rect 206600 26240 206760 26400
rect 206600 26400 206760 26560
rect 206600 26560 206760 26720
rect 206600 26720 206760 26880
rect 206600 26880 206760 27040
rect 206600 27040 206760 27200
rect 206600 27200 206760 27360
rect 206600 27360 206760 27520
rect 206600 27520 206760 27680
rect 206600 27680 206760 27840
rect 206600 27840 206760 28000
rect 206600 28000 206760 28160
rect 206600 28160 206760 28320
rect 206600 28320 206760 28480
rect 206600 28480 206760 28640
rect 206600 28640 206760 28800
rect 206600 28800 206760 28960
rect 206600 28960 206760 29120
rect 206600 29120 206760 29280
rect 206600 29280 206760 29440
rect 206600 29440 206760 29600
rect 206600 29600 206760 29760
rect 206600 29760 206760 29920
rect 206600 29920 206760 30080
rect 206600 30080 206760 30240
rect 206600 30240 206760 30400
rect 206600 30400 206760 30560
rect 206600 30560 206760 30720
rect 206600 30720 206760 30880
rect 206600 30880 206760 31040
rect 206600 31040 206760 31200
rect 206600 31200 206760 31360
rect 206600 31360 206760 31520
rect 206600 31520 206760 31680
rect 206600 31680 206760 31840
rect 206600 31840 206760 32000
rect 206600 32000 206760 32160
rect 206600 32160 206760 32320
rect 206600 32320 206760 32480
rect 206600 32480 206760 32640
rect 206600 32640 206760 32800
rect 206600 32800 206760 32960
rect 206600 32960 206760 33120
rect 206600 33120 206760 33280
rect 206600 33280 206760 33440
rect 206600 33440 206760 33600
rect 206600 33600 206760 33760
rect 206600 33760 206760 33920
rect 206600 33920 206760 34080
rect 206600 34080 206760 34240
rect 206600 34240 206760 34400
rect 206600 34400 206760 34560
rect 206600 34560 206760 34720
rect 206600 34720 206760 34880
rect 206600 34880 206760 35040
rect 206600 35040 206760 35200
rect 206600 35200 206760 35360
rect 206600 35360 206760 35520
rect 206600 35520 206760 35680
rect 206600 35680 206760 35840
rect 206600 35840 206760 36000
rect 206600 36000 206760 36160
rect 206600 36160 206760 36320
rect 206600 36320 206760 36480
rect 206600 36480 206760 36640
rect 206600 36640 206760 36800
rect 206600 36800 206760 36960
rect 206600 36960 206760 37120
rect 206600 37120 206760 37280
rect 206600 37280 206760 37440
rect 206600 37440 206760 37600
rect 206600 37600 206760 37760
rect 206600 37760 206760 37920
rect 206600 37920 206760 38080
rect 206600 38080 206760 38240
rect 206600 38240 206760 38400
rect 206600 38400 206760 38560
rect 206600 38560 206760 38720
rect 206600 38720 206760 38880
rect 206600 38880 206760 39040
rect 206600 39040 206760 39200
rect 206600 39200 206760 39360
rect 206600 39360 206760 39520
rect 206600 39520 206760 39680
rect 206600 39680 206760 39840
rect 206600 39840 206760 40000
rect 206600 40000 206760 40160
rect 206600 40160 206760 40320
rect 206600 40320 206760 40480
rect 206600 40480 206760 40640
rect 206600 40640 206760 40800
rect 206600 40800 206760 40960
rect 206600 40960 206760 41120
rect 206600 41120 206760 41280
rect 206600 41280 206760 41440
rect 206600 41440 206760 41600
rect 206600 41600 206760 41760
rect 206600 41760 206760 41920
rect 206600 41920 206760 42080
rect 206600 42080 206760 42240
rect 206600 42240 206760 42400
rect 206600 42400 206760 42560
rect 206600 42560 206760 42720
rect 206600 42720 206760 42880
rect 206600 42880 206760 43040
rect 206600 43040 206760 43200
rect 206600 43200 206760 43360
rect 206600 43360 206760 43520
rect 206600 48320 206760 48480
rect 206600 48480 206760 48640
rect 206600 48640 206760 48800
rect 206600 48800 206760 48960
rect 206600 48960 206760 49120
rect 206600 49120 206760 49280
rect 206600 49280 206760 49440
rect 206600 49440 206760 49600
rect 206600 49600 206760 49760
rect 206600 49760 206760 49920
rect 206600 49920 206760 50080
rect 206600 50080 206760 50240
rect 206600 50240 206760 50400
rect 206600 50400 206760 50560
rect 206600 50560 206760 50720
rect 206600 50720 206760 50880
rect 206600 50880 206760 51040
rect 206600 51040 206760 51200
rect 206600 51200 206760 51360
rect 206600 51360 206760 51520
rect 206600 51520 206760 51680
rect 206600 51680 206760 51840
rect 206600 51840 206760 52000
rect 206600 52000 206760 52160
rect 206600 52160 206760 52320
rect 206600 52320 206760 52480
rect 206600 52480 206760 52640
rect 206600 52640 206760 52800
rect 206600 52800 206760 52960
rect 206600 52960 206760 53120
rect 206760 25920 206920 26080
rect 206760 26080 206920 26240
rect 206760 26240 206920 26400
rect 206760 26400 206920 26560
rect 206760 26560 206920 26720
rect 206760 26720 206920 26880
rect 206760 26880 206920 27040
rect 206760 27040 206920 27200
rect 206760 27200 206920 27360
rect 206760 27360 206920 27520
rect 206760 27520 206920 27680
rect 206760 27680 206920 27840
rect 206760 27840 206920 28000
rect 206760 28000 206920 28160
rect 206760 28160 206920 28320
rect 206760 28320 206920 28480
rect 206760 28480 206920 28640
rect 206760 28640 206920 28800
rect 206760 28800 206920 28960
rect 206760 28960 206920 29120
rect 206760 29120 206920 29280
rect 206760 29280 206920 29440
rect 206760 29440 206920 29600
rect 206760 29600 206920 29760
rect 206760 29760 206920 29920
rect 206760 29920 206920 30080
rect 206760 30080 206920 30240
rect 206760 30240 206920 30400
rect 206760 30400 206920 30560
rect 206760 30560 206920 30720
rect 206760 30720 206920 30880
rect 206760 30880 206920 31040
rect 206760 31040 206920 31200
rect 206760 31200 206920 31360
rect 206760 31360 206920 31520
rect 206760 31520 206920 31680
rect 206760 31680 206920 31840
rect 206760 31840 206920 32000
rect 206760 32000 206920 32160
rect 206760 32160 206920 32320
rect 206760 32320 206920 32480
rect 206760 32480 206920 32640
rect 206760 32640 206920 32800
rect 206760 32800 206920 32960
rect 206760 32960 206920 33120
rect 206760 33120 206920 33280
rect 206760 33280 206920 33440
rect 206760 33440 206920 33600
rect 206760 33600 206920 33760
rect 206760 33760 206920 33920
rect 206760 33920 206920 34080
rect 206760 34080 206920 34240
rect 206760 34240 206920 34400
rect 206760 34400 206920 34560
rect 206760 34560 206920 34720
rect 206760 34720 206920 34880
rect 206760 34880 206920 35040
rect 206760 35040 206920 35200
rect 206760 35200 206920 35360
rect 206760 35360 206920 35520
rect 206760 35520 206920 35680
rect 206760 35680 206920 35840
rect 206760 35840 206920 36000
rect 206760 36000 206920 36160
rect 206760 36160 206920 36320
rect 206760 36320 206920 36480
rect 206760 36480 206920 36640
rect 206760 36640 206920 36800
rect 206760 36800 206920 36960
rect 206760 36960 206920 37120
rect 206760 37120 206920 37280
rect 206760 37280 206920 37440
rect 206760 37440 206920 37600
rect 206760 37600 206920 37760
rect 206760 37760 206920 37920
rect 206760 37920 206920 38080
rect 206760 38080 206920 38240
rect 206760 38240 206920 38400
rect 206760 38400 206920 38560
rect 206760 38560 206920 38720
rect 206760 38720 206920 38880
rect 206760 38880 206920 39040
rect 206760 39040 206920 39200
rect 206760 39200 206920 39360
rect 206760 39360 206920 39520
rect 206760 39520 206920 39680
rect 206760 39680 206920 39840
rect 206760 39840 206920 40000
rect 206760 40000 206920 40160
rect 206760 40160 206920 40320
rect 206760 40320 206920 40480
rect 206760 40480 206920 40640
rect 206760 40640 206920 40800
rect 206760 40800 206920 40960
rect 206760 40960 206920 41120
rect 206760 41120 206920 41280
rect 206760 41280 206920 41440
rect 206760 41440 206920 41600
rect 206760 41600 206920 41760
rect 206760 41760 206920 41920
rect 206760 41920 206920 42080
rect 206760 42080 206920 42240
rect 206760 42240 206920 42400
rect 206760 42400 206920 42560
rect 206760 42560 206920 42720
rect 206760 42720 206920 42880
rect 206760 42880 206920 43040
rect 206760 43040 206920 43200
rect 206760 43200 206920 43360
rect 206760 43360 206920 43520
rect 206760 43520 206920 43680
rect 206760 43680 206920 43840
rect 206760 48160 206920 48320
rect 206760 48320 206920 48480
rect 206760 48480 206920 48640
rect 206760 48640 206920 48800
rect 206760 48800 206920 48960
rect 206760 48960 206920 49120
rect 206760 49120 206920 49280
rect 206760 49280 206920 49440
rect 206760 49440 206920 49600
rect 206760 49600 206920 49760
rect 206760 49760 206920 49920
rect 206760 49920 206920 50080
rect 206760 50080 206920 50240
rect 206760 50240 206920 50400
rect 206760 50400 206920 50560
rect 206760 50560 206920 50720
rect 206760 50720 206920 50880
rect 206760 50880 206920 51040
rect 206760 51040 206920 51200
rect 206760 51200 206920 51360
rect 206760 51360 206920 51520
rect 206760 51520 206920 51680
rect 206760 51680 206920 51840
rect 206760 51840 206920 52000
rect 206760 52000 206920 52160
rect 206760 52160 206920 52320
rect 206760 52320 206920 52480
rect 206760 52480 206920 52640
rect 206760 52640 206920 52800
rect 206760 52800 206920 52960
rect 206760 52960 206920 53120
rect 206760 53120 206920 53280
rect 206920 25920 207080 26080
rect 206920 26080 207080 26240
rect 206920 26240 207080 26400
rect 206920 26400 207080 26560
rect 206920 26560 207080 26720
rect 206920 26720 207080 26880
rect 206920 26880 207080 27040
rect 206920 27040 207080 27200
rect 206920 27200 207080 27360
rect 206920 27360 207080 27520
rect 206920 27520 207080 27680
rect 206920 27680 207080 27840
rect 206920 27840 207080 28000
rect 206920 28000 207080 28160
rect 206920 28160 207080 28320
rect 206920 28320 207080 28480
rect 206920 28480 207080 28640
rect 206920 28640 207080 28800
rect 206920 28800 207080 28960
rect 206920 28960 207080 29120
rect 206920 29120 207080 29280
rect 206920 29280 207080 29440
rect 206920 29440 207080 29600
rect 206920 29600 207080 29760
rect 206920 29760 207080 29920
rect 206920 29920 207080 30080
rect 206920 30080 207080 30240
rect 206920 30240 207080 30400
rect 206920 30400 207080 30560
rect 206920 30560 207080 30720
rect 206920 30720 207080 30880
rect 206920 30880 207080 31040
rect 206920 31040 207080 31200
rect 206920 31200 207080 31360
rect 206920 31360 207080 31520
rect 206920 31520 207080 31680
rect 206920 31680 207080 31840
rect 206920 31840 207080 32000
rect 206920 32000 207080 32160
rect 206920 32160 207080 32320
rect 206920 32320 207080 32480
rect 206920 32480 207080 32640
rect 206920 32640 207080 32800
rect 206920 32800 207080 32960
rect 206920 32960 207080 33120
rect 206920 33120 207080 33280
rect 206920 33280 207080 33440
rect 206920 33440 207080 33600
rect 206920 33600 207080 33760
rect 206920 33760 207080 33920
rect 206920 33920 207080 34080
rect 206920 34080 207080 34240
rect 206920 34240 207080 34400
rect 206920 34400 207080 34560
rect 206920 34560 207080 34720
rect 206920 34720 207080 34880
rect 206920 34880 207080 35040
rect 206920 35040 207080 35200
rect 206920 35200 207080 35360
rect 206920 35360 207080 35520
rect 206920 35520 207080 35680
rect 206920 35680 207080 35840
rect 206920 35840 207080 36000
rect 206920 36000 207080 36160
rect 206920 36160 207080 36320
rect 206920 36320 207080 36480
rect 206920 36480 207080 36640
rect 206920 36640 207080 36800
rect 206920 36800 207080 36960
rect 206920 36960 207080 37120
rect 206920 37120 207080 37280
rect 206920 37280 207080 37440
rect 206920 37440 207080 37600
rect 206920 37600 207080 37760
rect 206920 37760 207080 37920
rect 206920 37920 207080 38080
rect 206920 38080 207080 38240
rect 206920 38240 207080 38400
rect 206920 38400 207080 38560
rect 206920 38560 207080 38720
rect 206920 38720 207080 38880
rect 206920 38880 207080 39040
rect 206920 39040 207080 39200
rect 206920 39200 207080 39360
rect 206920 39360 207080 39520
rect 206920 39520 207080 39680
rect 206920 39680 207080 39840
rect 206920 39840 207080 40000
rect 206920 40000 207080 40160
rect 206920 40160 207080 40320
rect 206920 40320 207080 40480
rect 206920 40480 207080 40640
rect 206920 40640 207080 40800
rect 206920 40800 207080 40960
rect 206920 40960 207080 41120
rect 206920 41120 207080 41280
rect 206920 41280 207080 41440
rect 206920 41440 207080 41600
rect 206920 41600 207080 41760
rect 206920 41760 207080 41920
rect 206920 41920 207080 42080
rect 206920 42080 207080 42240
rect 206920 42240 207080 42400
rect 206920 42400 207080 42560
rect 206920 42560 207080 42720
rect 206920 42720 207080 42880
rect 206920 42880 207080 43040
rect 206920 43040 207080 43200
rect 206920 43200 207080 43360
rect 206920 43360 207080 43520
rect 206920 43520 207080 43680
rect 206920 43680 207080 43840
rect 206920 43840 207080 44000
rect 206920 48000 207080 48160
rect 206920 48160 207080 48320
rect 206920 48320 207080 48480
rect 206920 48480 207080 48640
rect 206920 48640 207080 48800
rect 206920 48800 207080 48960
rect 206920 48960 207080 49120
rect 206920 49120 207080 49280
rect 206920 49280 207080 49440
rect 206920 49440 207080 49600
rect 206920 49600 207080 49760
rect 206920 49760 207080 49920
rect 206920 49920 207080 50080
rect 206920 50080 207080 50240
rect 206920 50240 207080 50400
rect 206920 50400 207080 50560
rect 206920 50560 207080 50720
rect 206920 50720 207080 50880
rect 206920 50880 207080 51040
rect 206920 51040 207080 51200
rect 206920 51200 207080 51360
rect 206920 51360 207080 51520
rect 206920 51520 207080 51680
rect 206920 51680 207080 51840
rect 206920 51840 207080 52000
rect 206920 52000 207080 52160
rect 206920 52160 207080 52320
rect 206920 52320 207080 52480
rect 206920 52480 207080 52640
rect 206920 52640 207080 52800
rect 206920 52800 207080 52960
rect 206920 52960 207080 53120
rect 206920 53120 207080 53280
rect 206920 53280 207080 53440
rect 207080 25920 207240 26080
rect 207080 26080 207240 26240
rect 207080 26240 207240 26400
rect 207080 26400 207240 26560
rect 207080 26560 207240 26720
rect 207080 26720 207240 26880
rect 207080 26880 207240 27040
rect 207080 27040 207240 27200
rect 207080 27200 207240 27360
rect 207080 27360 207240 27520
rect 207080 27520 207240 27680
rect 207080 27680 207240 27840
rect 207080 27840 207240 28000
rect 207080 28000 207240 28160
rect 207080 28160 207240 28320
rect 207080 28320 207240 28480
rect 207080 28480 207240 28640
rect 207080 28640 207240 28800
rect 207080 28800 207240 28960
rect 207080 28960 207240 29120
rect 207080 29120 207240 29280
rect 207080 29280 207240 29440
rect 207080 29440 207240 29600
rect 207080 29600 207240 29760
rect 207080 29760 207240 29920
rect 207080 29920 207240 30080
rect 207080 30080 207240 30240
rect 207080 30240 207240 30400
rect 207080 30400 207240 30560
rect 207080 30560 207240 30720
rect 207080 30720 207240 30880
rect 207080 30880 207240 31040
rect 207080 31040 207240 31200
rect 207080 31200 207240 31360
rect 207080 31360 207240 31520
rect 207080 31520 207240 31680
rect 207080 31680 207240 31840
rect 207080 31840 207240 32000
rect 207080 32000 207240 32160
rect 207080 32160 207240 32320
rect 207080 32320 207240 32480
rect 207080 32480 207240 32640
rect 207080 32640 207240 32800
rect 207080 32800 207240 32960
rect 207080 32960 207240 33120
rect 207080 33120 207240 33280
rect 207080 33280 207240 33440
rect 207080 33440 207240 33600
rect 207080 33600 207240 33760
rect 207080 33760 207240 33920
rect 207080 33920 207240 34080
rect 207080 34080 207240 34240
rect 207080 34240 207240 34400
rect 207080 34400 207240 34560
rect 207080 34560 207240 34720
rect 207080 34720 207240 34880
rect 207080 34880 207240 35040
rect 207080 35040 207240 35200
rect 207080 35200 207240 35360
rect 207080 35360 207240 35520
rect 207080 35520 207240 35680
rect 207080 35680 207240 35840
rect 207080 35840 207240 36000
rect 207080 36000 207240 36160
rect 207080 36160 207240 36320
rect 207080 36320 207240 36480
rect 207080 36480 207240 36640
rect 207080 36640 207240 36800
rect 207080 36800 207240 36960
rect 207080 36960 207240 37120
rect 207080 37120 207240 37280
rect 207080 37280 207240 37440
rect 207080 37440 207240 37600
rect 207080 37600 207240 37760
rect 207080 37760 207240 37920
rect 207080 37920 207240 38080
rect 207080 38080 207240 38240
rect 207080 38240 207240 38400
rect 207080 38400 207240 38560
rect 207080 38560 207240 38720
rect 207080 38720 207240 38880
rect 207080 38880 207240 39040
rect 207080 39040 207240 39200
rect 207080 39200 207240 39360
rect 207080 39360 207240 39520
rect 207080 39520 207240 39680
rect 207080 39680 207240 39840
rect 207080 39840 207240 40000
rect 207080 40000 207240 40160
rect 207080 40160 207240 40320
rect 207080 40320 207240 40480
rect 207080 40480 207240 40640
rect 207080 40640 207240 40800
rect 207080 40800 207240 40960
rect 207080 40960 207240 41120
rect 207080 41120 207240 41280
rect 207080 41280 207240 41440
rect 207080 41440 207240 41600
rect 207080 41600 207240 41760
rect 207080 41760 207240 41920
rect 207080 41920 207240 42080
rect 207080 42080 207240 42240
rect 207080 42240 207240 42400
rect 207080 42400 207240 42560
rect 207080 42560 207240 42720
rect 207080 42720 207240 42880
rect 207080 42880 207240 43040
rect 207080 43040 207240 43200
rect 207080 43200 207240 43360
rect 207080 43360 207240 43520
rect 207080 43520 207240 43680
rect 207080 43680 207240 43840
rect 207080 43840 207240 44000
rect 207080 44000 207240 44160
rect 207080 44160 207240 44320
rect 207080 47840 207240 48000
rect 207080 48000 207240 48160
rect 207080 48160 207240 48320
rect 207080 48320 207240 48480
rect 207080 48480 207240 48640
rect 207080 48640 207240 48800
rect 207080 48800 207240 48960
rect 207080 48960 207240 49120
rect 207080 49120 207240 49280
rect 207080 49280 207240 49440
rect 207080 49440 207240 49600
rect 207080 49600 207240 49760
rect 207080 49760 207240 49920
rect 207080 49920 207240 50080
rect 207080 50080 207240 50240
rect 207080 50240 207240 50400
rect 207080 50400 207240 50560
rect 207080 50560 207240 50720
rect 207080 50720 207240 50880
rect 207080 50880 207240 51040
rect 207080 51040 207240 51200
rect 207080 51200 207240 51360
rect 207080 51360 207240 51520
rect 207080 51520 207240 51680
rect 207080 51680 207240 51840
rect 207080 51840 207240 52000
rect 207080 52000 207240 52160
rect 207080 52160 207240 52320
rect 207080 52320 207240 52480
rect 207080 52480 207240 52640
rect 207080 52640 207240 52800
rect 207080 52800 207240 52960
rect 207080 52960 207240 53120
rect 207080 53120 207240 53280
rect 207080 53280 207240 53440
rect 207080 53440 207240 53600
rect 207240 25920 207400 26080
rect 207240 26080 207400 26240
rect 207240 26240 207400 26400
rect 207240 26400 207400 26560
rect 207240 26560 207400 26720
rect 207240 26720 207400 26880
rect 207240 26880 207400 27040
rect 207240 27040 207400 27200
rect 207240 27200 207400 27360
rect 207240 27360 207400 27520
rect 207240 27520 207400 27680
rect 207240 27680 207400 27840
rect 207240 27840 207400 28000
rect 207240 28000 207400 28160
rect 207240 28160 207400 28320
rect 207240 28320 207400 28480
rect 207240 28480 207400 28640
rect 207240 28640 207400 28800
rect 207240 28800 207400 28960
rect 207240 28960 207400 29120
rect 207240 29120 207400 29280
rect 207240 29280 207400 29440
rect 207240 29440 207400 29600
rect 207240 29600 207400 29760
rect 207240 29760 207400 29920
rect 207240 29920 207400 30080
rect 207240 30080 207400 30240
rect 207240 30240 207400 30400
rect 207240 30400 207400 30560
rect 207240 30560 207400 30720
rect 207240 30720 207400 30880
rect 207240 30880 207400 31040
rect 207240 31040 207400 31200
rect 207240 31200 207400 31360
rect 207240 31360 207400 31520
rect 207240 31520 207400 31680
rect 207240 31680 207400 31840
rect 207240 31840 207400 32000
rect 207240 32000 207400 32160
rect 207240 32160 207400 32320
rect 207240 32320 207400 32480
rect 207240 32480 207400 32640
rect 207240 32640 207400 32800
rect 207240 32800 207400 32960
rect 207240 32960 207400 33120
rect 207240 33120 207400 33280
rect 207240 33280 207400 33440
rect 207240 33440 207400 33600
rect 207240 33600 207400 33760
rect 207240 33760 207400 33920
rect 207240 33920 207400 34080
rect 207240 34080 207400 34240
rect 207240 34240 207400 34400
rect 207240 34400 207400 34560
rect 207240 34560 207400 34720
rect 207240 34720 207400 34880
rect 207240 34880 207400 35040
rect 207240 35040 207400 35200
rect 207240 35200 207400 35360
rect 207240 35360 207400 35520
rect 207240 35520 207400 35680
rect 207240 35680 207400 35840
rect 207240 35840 207400 36000
rect 207240 36000 207400 36160
rect 207240 36160 207400 36320
rect 207240 36320 207400 36480
rect 207240 36480 207400 36640
rect 207240 36640 207400 36800
rect 207240 36800 207400 36960
rect 207240 36960 207400 37120
rect 207240 37120 207400 37280
rect 207240 37280 207400 37440
rect 207240 37440 207400 37600
rect 207240 37600 207400 37760
rect 207240 37760 207400 37920
rect 207240 37920 207400 38080
rect 207240 38080 207400 38240
rect 207240 38240 207400 38400
rect 207240 38400 207400 38560
rect 207240 38560 207400 38720
rect 207240 38720 207400 38880
rect 207240 38880 207400 39040
rect 207240 39040 207400 39200
rect 207240 39200 207400 39360
rect 207240 39360 207400 39520
rect 207240 39520 207400 39680
rect 207240 39680 207400 39840
rect 207240 39840 207400 40000
rect 207240 40000 207400 40160
rect 207240 40160 207400 40320
rect 207240 40320 207400 40480
rect 207240 40480 207400 40640
rect 207240 40640 207400 40800
rect 207240 40800 207400 40960
rect 207240 40960 207400 41120
rect 207240 41120 207400 41280
rect 207240 41280 207400 41440
rect 207240 41440 207400 41600
rect 207240 41600 207400 41760
rect 207240 41760 207400 41920
rect 207240 41920 207400 42080
rect 207240 42080 207400 42240
rect 207240 42240 207400 42400
rect 207240 42400 207400 42560
rect 207240 42560 207400 42720
rect 207240 42720 207400 42880
rect 207240 42880 207400 43040
rect 207240 43040 207400 43200
rect 207240 43200 207400 43360
rect 207240 43360 207400 43520
rect 207240 43520 207400 43680
rect 207240 43680 207400 43840
rect 207240 43840 207400 44000
rect 207240 44000 207400 44160
rect 207240 44160 207400 44320
rect 207240 44320 207400 44480
rect 207240 47680 207400 47840
rect 207240 47840 207400 48000
rect 207240 48000 207400 48160
rect 207240 48160 207400 48320
rect 207240 48320 207400 48480
rect 207240 48480 207400 48640
rect 207240 48640 207400 48800
rect 207240 48800 207400 48960
rect 207240 48960 207400 49120
rect 207240 49120 207400 49280
rect 207240 49280 207400 49440
rect 207240 49440 207400 49600
rect 207240 49600 207400 49760
rect 207240 49760 207400 49920
rect 207240 49920 207400 50080
rect 207240 50080 207400 50240
rect 207240 50240 207400 50400
rect 207240 50400 207400 50560
rect 207240 50560 207400 50720
rect 207240 50720 207400 50880
rect 207240 50880 207400 51040
rect 207240 51040 207400 51200
rect 207240 51200 207400 51360
rect 207240 51360 207400 51520
rect 207240 51520 207400 51680
rect 207240 51680 207400 51840
rect 207240 51840 207400 52000
rect 207240 52000 207400 52160
rect 207240 52160 207400 52320
rect 207240 52320 207400 52480
rect 207240 52480 207400 52640
rect 207240 52640 207400 52800
rect 207240 52800 207400 52960
rect 207240 52960 207400 53120
rect 207240 53120 207400 53280
rect 207240 53280 207400 53440
rect 207240 53440 207400 53600
rect 207240 53600 207400 53760
rect 207400 25920 207560 26080
rect 207400 26080 207560 26240
rect 207400 26240 207560 26400
rect 207400 26400 207560 26560
rect 207400 26560 207560 26720
rect 207400 26720 207560 26880
rect 207400 26880 207560 27040
rect 207400 27040 207560 27200
rect 207400 27200 207560 27360
rect 207400 27360 207560 27520
rect 207400 27520 207560 27680
rect 207400 27680 207560 27840
rect 207400 27840 207560 28000
rect 207400 28000 207560 28160
rect 207400 28160 207560 28320
rect 207400 28320 207560 28480
rect 207400 28480 207560 28640
rect 207400 28640 207560 28800
rect 207400 28800 207560 28960
rect 207400 28960 207560 29120
rect 207400 29120 207560 29280
rect 207400 29280 207560 29440
rect 207400 29440 207560 29600
rect 207400 29600 207560 29760
rect 207400 29760 207560 29920
rect 207400 29920 207560 30080
rect 207400 30080 207560 30240
rect 207400 30240 207560 30400
rect 207400 30400 207560 30560
rect 207400 30560 207560 30720
rect 207400 30720 207560 30880
rect 207400 30880 207560 31040
rect 207400 31040 207560 31200
rect 207400 31200 207560 31360
rect 207400 31360 207560 31520
rect 207400 31520 207560 31680
rect 207400 31680 207560 31840
rect 207400 31840 207560 32000
rect 207400 32000 207560 32160
rect 207400 32160 207560 32320
rect 207400 32320 207560 32480
rect 207400 32480 207560 32640
rect 207400 32640 207560 32800
rect 207400 32800 207560 32960
rect 207400 32960 207560 33120
rect 207400 33120 207560 33280
rect 207400 33280 207560 33440
rect 207400 33440 207560 33600
rect 207400 33600 207560 33760
rect 207400 33760 207560 33920
rect 207400 33920 207560 34080
rect 207400 34080 207560 34240
rect 207400 34240 207560 34400
rect 207400 34400 207560 34560
rect 207400 34560 207560 34720
rect 207400 34720 207560 34880
rect 207400 34880 207560 35040
rect 207400 35040 207560 35200
rect 207400 35200 207560 35360
rect 207400 35360 207560 35520
rect 207400 35520 207560 35680
rect 207400 35680 207560 35840
rect 207400 35840 207560 36000
rect 207400 36000 207560 36160
rect 207400 36160 207560 36320
rect 207400 36320 207560 36480
rect 207400 36480 207560 36640
rect 207400 36640 207560 36800
rect 207400 36800 207560 36960
rect 207400 36960 207560 37120
rect 207400 37120 207560 37280
rect 207400 37280 207560 37440
rect 207400 37440 207560 37600
rect 207400 37600 207560 37760
rect 207400 37760 207560 37920
rect 207400 37920 207560 38080
rect 207400 38080 207560 38240
rect 207400 38240 207560 38400
rect 207400 38400 207560 38560
rect 207400 38560 207560 38720
rect 207400 38720 207560 38880
rect 207400 38880 207560 39040
rect 207400 39040 207560 39200
rect 207400 39200 207560 39360
rect 207400 39360 207560 39520
rect 207400 39520 207560 39680
rect 207400 39680 207560 39840
rect 207400 39840 207560 40000
rect 207400 40000 207560 40160
rect 207400 40160 207560 40320
rect 207400 40320 207560 40480
rect 207400 40480 207560 40640
rect 207400 40640 207560 40800
rect 207400 40800 207560 40960
rect 207400 40960 207560 41120
rect 207400 41120 207560 41280
rect 207400 41280 207560 41440
rect 207400 41440 207560 41600
rect 207400 41600 207560 41760
rect 207400 41760 207560 41920
rect 207400 41920 207560 42080
rect 207400 42080 207560 42240
rect 207400 42240 207560 42400
rect 207400 42400 207560 42560
rect 207400 42560 207560 42720
rect 207400 42720 207560 42880
rect 207400 42880 207560 43040
rect 207400 43040 207560 43200
rect 207400 43200 207560 43360
rect 207400 43360 207560 43520
rect 207400 43520 207560 43680
rect 207400 43680 207560 43840
rect 207400 43840 207560 44000
rect 207400 44000 207560 44160
rect 207400 44160 207560 44320
rect 207400 44320 207560 44480
rect 207400 44480 207560 44640
rect 207400 47520 207560 47680
rect 207400 47680 207560 47840
rect 207400 47840 207560 48000
rect 207400 48000 207560 48160
rect 207400 48160 207560 48320
rect 207400 48320 207560 48480
rect 207400 48480 207560 48640
rect 207400 48640 207560 48800
rect 207400 48800 207560 48960
rect 207400 48960 207560 49120
rect 207400 49120 207560 49280
rect 207400 49280 207560 49440
rect 207400 49440 207560 49600
rect 207400 49600 207560 49760
rect 207400 49760 207560 49920
rect 207400 49920 207560 50080
rect 207400 50080 207560 50240
rect 207400 50240 207560 50400
rect 207400 50400 207560 50560
rect 207400 50560 207560 50720
rect 207400 50720 207560 50880
rect 207400 50880 207560 51040
rect 207400 51040 207560 51200
rect 207400 51200 207560 51360
rect 207400 51360 207560 51520
rect 207400 51520 207560 51680
rect 207400 51680 207560 51840
rect 207400 51840 207560 52000
rect 207400 52000 207560 52160
rect 207400 52160 207560 52320
rect 207400 52320 207560 52480
rect 207400 52480 207560 52640
rect 207400 52640 207560 52800
rect 207400 52800 207560 52960
rect 207400 52960 207560 53120
rect 207400 53120 207560 53280
rect 207400 53280 207560 53440
rect 207400 53440 207560 53600
rect 207400 53600 207560 53760
rect 207400 53760 207560 53920
rect 207560 25920 207720 26080
rect 207560 26080 207720 26240
rect 207560 26240 207720 26400
rect 207560 26400 207720 26560
rect 207560 26560 207720 26720
rect 207560 26720 207720 26880
rect 207560 26880 207720 27040
rect 207560 27040 207720 27200
rect 207560 27200 207720 27360
rect 207560 27360 207720 27520
rect 207560 27520 207720 27680
rect 207560 27680 207720 27840
rect 207560 27840 207720 28000
rect 207560 28000 207720 28160
rect 207560 28160 207720 28320
rect 207560 28320 207720 28480
rect 207560 28480 207720 28640
rect 207560 28640 207720 28800
rect 207560 28800 207720 28960
rect 207560 28960 207720 29120
rect 207560 29120 207720 29280
rect 207560 29280 207720 29440
rect 207560 29440 207720 29600
rect 207560 29600 207720 29760
rect 207560 29760 207720 29920
rect 207560 29920 207720 30080
rect 207560 30080 207720 30240
rect 207560 30240 207720 30400
rect 207560 30400 207720 30560
rect 207560 30560 207720 30720
rect 207560 30720 207720 30880
rect 207560 30880 207720 31040
rect 207560 31040 207720 31200
rect 207560 31200 207720 31360
rect 207560 31360 207720 31520
rect 207560 31520 207720 31680
rect 207560 31680 207720 31840
rect 207560 31840 207720 32000
rect 207560 32000 207720 32160
rect 207560 32160 207720 32320
rect 207560 32320 207720 32480
rect 207560 32480 207720 32640
rect 207560 32640 207720 32800
rect 207560 32800 207720 32960
rect 207560 32960 207720 33120
rect 207560 33120 207720 33280
rect 207560 33280 207720 33440
rect 207560 33440 207720 33600
rect 207560 33600 207720 33760
rect 207560 33760 207720 33920
rect 207560 33920 207720 34080
rect 207560 34080 207720 34240
rect 207560 34240 207720 34400
rect 207560 34400 207720 34560
rect 207560 34560 207720 34720
rect 207560 34720 207720 34880
rect 207560 34880 207720 35040
rect 207560 35040 207720 35200
rect 207560 35200 207720 35360
rect 207560 35360 207720 35520
rect 207560 35520 207720 35680
rect 207560 35680 207720 35840
rect 207560 35840 207720 36000
rect 207560 36000 207720 36160
rect 207560 36160 207720 36320
rect 207560 36320 207720 36480
rect 207560 36480 207720 36640
rect 207560 36640 207720 36800
rect 207560 36800 207720 36960
rect 207560 36960 207720 37120
rect 207560 37120 207720 37280
rect 207560 37280 207720 37440
rect 207560 37440 207720 37600
rect 207560 37600 207720 37760
rect 207560 37760 207720 37920
rect 207560 37920 207720 38080
rect 207560 38080 207720 38240
rect 207560 38240 207720 38400
rect 207560 38400 207720 38560
rect 207560 38560 207720 38720
rect 207560 38720 207720 38880
rect 207560 38880 207720 39040
rect 207560 39040 207720 39200
rect 207560 39200 207720 39360
rect 207560 39360 207720 39520
rect 207560 39520 207720 39680
rect 207560 39680 207720 39840
rect 207560 39840 207720 40000
rect 207560 40000 207720 40160
rect 207560 40160 207720 40320
rect 207560 40320 207720 40480
rect 207560 40480 207720 40640
rect 207560 40640 207720 40800
rect 207560 40800 207720 40960
rect 207560 40960 207720 41120
rect 207560 41120 207720 41280
rect 207560 41280 207720 41440
rect 207560 41440 207720 41600
rect 207560 41600 207720 41760
rect 207560 41760 207720 41920
rect 207560 41920 207720 42080
rect 207560 42080 207720 42240
rect 207560 42240 207720 42400
rect 207560 42400 207720 42560
rect 207560 42560 207720 42720
rect 207560 42720 207720 42880
rect 207560 42880 207720 43040
rect 207560 43040 207720 43200
rect 207560 43200 207720 43360
rect 207560 43360 207720 43520
rect 207560 43520 207720 43680
rect 207560 43680 207720 43840
rect 207560 43840 207720 44000
rect 207560 44000 207720 44160
rect 207560 44160 207720 44320
rect 207560 44320 207720 44480
rect 207560 44480 207720 44640
rect 207560 44640 207720 44800
rect 207560 47520 207720 47680
rect 207560 47680 207720 47840
rect 207560 47840 207720 48000
rect 207560 48000 207720 48160
rect 207560 48160 207720 48320
rect 207560 48320 207720 48480
rect 207560 48480 207720 48640
rect 207560 48640 207720 48800
rect 207560 48800 207720 48960
rect 207560 48960 207720 49120
rect 207560 49120 207720 49280
rect 207560 49280 207720 49440
rect 207560 49440 207720 49600
rect 207560 49600 207720 49760
rect 207560 49760 207720 49920
rect 207560 49920 207720 50080
rect 207560 50080 207720 50240
rect 207560 50240 207720 50400
rect 207560 50400 207720 50560
rect 207560 50560 207720 50720
rect 207560 50720 207720 50880
rect 207560 50880 207720 51040
rect 207560 51040 207720 51200
rect 207560 51200 207720 51360
rect 207560 51360 207720 51520
rect 207560 51520 207720 51680
rect 207560 51680 207720 51840
rect 207560 51840 207720 52000
rect 207560 52000 207720 52160
rect 207560 52160 207720 52320
rect 207560 52320 207720 52480
rect 207560 52480 207720 52640
rect 207560 52640 207720 52800
rect 207560 52800 207720 52960
rect 207560 52960 207720 53120
rect 207560 53120 207720 53280
rect 207560 53280 207720 53440
rect 207560 53440 207720 53600
rect 207560 53600 207720 53760
rect 207560 53760 207720 53920
rect 207560 53920 207720 54080
rect 207720 25920 207880 26080
rect 207720 26080 207880 26240
rect 207720 26240 207880 26400
rect 207720 26400 207880 26560
rect 207720 26560 207880 26720
rect 207720 26720 207880 26880
rect 207720 26880 207880 27040
rect 207720 27040 207880 27200
rect 207720 27200 207880 27360
rect 207720 27360 207880 27520
rect 207720 27520 207880 27680
rect 207720 27680 207880 27840
rect 207720 27840 207880 28000
rect 207720 28000 207880 28160
rect 207720 28160 207880 28320
rect 207720 28320 207880 28480
rect 207720 28480 207880 28640
rect 207720 28640 207880 28800
rect 207720 28800 207880 28960
rect 207720 28960 207880 29120
rect 207720 29120 207880 29280
rect 207720 29280 207880 29440
rect 207720 29440 207880 29600
rect 207720 29600 207880 29760
rect 207720 29760 207880 29920
rect 207720 29920 207880 30080
rect 207720 30080 207880 30240
rect 207720 30240 207880 30400
rect 207720 30400 207880 30560
rect 207720 30560 207880 30720
rect 207720 30720 207880 30880
rect 207720 30880 207880 31040
rect 207720 31040 207880 31200
rect 207720 31200 207880 31360
rect 207720 31360 207880 31520
rect 207720 31520 207880 31680
rect 207720 31680 207880 31840
rect 207720 31840 207880 32000
rect 207720 32000 207880 32160
rect 207720 32160 207880 32320
rect 207720 32320 207880 32480
rect 207720 32480 207880 32640
rect 207720 32640 207880 32800
rect 207720 32800 207880 32960
rect 207720 32960 207880 33120
rect 207720 33120 207880 33280
rect 207720 33280 207880 33440
rect 207720 33440 207880 33600
rect 207720 33600 207880 33760
rect 207720 33760 207880 33920
rect 207720 33920 207880 34080
rect 207720 34080 207880 34240
rect 207720 34240 207880 34400
rect 207720 34400 207880 34560
rect 207720 34560 207880 34720
rect 207720 34720 207880 34880
rect 207720 34880 207880 35040
rect 207720 35040 207880 35200
rect 207720 35200 207880 35360
rect 207720 35360 207880 35520
rect 207720 35520 207880 35680
rect 207720 35680 207880 35840
rect 207720 35840 207880 36000
rect 207720 36000 207880 36160
rect 207720 36160 207880 36320
rect 207720 36320 207880 36480
rect 207720 36480 207880 36640
rect 207720 36640 207880 36800
rect 207720 36800 207880 36960
rect 207720 36960 207880 37120
rect 207720 37120 207880 37280
rect 207720 37280 207880 37440
rect 207720 37440 207880 37600
rect 207720 37600 207880 37760
rect 207720 37760 207880 37920
rect 207720 37920 207880 38080
rect 207720 38080 207880 38240
rect 207720 38240 207880 38400
rect 207720 38400 207880 38560
rect 207720 38560 207880 38720
rect 207720 38720 207880 38880
rect 207720 38880 207880 39040
rect 207720 39040 207880 39200
rect 207720 39200 207880 39360
rect 207720 39360 207880 39520
rect 207720 39520 207880 39680
rect 207720 39680 207880 39840
rect 207720 39840 207880 40000
rect 207720 40000 207880 40160
rect 207720 40160 207880 40320
rect 207720 40320 207880 40480
rect 207720 40480 207880 40640
rect 207720 40640 207880 40800
rect 207720 40800 207880 40960
rect 207720 40960 207880 41120
rect 207720 41120 207880 41280
rect 207720 41280 207880 41440
rect 207720 41440 207880 41600
rect 207720 41600 207880 41760
rect 207720 41760 207880 41920
rect 207720 41920 207880 42080
rect 207720 42080 207880 42240
rect 207720 42240 207880 42400
rect 207720 42400 207880 42560
rect 207720 42560 207880 42720
rect 207720 42720 207880 42880
rect 207720 42880 207880 43040
rect 207720 43040 207880 43200
rect 207720 43200 207880 43360
rect 207720 43360 207880 43520
rect 207720 43520 207880 43680
rect 207720 43680 207880 43840
rect 207720 43840 207880 44000
rect 207720 44000 207880 44160
rect 207720 44160 207880 44320
rect 207720 44320 207880 44480
rect 207720 44480 207880 44640
rect 207720 44640 207880 44800
rect 207720 44800 207880 44960
rect 207720 47360 207880 47520
rect 207720 47520 207880 47680
rect 207720 47680 207880 47840
rect 207720 47840 207880 48000
rect 207720 48000 207880 48160
rect 207720 48160 207880 48320
rect 207720 48320 207880 48480
rect 207720 48480 207880 48640
rect 207720 48640 207880 48800
rect 207720 48800 207880 48960
rect 207720 48960 207880 49120
rect 207720 49120 207880 49280
rect 207720 49280 207880 49440
rect 207720 49440 207880 49600
rect 207720 49600 207880 49760
rect 207720 49760 207880 49920
rect 207720 49920 207880 50080
rect 207720 50080 207880 50240
rect 207720 50240 207880 50400
rect 207720 50400 207880 50560
rect 207720 50560 207880 50720
rect 207720 50720 207880 50880
rect 207720 50880 207880 51040
rect 207720 51040 207880 51200
rect 207720 51200 207880 51360
rect 207720 51360 207880 51520
rect 207720 51520 207880 51680
rect 207720 51680 207880 51840
rect 207720 51840 207880 52000
rect 207720 52000 207880 52160
rect 207720 52160 207880 52320
rect 207720 52320 207880 52480
rect 207720 52480 207880 52640
rect 207720 52640 207880 52800
rect 207720 52800 207880 52960
rect 207720 52960 207880 53120
rect 207720 53120 207880 53280
rect 207720 53280 207880 53440
rect 207720 53440 207880 53600
rect 207720 53600 207880 53760
rect 207720 53760 207880 53920
rect 207720 53920 207880 54080
rect 207720 54080 207880 54240
rect 207880 25920 208040 26080
rect 207880 26080 208040 26240
rect 207880 26240 208040 26400
rect 207880 26400 208040 26560
rect 207880 26560 208040 26720
rect 207880 26720 208040 26880
rect 207880 26880 208040 27040
rect 207880 27040 208040 27200
rect 207880 27200 208040 27360
rect 207880 27360 208040 27520
rect 207880 27520 208040 27680
rect 207880 27680 208040 27840
rect 207880 27840 208040 28000
rect 207880 28000 208040 28160
rect 207880 28160 208040 28320
rect 207880 28320 208040 28480
rect 207880 28480 208040 28640
rect 207880 28640 208040 28800
rect 207880 28800 208040 28960
rect 207880 28960 208040 29120
rect 207880 29120 208040 29280
rect 207880 29280 208040 29440
rect 207880 29440 208040 29600
rect 207880 29600 208040 29760
rect 207880 29760 208040 29920
rect 207880 29920 208040 30080
rect 207880 30080 208040 30240
rect 207880 30240 208040 30400
rect 207880 30400 208040 30560
rect 207880 30560 208040 30720
rect 207880 30720 208040 30880
rect 207880 30880 208040 31040
rect 207880 31040 208040 31200
rect 207880 31200 208040 31360
rect 207880 31360 208040 31520
rect 207880 31520 208040 31680
rect 207880 31680 208040 31840
rect 207880 31840 208040 32000
rect 207880 32000 208040 32160
rect 207880 32160 208040 32320
rect 207880 32320 208040 32480
rect 207880 32480 208040 32640
rect 207880 32640 208040 32800
rect 207880 32800 208040 32960
rect 207880 32960 208040 33120
rect 207880 33120 208040 33280
rect 207880 33280 208040 33440
rect 207880 33440 208040 33600
rect 207880 33600 208040 33760
rect 207880 33760 208040 33920
rect 207880 33920 208040 34080
rect 207880 34080 208040 34240
rect 207880 34240 208040 34400
rect 207880 34400 208040 34560
rect 207880 34560 208040 34720
rect 207880 34720 208040 34880
rect 207880 34880 208040 35040
rect 207880 35040 208040 35200
rect 207880 35200 208040 35360
rect 207880 35360 208040 35520
rect 207880 35520 208040 35680
rect 207880 35680 208040 35840
rect 207880 35840 208040 36000
rect 207880 36000 208040 36160
rect 207880 36160 208040 36320
rect 207880 36320 208040 36480
rect 207880 36480 208040 36640
rect 207880 36640 208040 36800
rect 207880 36800 208040 36960
rect 207880 36960 208040 37120
rect 207880 37120 208040 37280
rect 207880 37280 208040 37440
rect 207880 37440 208040 37600
rect 207880 37600 208040 37760
rect 207880 37760 208040 37920
rect 207880 37920 208040 38080
rect 207880 38080 208040 38240
rect 207880 38240 208040 38400
rect 207880 38400 208040 38560
rect 207880 38560 208040 38720
rect 207880 38720 208040 38880
rect 207880 38880 208040 39040
rect 207880 39040 208040 39200
rect 207880 39200 208040 39360
rect 207880 39360 208040 39520
rect 207880 39520 208040 39680
rect 207880 39680 208040 39840
rect 207880 39840 208040 40000
rect 207880 40000 208040 40160
rect 207880 40160 208040 40320
rect 207880 40320 208040 40480
rect 207880 40480 208040 40640
rect 207880 40640 208040 40800
rect 207880 40800 208040 40960
rect 207880 40960 208040 41120
rect 207880 41120 208040 41280
rect 207880 41280 208040 41440
rect 207880 41440 208040 41600
rect 207880 41600 208040 41760
rect 207880 41760 208040 41920
rect 207880 41920 208040 42080
rect 207880 42080 208040 42240
rect 207880 42240 208040 42400
rect 207880 42400 208040 42560
rect 207880 42560 208040 42720
rect 207880 42720 208040 42880
rect 207880 42880 208040 43040
rect 207880 43040 208040 43200
rect 207880 43200 208040 43360
rect 207880 43360 208040 43520
rect 207880 43520 208040 43680
rect 207880 43680 208040 43840
rect 207880 43840 208040 44000
rect 207880 44000 208040 44160
rect 207880 44160 208040 44320
rect 207880 44320 208040 44480
rect 207880 44480 208040 44640
rect 207880 44640 208040 44800
rect 207880 44800 208040 44960
rect 207880 44960 208040 45120
rect 207880 47360 208040 47520
rect 207880 47520 208040 47680
rect 207880 47680 208040 47840
rect 207880 47840 208040 48000
rect 207880 48000 208040 48160
rect 207880 48160 208040 48320
rect 207880 48320 208040 48480
rect 207880 48480 208040 48640
rect 207880 48640 208040 48800
rect 207880 48800 208040 48960
rect 207880 48960 208040 49120
rect 207880 49120 208040 49280
rect 207880 49280 208040 49440
rect 207880 49440 208040 49600
rect 207880 49600 208040 49760
rect 207880 49760 208040 49920
rect 207880 49920 208040 50080
rect 207880 50080 208040 50240
rect 207880 50240 208040 50400
rect 207880 50400 208040 50560
rect 207880 50560 208040 50720
rect 207880 50720 208040 50880
rect 207880 50880 208040 51040
rect 207880 51040 208040 51200
rect 207880 51200 208040 51360
rect 207880 51360 208040 51520
rect 207880 51520 208040 51680
rect 207880 51680 208040 51840
rect 207880 51840 208040 52000
rect 207880 52000 208040 52160
rect 207880 52160 208040 52320
rect 207880 52320 208040 52480
rect 207880 52480 208040 52640
rect 207880 52640 208040 52800
rect 207880 52800 208040 52960
rect 207880 52960 208040 53120
rect 207880 53120 208040 53280
rect 207880 53280 208040 53440
rect 207880 53440 208040 53600
rect 207880 53600 208040 53760
rect 207880 53760 208040 53920
rect 207880 53920 208040 54080
rect 207880 54080 208040 54240
rect 208040 26080 208200 26240
rect 208040 26240 208200 26400
rect 208040 26400 208200 26560
rect 208040 26560 208200 26720
rect 208040 26720 208200 26880
rect 208040 26880 208200 27040
rect 208040 27040 208200 27200
rect 208040 27200 208200 27360
rect 208040 27360 208200 27520
rect 208040 27520 208200 27680
rect 208040 27680 208200 27840
rect 208040 27840 208200 28000
rect 208040 28000 208200 28160
rect 208040 28160 208200 28320
rect 208040 28320 208200 28480
rect 208040 28480 208200 28640
rect 208040 28640 208200 28800
rect 208040 28800 208200 28960
rect 208040 28960 208200 29120
rect 208040 29120 208200 29280
rect 208040 29280 208200 29440
rect 208040 29440 208200 29600
rect 208040 29600 208200 29760
rect 208040 29760 208200 29920
rect 208040 29920 208200 30080
rect 208040 30080 208200 30240
rect 208040 30240 208200 30400
rect 208040 30400 208200 30560
rect 208040 30560 208200 30720
rect 208040 30720 208200 30880
rect 208040 30880 208200 31040
rect 208040 31040 208200 31200
rect 208040 31200 208200 31360
rect 208040 31360 208200 31520
rect 208040 31520 208200 31680
rect 208040 31680 208200 31840
rect 208040 31840 208200 32000
rect 208040 32000 208200 32160
rect 208040 32160 208200 32320
rect 208040 32320 208200 32480
rect 208040 32480 208200 32640
rect 208040 32640 208200 32800
rect 208040 32800 208200 32960
rect 208040 32960 208200 33120
rect 208040 33120 208200 33280
rect 208040 33280 208200 33440
rect 208040 33440 208200 33600
rect 208040 33600 208200 33760
rect 208040 33760 208200 33920
rect 208040 33920 208200 34080
rect 208040 34080 208200 34240
rect 208040 34240 208200 34400
rect 208040 34400 208200 34560
rect 208040 34560 208200 34720
rect 208040 34720 208200 34880
rect 208040 34880 208200 35040
rect 208040 35040 208200 35200
rect 208040 35200 208200 35360
rect 208040 35360 208200 35520
rect 208040 35520 208200 35680
rect 208040 35680 208200 35840
rect 208040 35840 208200 36000
rect 208040 36000 208200 36160
rect 208040 36160 208200 36320
rect 208040 36320 208200 36480
rect 208040 36480 208200 36640
rect 208040 36640 208200 36800
rect 208040 36800 208200 36960
rect 208040 36960 208200 37120
rect 208040 37120 208200 37280
rect 208040 37280 208200 37440
rect 208040 37440 208200 37600
rect 208040 37600 208200 37760
rect 208040 37760 208200 37920
rect 208040 37920 208200 38080
rect 208040 38080 208200 38240
rect 208040 38240 208200 38400
rect 208040 38400 208200 38560
rect 208040 38560 208200 38720
rect 208040 38720 208200 38880
rect 208040 38880 208200 39040
rect 208040 39040 208200 39200
rect 208040 39200 208200 39360
rect 208040 39360 208200 39520
rect 208040 39520 208200 39680
rect 208040 39680 208200 39840
rect 208040 39840 208200 40000
rect 208040 40000 208200 40160
rect 208040 40160 208200 40320
rect 208040 40320 208200 40480
rect 208040 40480 208200 40640
rect 208040 40640 208200 40800
rect 208040 40800 208200 40960
rect 208040 40960 208200 41120
rect 208040 41120 208200 41280
rect 208040 41280 208200 41440
rect 208040 41440 208200 41600
rect 208040 41600 208200 41760
rect 208040 41760 208200 41920
rect 208040 41920 208200 42080
rect 208040 42080 208200 42240
rect 208040 42240 208200 42400
rect 208040 42400 208200 42560
rect 208040 42560 208200 42720
rect 208040 42720 208200 42880
rect 208040 42880 208200 43040
rect 208040 43040 208200 43200
rect 208040 43200 208200 43360
rect 208040 43360 208200 43520
rect 208040 43520 208200 43680
rect 208040 43680 208200 43840
rect 208040 43840 208200 44000
rect 208040 44000 208200 44160
rect 208040 44160 208200 44320
rect 208040 44320 208200 44480
rect 208040 44480 208200 44640
rect 208040 44640 208200 44800
rect 208040 44800 208200 44960
rect 208040 44960 208200 45120
rect 208040 45120 208200 45280
rect 208040 47200 208200 47360
rect 208040 47360 208200 47520
rect 208040 47520 208200 47680
rect 208040 47680 208200 47840
rect 208040 47840 208200 48000
rect 208040 48000 208200 48160
rect 208040 48160 208200 48320
rect 208040 48320 208200 48480
rect 208040 48480 208200 48640
rect 208040 48640 208200 48800
rect 208040 48800 208200 48960
rect 208040 48960 208200 49120
rect 208040 49120 208200 49280
rect 208040 49280 208200 49440
rect 208040 49440 208200 49600
rect 208040 49600 208200 49760
rect 208040 49760 208200 49920
rect 208040 49920 208200 50080
rect 208040 50080 208200 50240
rect 208040 50240 208200 50400
rect 208040 50400 208200 50560
rect 208040 50560 208200 50720
rect 208040 50720 208200 50880
rect 208040 50880 208200 51040
rect 208040 51040 208200 51200
rect 208040 51200 208200 51360
rect 208040 51360 208200 51520
rect 208040 51520 208200 51680
rect 208040 51680 208200 51840
rect 208040 51840 208200 52000
rect 208040 52000 208200 52160
rect 208040 52160 208200 52320
rect 208040 52320 208200 52480
rect 208040 52480 208200 52640
rect 208040 52640 208200 52800
rect 208040 52800 208200 52960
rect 208040 52960 208200 53120
rect 208040 53120 208200 53280
rect 208040 53280 208200 53440
rect 208040 53440 208200 53600
rect 208040 53600 208200 53760
rect 208040 53760 208200 53920
rect 208040 53920 208200 54080
rect 208040 54080 208200 54240
rect 208040 54240 208200 54400
rect 208200 26080 208360 26240
rect 208200 26240 208360 26400
rect 208200 26400 208360 26560
rect 208200 26560 208360 26720
rect 208200 26720 208360 26880
rect 208200 26880 208360 27040
rect 208200 27040 208360 27200
rect 208200 27200 208360 27360
rect 208200 27360 208360 27520
rect 208200 27520 208360 27680
rect 208200 27680 208360 27840
rect 208200 27840 208360 28000
rect 208200 28000 208360 28160
rect 208200 28160 208360 28320
rect 208200 28320 208360 28480
rect 208200 28480 208360 28640
rect 208200 28640 208360 28800
rect 208200 28800 208360 28960
rect 208200 28960 208360 29120
rect 208200 29120 208360 29280
rect 208200 29280 208360 29440
rect 208200 29440 208360 29600
rect 208200 29600 208360 29760
rect 208200 29760 208360 29920
rect 208200 29920 208360 30080
rect 208200 30080 208360 30240
rect 208200 30240 208360 30400
rect 208200 30400 208360 30560
rect 208200 30560 208360 30720
rect 208200 30720 208360 30880
rect 208200 30880 208360 31040
rect 208200 31040 208360 31200
rect 208200 31200 208360 31360
rect 208200 31360 208360 31520
rect 208200 31520 208360 31680
rect 208200 31680 208360 31840
rect 208200 31840 208360 32000
rect 208200 32000 208360 32160
rect 208200 32160 208360 32320
rect 208200 32320 208360 32480
rect 208200 32480 208360 32640
rect 208200 32640 208360 32800
rect 208200 32800 208360 32960
rect 208200 32960 208360 33120
rect 208200 33120 208360 33280
rect 208200 33280 208360 33440
rect 208200 33440 208360 33600
rect 208200 33600 208360 33760
rect 208200 33760 208360 33920
rect 208200 33920 208360 34080
rect 208200 34080 208360 34240
rect 208200 34240 208360 34400
rect 208200 34400 208360 34560
rect 208200 34560 208360 34720
rect 208200 34720 208360 34880
rect 208200 34880 208360 35040
rect 208200 35040 208360 35200
rect 208200 35200 208360 35360
rect 208200 35360 208360 35520
rect 208200 35520 208360 35680
rect 208200 35680 208360 35840
rect 208200 35840 208360 36000
rect 208200 36000 208360 36160
rect 208200 36160 208360 36320
rect 208200 36320 208360 36480
rect 208200 36480 208360 36640
rect 208200 36640 208360 36800
rect 208200 36800 208360 36960
rect 208200 36960 208360 37120
rect 208200 37120 208360 37280
rect 208200 37280 208360 37440
rect 208200 37440 208360 37600
rect 208200 37600 208360 37760
rect 208200 37760 208360 37920
rect 208200 37920 208360 38080
rect 208200 38080 208360 38240
rect 208200 38240 208360 38400
rect 208200 38400 208360 38560
rect 208200 38560 208360 38720
rect 208200 38720 208360 38880
rect 208200 38880 208360 39040
rect 208200 39040 208360 39200
rect 208200 39200 208360 39360
rect 208200 39360 208360 39520
rect 208200 39520 208360 39680
rect 208200 39680 208360 39840
rect 208200 39840 208360 40000
rect 208200 40000 208360 40160
rect 208200 40160 208360 40320
rect 208200 40320 208360 40480
rect 208200 40480 208360 40640
rect 208200 40640 208360 40800
rect 208200 40800 208360 40960
rect 208200 40960 208360 41120
rect 208200 41120 208360 41280
rect 208200 41280 208360 41440
rect 208200 41440 208360 41600
rect 208200 41600 208360 41760
rect 208200 41760 208360 41920
rect 208200 41920 208360 42080
rect 208200 42080 208360 42240
rect 208200 42240 208360 42400
rect 208200 42400 208360 42560
rect 208200 42560 208360 42720
rect 208200 42720 208360 42880
rect 208200 42880 208360 43040
rect 208200 43040 208360 43200
rect 208200 43200 208360 43360
rect 208200 43360 208360 43520
rect 208200 43520 208360 43680
rect 208200 43680 208360 43840
rect 208200 43840 208360 44000
rect 208200 44000 208360 44160
rect 208200 44160 208360 44320
rect 208200 44320 208360 44480
rect 208200 44480 208360 44640
rect 208200 44640 208360 44800
rect 208200 44800 208360 44960
rect 208200 44960 208360 45120
rect 208200 45120 208360 45280
rect 208200 45280 208360 45440
rect 208200 47200 208360 47360
rect 208200 47360 208360 47520
rect 208200 47520 208360 47680
rect 208200 47680 208360 47840
rect 208200 47840 208360 48000
rect 208200 48000 208360 48160
rect 208200 48160 208360 48320
rect 208200 48320 208360 48480
rect 208200 48480 208360 48640
rect 208200 48640 208360 48800
rect 208200 48800 208360 48960
rect 208200 48960 208360 49120
rect 208200 49120 208360 49280
rect 208200 49280 208360 49440
rect 208200 49440 208360 49600
rect 208200 49600 208360 49760
rect 208200 49760 208360 49920
rect 208200 49920 208360 50080
rect 208200 50080 208360 50240
rect 208200 50240 208360 50400
rect 208200 50400 208360 50560
rect 208200 50560 208360 50720
rect 208200 50720 208360 50880
rect 208200 50880 208360 51040
rect 208200 51040 208360 51200
rect 208200 51200 208360 51360
rect 208200 51360 208360 51520
rect 208200 51520 208360 51680
rect 208200 51680 208360 51840
rect 208200 51840 208360 52000
rect 208200 52000 208360 52160
rect 208200 52160 208360 52320
rect 208200 52320 208360 52480
rect 208200 52480 208360 52640
rect 208200 52640 208360 52800
rect 208200 52800 208360 52960
rect 208200 52960 208360 53120
rect 208200 53120 208360 53280
rect 208200 53280 208360 53440
rect 208200 53440 208360 53600
rect 208200 53600 208360 53760
rect 208200 53760 208360 53920
rect 208200 53920 208360 54080
rect 208200 54080 208360 54240
rect 208200 54240 208360 54400
rect 208360 26240 208520 26400
rect 208360 26400 208520 26560
rect 208360 26560 208520 26720
rect 208360 26720 208520 26880
rect 208360 26880 208520 27040
rect 208360 27040 208520 27200
rect 208360 27200 208520 27360
rect 208360 27360 208520 27520
rect 208360 27520 208520 27680
rect 208360 27680 208520 27840
rect 208360 27840 208520 28000
rect 208360 28000 208520 28160
rect 208360 28160 208520 28320
rect 208360 28320 208520 28480
rect 208360 28480 208520 28640
rect 208360 28640 208520 28800
rect 208360 28800 208520 28960
rect 208360 28960 208520 29120
rect 208360 29120 208520 29280
rect 208360 29280 208520 29440
rect 208360 29440 208520 29600
rect 208360 29600 208520 29760
rect 208360 29760 208520 29920
rect 208360 29920 208520 30080
rect 208360 30080 208520 30240
rect 208360 30240 208520 30400
rect 208360 30400 208520 30560
rect 208360 30560 208520 30720
rect 208360 30720 208520 30880
rect 208360 30880 208520 31040
rect 208360 31040 208520 31200
rect 208360 31200 208520 31360
rect 208360 31360 208520 31520
rect 208360 31520 208520 31680
rect 208360 31680 208520 31840
rect 208360 31840 208520 32000
rect 208360 32000 208520 32160
rect 208360 32160 208520 32320
rect 208360 32320 208520 32480
rect 208360 32480 208520 32640
rect 208360 32640 208520 32800
rect 208360 32800 208520 32960
rect 208360 32960 208520 33120
rect 208360 33120 208520 33280
rect 208360 33280 208520 33440
rect 208360 33440 208520 33600
rect 208360 33600 208520 33760
rect 208360 33760 208520 33920
rect 208360 33920 208520 34080
rect 208360 34080 208520 34240
rect 208360 34240 208520 34400
rect 208360 34400 208520 34560
rect 208360 34560 208520 34720
rect 208360 34720 208520 34880
rect 208360 34880 208520 35040
rect 208360 35040 208520 35200
rect 208360 35200 208520 35360
rect 208360 35360 208520 35520
rect 208360 35520 208520 35680
rect 208360 35680 208520 35840
rect 208360 35840 208520 36000
rect 208360 36000 208520 36160
rect 208360 36160 208520 36320
rect 208360 36320 208520 36480
rect 208360 36480 208520 36640
rect 208360 36640 208520 36800
rect 208360 36800 208520 36960
rect 208360 36960 208520 37120
rect 208360 37120 208520 37280
rect 208360 37280 208520 37440
rect 208360 37440 208520 37600
rect 208360 37600 208520 37760
rect 208360 37760 208520 37920
rect 208360 37920 208520 38080
rect 208360 38080 208520 38240
rect 208360 38240 208520 38400
rect 208360 38400 208520 38560
rect 208360 38560 208520 38720
rect 208360 38720 208520 38880
rect 208360 38880 208520 39040
rect 208360 39040 208520 39200
rect 208360 39200 208520 39360
rect 208360 39360 208520 39520
rect 208360 39520 208520 39680
rect 208360 39680 208520 39840
rect 208360 39840 208520 40000
rect 208360 40000 208520 40160
rect 208360 40160 208520 40320
rect 208360 40320 208520 40480
rect 208360 40480 208520 40640
rect 208360 40640 208520 40800
rect 208360 40800 208520 40960
rect 208360 40960 208520 41120
rect 208360 41120 208520 41280
rect 208360 41280 208520 41440
rect 208360 41440 208520 41600
rect 208360 41600 208520 41760
rect 208360 41760 208520 41920
rect 208360 41920 208520 42080
rect 208360 42080 208520 42240
rect 208360 42240 208520 42400
rect 208360 42400 208520 42560
rect 208360 42560 208520 42720
rect 208360 42720 208520 42880
rect 208360 42880 208520 43040
rect 208360 43040 208520 43200
rect 208360 43200 208520 43360
rect 208360 43360 208520 43520
rect 208360 43520 208520 43680
rect 208360 43680 208520 43840
rect 208360 43840 208520 44000
rect 208360 44000 208520 44160
rect 208360 44160 208520 44320
rect 208360 44320 208520 44480
rect 208360 44480 208520 44640
rect 208360 44640 208520 44800
rect 208360 44800 208520 44960
rect 208360 44960 208520 45120
rect 208360 45120 208520 45280
rect 208360 45280 208520 45440
rect 208360 47040 208520 47200
rect 208360 47200 208520 47360
rect 208360 47360 208520 47520
rect 208360 47520 208520 47680
rect 208360 47680 208520 47840
rect 208360 47840 208520 48000
rect 208360 48000 208520 48160
rect 208360 48160 208520 48320
rect 208360 48320 208520 48480
rect 208360 48480 208520 48640
rect 208360 48640 208520 48800
rect 208360 48800 208520 48960
rect 208360 48960 208520 49120
rect 208360 49120 208520 49280
rect 208360 49280 208520 49440
rect 208360 49440 208520 49600
rect 208360 49600 208520 49760
rect 208360 49760 208520 49920
rect 208360 49920 208520 50080
rect 208360 50080 208520 50240
rect 208360 50240 208520 50400
rect 208360 50880 208520 51040
rect 208360 51040 208520 51200
rect 208360 51200 208520 51360
rect 208360 51360 208520 51520
rect 208360 51520 208520 51680
rect 208360 51680 208520 51840
rect 208360 51840 208520 52000
rect 208360 52000 208520 52160
rect 208360 52160 208520 52320
rect 208360 52320 208520 52480
rect 208360 52480 208520 52640
rect 208360 52640 208520 52800
rect 208360 52800 208520 52960
rect 208360 52960 208520 53120
rect 208360 53120 208520 53280
rect 208360 53280 208520 53440
rect 208360 53440 208520 53600
rect 208360 53600 208520 53760
rect 208360 53760 208520 53920
rect 208360 53920 208520 54080
rect 208360 54080 208520 54240
rect 208360 54240 208520 54400
rect 208520 26400 208680 26560
rect 208520 26560 208680 26720
rect 208520 26720 208680 26880
rect 208520 26880 208680 27040
rect 208520 27040 208680 27200
rect 208520 27200 208680 27360
rect 208520 27360 208680 27520
rect 208520 27520 208680 27680
rect 208520 27680 208680 27840
rect 208520 27840 208680 28000
rect 208520 28000 208680 28160
rect 208520 28160 208680 28320
rect 208520 28320 208680 28480
rect 208520 28480 208680 28640
rect 208520 28640 208680 28800
rect 208520 28800 208680 28960
rect 208520 28960 208680 29120
rect 208520 29120 208680 29280
rect 208520 29280 208680 29440
rect 208520 29440 208680 29600
rect 208520 29600 208680 29760
rect 208520 29760 208680 29920
rect 208520 29920 208680 30080
rect 208520 30080 208680 30240
rect 208520 30240 208680 30400
rect 208520 30400 208680 30560
rect 208520 30560 208680 30720
rect 208520 30720 208680 30880
rect 208520 30880 208680 31040
rect 208520 31040 208680 31200
rect 208520 31200 208680 31360
rect 208520 31360 208680 31520
rect 208520 31520 208680 31680
rect 208520 31680 208680 31840
rect 208520 31840 208680 32000
rect 208520 32000 208680 32160
rect 208520 32160 208680 32320
rect 208520 32320 208680 32480
rect 208520 32480 208680 32640
rect 208520 32640 208680 32800
rect 208520 32800 208680 32960
rect 208520 32960 208680 33120
rect 208520 33120 208680 33280
rect 208520 33280 208680 33440
rect 208520 33440 208680 33600
rect 208520 33600 208680 33760
rect 208520 33760 208680 33920
rect 208520 33920 208680 34080
rect 208520 34080 208680 34240
rect 208520 34240 208680 34400
rect 208520 34400 208680 34560
rect 208520 34560 208680 34720
rect 208520 34720 208680 34880
rect 208520 34880 208680 35040
rect 208520 35040 208680 35200
rect 208520 35200 208680 35360
rect 208520 35360 208680 35520
rect 208520 35520 208680 35680
rect 208520 35680 208680 35840
rect 208520 35840 208680 36000
rect 208520 36000 208680 36160
rect 208520 36160 208680 36320
rect 208520 36320 208680 36480
rect 208520 36480 208680 36640
rect 208520 36640 208680 36800
rect 208520 36800 208680 36960
rect 208520 36960 208680 37120
rect 208520 37120 208680 37280
rect 208520 37280 208680 37440
rect 208520 37440 208680 37600
rect 208520 37600 208680 37760
rect 208520 37760 208680 37920
rect 208520 37920 208680 38080
rect 208520 38080 208680 38240
rect 208520 38240 208680 38400
rect 208520 38400 208680 38560
rect 208520 38560 208680 38720
rect 208520 38720 208680 38880
rect 208520 38880 208680 39040
rect 208520 39040 208680 39200
rect 208520 39200 208680 39360
rect 208520 39360 208680 39520
rect 208520 39520 208680 39680
rect 208520 39680 208680 39840
rect 208520 39840 208680 40000
rect 208520 40000 208680 40160
rect 208520 40160 208680 40320
rect 208520 40320 208680 40480
rect 208520 40480 208680 40640
rect 208520 40640 208680 40800
rect 208520 40800 208680 40960
rect 208520 40960 208680 41120
rect 208520 41120 208680 41280
rect 208520 41280 208680 41440
rect 208520 41440 208680 41600
rect 208520 41600 208680 41760
rect 208520 41760 208680 41920
rect 208520 41920 208680 42080
rect 208520 42080 208680 42240
rect 208520 42240 208680 42400
rect 208520 42400 208680 42560
rect 208520 42560 208680 42720
rect 208520 42720 208680 42880
rect 208520 42880 208680 43040
rect 208520 43040 208680 43200
rect 208520 43200 208680 43360
rect 208520 43360 208680 43520
rect 208520 43520 208680 43680
rect 208520 43680 208680 43840
rect 208520 43840 208680 44000
rect 208520 44000 208680 44160
rect 208520 44160 208680 44320
rect 208520 44320 208680 44480
rect 208520 44480 208680 44640
rect 208520 44640 208680 44800
rect 208520 44800 208680 44960
rect 208520 44960 208680 45120
rect 208520 45120 208680 45280
rect 208520 45280 208680 45440
rect 208520 45440 208680 45600
rect 208520 47040 208680 47200
rect 208520 47200 208680 47360
rect 208520 47360 208680 47520
rect 208520 47520 208680 47680
rect 208520 47680 208680 47840
rect 208520 47840 208680 48000
rect 208520 48000 208680 48160
rect 208520 48160 208680 48320
rect 208520 48320 208680 48480
rect 208520 48480 208680 48640
rect 208520 48640 208680 48800
rect 208520 48800 208680 48960
rect 208520 48960 208680 49120
rect 208520 49120 208680 49280
rect 208520 49280 208680 49440
rect 208520 49440 208680 49600
rect 208520 49600 208680 49760
rect 208520 49760 208680 49920
rect 208520 51360 208680 51520
rect 208520 51520 208680 51680
rect 208520 51680 208680 51840
rect 208520 51840 208680 52000
rect 208520 52000 208680 52160
rect 208520 52160 208680 52320
rect 208520 52320 208680 52480
rect 208520 52480 208680 52640
rect 208520 52640 208680 52800
rect 208520 52800 208680 52960
rect 208520 52960 208680 53120
rect 208520 53120 208680 53280
rect 208520 53280 208680 53440
rect 208520 53440 208680 53600
rect 208520 53600 208680 53760
rect 208520 53760 208680 53920
rect 208520 53920 208680 54080
rect 208520 54080 208680 54240
rect 208520 54240 208680 54400
rect 208520 54400 208680 54560
rect 208680 26560 208840 26720
rect 208680 26720 208840 26880
rect 208680 26880 208840 27040
rect 208680 27040 208840 27200
rect 208680 27200 208840 27360
rect 208680 27360 208840 27520
rect 208680 27520 208840 27680
rect 208680 27680 208840 27840
rect 208680 27840 208840 28000
rect 208680 28000 208840 28160
rect 208680 28160 208840 28320
rect 208680 28320 208840 28480
rect 208680 28480 208840 28640
rect 208680 28640 208840 28800
rect 208680 28800 208840 28960
rect 208680 28960 208840 29120
rect 208680 29120 208840 29280
rect 208680 29280 208840 29440
rect 208680 29440 208840 29600
rect 208680 29600 208840 29760
rect 208680 29760 208840 29920
rect 208680 29920 208840 30080
rect 208680 30080 208840 30240
rect 208680 30240 208840 30400
rect 208680 30400 208840 30560
rect 208680 30560 208840 30720
rect 208680 30720 208840 30880
rect 208680 30880 208840 31040
rect 208680 31040 208840 31200
rect 208680 31200 208840 31360
rect 208680 31360 208840 31520
rect 208680 31520 208840 31680
rect 208680 31680 208840 31840
rect 208680 31840 208840 32000
rect 208680 32000 208840 32160
rect 208680 32160 208840 32320
rect 208680 32320 208840 32480
rect 208680 32480 208840 32640
rect 208680 32640 208840 32800
rect 208680 32800 208840 32960
rect 208680 32960 208840 33120
rect 208680 33120 208840 33280
rect 208680 33280 208840 33440
rect 208680 33440 208840 33600
rect 208680 33600 208840 33760
rect 208680 33760 208840 33920
rect 208680 33920 208840 34080
rect 208680 34080 208840 34240
rect 208680 34240 208840 34400
rect 208680 34400 208840 34560
rect 208680 34560 208840 34720
rect 208680 34720 208840 34880
rect 208680 34880 208840 35040
rect 208680 35040 208840 35200
rect 208680 35200 208840 35360
rect 208680 35360 208840 35520
rect 208680 35520 208840 35680
rect 208680 35680 208840 35840
rect 208680 35840 208840 36000
rect 208680 36000 208840 36160
rect 208680 36160 208840 36320
rect 208680 36320 208840 36480
rect 208680 36480 208840 36640
rect 208680 36640 208840 36800
rect 208680 36800 208840 36960
rect 208680 36960 208840 37120
rect 208680 37120 208840 37280
rect 208680 37280 208840 37440
rect 208680 37440 208840 37600
rect 208680 37600 208840 37760
rect 208680 37760 208840 37920
rect 208680 37920 208840 38080
rect 208680 38080 208840 38240
rect 208680 38240 208840 38400
rect 208680 38400 208840 38560
rect 208680 38560 208840 38720
rect 208680 38720 208840 38880
rect 208680 38880 208840 39040
rect 208680 39040 208840 39200
rect 208680 39200 208840 39360
rect 208680 39360 208840 39520
rect 208680 39520 208840 39680
rect 208680 39680 208840 39840
rect 208680 39840 208840 40000
rect 208680 40000 208840 40160
rect 208680 40160 208840 40320
rect 208680 40320 208840 40480
rect 208680 40480 208840 40640
rect 208680 40640 208840 40800
rect 208680 40800 208840 40960
rect 208680 40960 208840 41120
rect 208680 41120 208840 41280
rect 208680 41280 208840 41440
rect 208680 41440 208840 41600
rect 208680 41600 208840 41760
rect 208680 41760 208840 41920
rect 208680 41920 208840 42080
rect 208680 42080 208840 42240
rect 208680 42240 208840 42400
rect 208680 42400 208840 42560
rect 208680 42560 208840 42720
rect 208680 42720 208840 42880
rect 208680 42880 208840 43040
rect 208680 43040 208840 43200
rect 208680 43200 208840 43360
rect 208680 43360 208840 43520
rect 208680 43520 208840 43680
rect 208680 43680 208840 43840
rect 208680 43840 208840 44000
rect 208680 44000 208840 44160
rect 208680 44160 208840 44320
rect 208680 44320 208840 44480
rect 208680 44480 208840 44640
rect 208680 44640 208840 44800
rect 208680 44800 208840 44960
rect 208680 44960 208840 45120
rect 208680 45120 208840 45280
rect 208680 45280 208840 45440
rect 208680 45440 208840 45600
rect 208680 47040 208840 47200
rect 208680 47200 208840 47360
rect 208680 47360 208840 47520
rect 208680 47520 208840 47680
rect 208680 47680 208840 47840
rect 208680 47840 208840 48000
rect 208680 48000 208840 48160
rect 208680 48160 208840 48320
rect 208680 48320 208840 48480
rect 208680 48480 208840 48640
rect 208680 48640 208840 48800
rect 208680 48800 208840 48960
rect 208680 48960 208840 49120
rect 208680 49120 208840 49280
rect 208680 49280 208840 49440
rect 208680 49440 208840 49600
rect 208680 49600 208840 49760
rect 208680 51520 208840 51680
rect 208680 51680 208840 51840
rect 208680 51840 208840 52000
rect 208680 52000 208840 52160
rect 208680 52160 208840 52320
rect 208680 52320 208840 52480
rect 208680 52480 208840 52640
rect 208680 52640 208840 52800
rect 208680 52800 208840 52960
rect 208680 52960 208840 53120
rect 208680 53120 208840 53280
rect 208680 53280 208840 53440
rect 208680 53440 208840 53600
rect 208680 53600 208840 53760
rect 208680 53760 208840 53920
rect 208680 53920 208840 54080
rect 208680 54080 208840 54240
rect 208680 54240 208840 54400
rect 208680 54400 208840 54560
rect 208840 26720 209000 26880
rect 208840 26880 209000 27040
rect 208840 27040 209000 27200
rect 208840 27200 209000 27360
rect 208840 27360 209000 27520
rect 208840 27520 209000 27680
rect 208840 27680 209000 27840
rect 208840 27840 209000 28000
rect 208840 28000 209000 28160
rect 208840 28160 209000 28320
rect 208840 28320 209000 28480
rect 208840 28480 209000 28640
rect 208840 28640 209000 28800
rect 208840 28800 209000 28960
rect 208840 28960 209000 29120
rect 208840 29120 209000 29280
rect 208840 29280 209000 29440
rect 208840 29440 209000 29600
rect 208840 29600 209000 29760
rect 208840 29760 209000 29920
rect 208840 29920 209000 30080
rect 208840 30080 209000 30240
rect 208840 30240 209000 30400
rect 208840 30400 209000 30560
rect 208840 30560 209000 30720
rect 208840 30720 209000 30880
rect 208840 30880 209000 31040
rect 208840 31040 209000 31200
rect 208840 31200 209000 31360
rect 208840 31360 209000 31520
rect 208840 31520 209000 31680
rect 208840 31680 209000 31840
rect 208840 31840 209000 32000
rect 208840 32000 209000 32160
rect 208840 32160 209000 32320
rect 208840 32320 209000 32480
rect 208840 32480 209000 32640
rect 208840 32640 209000 32800
rect 208840 32800 209000 32960
rect 208840 32960 209000 33120
rect 208840 33120 209000 33280
rect 208840 33280 209000 33440
rect 208840 33440 209000 33600
rect 208840 33600 209000 33760
rect 208840 33760 209000 33920
rect 208840 33920 209000 34080
rect 208840 34080 209000 34240
rect 208840 34240 209000 34400
rect 208840 34400 209000 34560
rect 208840 34560 209000 34720
rect 208840 34720 209000 34880
rect 208840 34880 209000 35040
rect 208840 35040 209000 35200
rect 208840 35200 209000 35360
rect 208840 35360 209000 35520
rect 208840 35520 209000 35680
rect 208840 35680 209000 35840
rect 208840 35840 209000 36000
rect 208840 36000 209000 36160
rect 208840 36160 209000 36320
rect 208840 36320 209000 36480
rect 208840 36480 209000 36640
rect 208840 36640 209000 36800
rect 208840 36800 209000 36960
rect 208840 36960 209000 37120
rect 208840 37120 209000 37280
rect 208840 37280 209000 37440
rect 208840 37440 209000 37600
rect 208840 37600 209000 37760
rect 208840 37760 209000 37920
rect 208840 37920 209000 38080
rect 208840 38080 209000 38240
rect 208840 38240 209000 38400
rect 208840 38400 209000 38560
rect 208840 38560 209000 38720
rect 208840 38720 209000 38880
rect 208840 38880 209000 39040
rect 208840 39040 209000 39200
rect 208840 39200 209000 39360
rect 208840 39360 209000 39520
rect 208840 39520 209000 39680
rect 208840 39680 209000 39840
rect 208840 39840 209000 40000
rect 208840 40000 209000 40160
rect 208840 40160 209000 40320
rect 208840 40320 209000 40480
rect 208840 40480 209000 40640
rect 208840 40640 209000 40800
rect 208840 40800 209000 40960
rect 208840 40960 209000 41120
rect 208840 41120 209000 41280
rect 208840 41280 209000 41440
rect 208840 41440 209000 41600
rect 208840 41600 209000 41760
rect 208840 41760 209000 41920
rect 208840 41920 209000 42080
rect 208840 42080 209000 42240
rect 208840 42240 209000 42400
rect 208840 42400 209000 42560
rect 208840 42560 209000 42720
rect 208840 42720 209000 42880
rect 208840 42880 209000 43040
rect 208840 43040 209000 43200
rect 208840 43200 209000 43360
rect 208840 43360 209000 43520
rect 208840 43520 209000 43680
rect 208840 43680 209000 43840
rect 208840 43840 209000 44000
rect 208840 44000 209000 44160
rect 208840 44160 209000 44320
rect 208840 44320 209000 44480
rect 208840 44480 209000 44640
rect 208840 44640 209000 44800
rect 208840 44800 209000 44960
rect 208840 44960 209000 45120
rect 208840 45120 209000 45280
rect 208840 45280 209000 45440
rect 208840 45440 209000 45600
rect 208840 45600 209000 45760
rect 208840 46880 209000 47040
rect 208840 47040 209000 47200
rect 208840 47200 209000 47360
rect 208840 47360 209000 47520
rect 208840 47520 209000 47680
rect 208840 47680 209000 47840
rect 208840 47840 209000 48000
rect 208840 48000 209000 48160
rect 208840 48160 209000 48320
rect 208840 48320 209000 48480
rect 208840 48480 209000 48640
rect 208840 48640 209000 48800
rect 208840 48800 209000 48960
rect 208840 48960 209000 49120
rect 208840 49120 209000 49280
rect 208840 49280 209000 49440
rect 208840 49440 209000 49600
rect 208840 51680 209000 51840
rect 208840 51840 209000 52000
rect 208840 52000 209000 52160
rect 208840 52160 209000 52320
rect 208840 52320 209000 52480
rect 208840 52480 209000 52640
rect 208840 52640 209000 52800
rect 208840 52800 209000 52960
rect 208840 52960 209000 53120
rect 208840 53120 209000 53280
rect 208840 53280 209000 53440
rect 208840 53440 209000 53600
rect 208840 53600 209000 53760
rect 208840 53760 209000 53920
rect 208840 53920 209000 54080
rect 208840 54080 209000 54240
rect 208840 54240 209000 54400
rect 208840 54400 209000 54560
rect 209000 26880 209160 27040
rect 209000 27040 209160 27200
rect 209000 27200 209160 27360
rect 209000 27360 209160 27520
rect 209000 27520 209160 27680
rect 209000 27680 209160 27840
rect 209000 27840 209160 28000
rect 209000 28000 209160 28160
rect 209000 28160 209160 28320
rect 209000 28320 209160 28480
rect 209000 28480 209160 28640
rect 209000 28640 209160 28800
rect 209000 28800 209160 28960
rect 209000 28960 209160 29120
rect 209000 29120 209160 29280
rect 209000 29280 209160 29440
rect 209000 29440 209160 29600
rect 209000 29600 209160 29760
rect 209000 29760 209160 29920
rect 209000 29920 209160 30080
rect 209000 30080 209160 30240
rect 209000 30240 209160 30400
rect 209000 30400 209160 30560
rect 209000 30560 209160 30720
rect 209000 30720 209160 30880
rect 209000 30880 209160 31040
rect 209000 31040 209160 31200
rect 209000 31200 209160 31360
rect 209000 31360 209160 31520
rect 209000 31520 209160 31680
rect 209000 31680 209160 31840
rect 209000 31840 209160 32000
rect 209000 32000 209160 32160
rect 209000 32160 209160 32320
rect 209000 32320 209160 32480
rect 209000 32480 209160 32640
rect 209000 32640 209160 32800
rect 209000 32800 209160 32960
rect 209000 32960 209160 33120
rect 209000 33120 209160 33280
rect 209000 33280 209160 33440
rect 209000 33440 209160 33600
rect 209000 33600 209160 33760
rect 209000 33760 209160 33920
rect 209000 33920 209160 34080
rect 209000 34080 209160 34240
rect 209000 34240 209160 34400
rect 209000 34400 209160 34560
rect 209000 34560 209160 34720
rect 209000 34720 209160 34880
rect 209000 34880 209160 35040
rect 209000 35040 209160 35200
rect 209000 35200 209160 35360
rect 209000 35360 209160 35520
rect 209000 35520 209160 35680
rect 209000 35680 209160 35840
rect 209000 35840 209160 36000
rect 209000 36000 209160 36160
rect 209000 36160 209160 36320
rect 209000 36320 209160 36480
rect 209000 36480 209160 36640
rect 209000 36640 209160 36800
rect 209000 36800 209160 36960
rect 209000 36960 209160 37120
rect 209000 37120 209160 37280
rect 209000 37280 209160 37440
rect 209000 37440 209160 37600
rect 209000 37600 209160 37760
rect 209000 37760 209160 37920
rect 209000 37920 209160 38080
rect 209000 38080 209160 38240
rect 209000 38240 209160 38400
rect 209000 38400 209160 38560
rect 209000 38560 209160 38720
rect 209000 38720 209160 38880
rect 209000 38880 209160 39040
rect 209000 39040 209160 39200
rect 209000 39200 209160 39360
rect 209000 39360 209160 39520
rect 209000 39520 209160 39680
rect 209000 39680 209160 39840
rect 209000 39840 209160 40000
rect 209000 40000 209160 40160
rect 209000 40160 209160 40320
rect 209000 40320 209160 40480
rect 209000 40480 209160 40640
rect 209000 40640 209160 40800
rect 209000 40800 209160 40960
rect 209000 40960 209160 41120
rect 209000 41120 209160 41280
rect 209000 41280 209160 41440
rect 209000 41440 209160 41600
rect 209000 41600 209160 41760
rect 209000 41760 209160 41920
rect 209000 41920 209160 42080
rect 209000 42080 209160 42240
rect 209000 42240 209160 42400
rect 209000 42400 209160 42560
rect 209000 42560 209160 42720
rect 209000 42720 209160 42880
rect 209000 42880 209160 43040
rect 209000 43040 209160 43200
rect 209000 43200 209160 43360
rect 209000 43360 209160 43520
rect 209000 43520 209160 43680
rect 209000 43680 209160 43840
rect 209000 43840 209160 44000
rect 209000 44000 209160 44160
rect 209000 44160 209160 44320
rect 209000 44320 209160 44480
rect 209000 44480 209160 44640
rect 209000 44640 209160 44800
rect 209000 44800 209160 44960
rect 209000 44960 209160 45120
rect 209000 45120 209160 45280
rect 209000 45280 209160 45440
rect 209000 45440 209160 45600
rect 209000 45600 209160 45760
rect 209000 46880 209160 47040
rect 209000 47040 209160 47200
rect 209000 47200 209160 47360
rect 209000 47360 209160 47520
rect 209000 47520 209160 47680
rect 209000 47680 209160 47840
rect 209000 47840 209160 48000
rect 209000 48000 209160 48160
rect 209000 48160 209160 48320
rect 209000 48320 209160 48480
rect 209000 48480 209160 48640
rect 209000 48640 209160 48800
rect 209000 48800 209160 48960
rect 209000 48960 209160 49120
rect 209000 49120 209160 49280
rect 209000 49280 209160 49440
rect 209000 51840 209160 52000
rect 209000 52000 209160 52160
rect 209000 52160 209160 52320
rect 209000 52320 209160 52480
rect 209000 52480 209160 52640
rect 209000 52640 209160 52800
rect 209000 52800 209160 52960
rect 209000 52960 209160 53120
rect 209000 53120 209160 53280
rect 209000 53280 209160 53440
rect 209000 53440 209160 53600
rect 209000 53600 209160 53760
rect 209000 53760 209160 53920
rect 209000 53920 209160 54080
rect 209000 54080 209160 54240
rect 209000 54240 209160 54400
rect 209000 54400 209160 54560
rect 209160 27200 209320 27360
rect 209160 27360 209320 27520
rect 209160 27520 209320 27680
rect 209160 27680 209320 27840
rect 209160 27840 209320 28000
rect 209160 28000 209320 28160
rect 209160 28160 209320 28320
rect 209160 28320 209320 28480
rect 209160 28480 209320 28640
rect 209160 28640 209320 28800
rect 209160 28800 209320 28960
rect 209160 28960 209320 29120
rect 209160 29120 209320 29280
rect 209160 29280 209320 29440
rect 209160 29600 209320 29760
rect 209160 36800 209320 36960
rect 209160 37120 209320 37280
rect 209160 37280 209320 37440
rect 209160 37440 209320 37600
rect 209160 37600 209320 37760
rect 209160 37760 209320 37920
rect 209160 37920 209320 38080
rect 209160 38080 209320 38240
rect 209160 38240 209320 38400
rect 209160 38400 209320 38560
rect 209160 38560 209320 38720
rect 209160 38720 209320 38880
rect 209160 38880 209320 39040
rect 209160 39040 209320 39200
rect 209160 39200 209320 39360
rect 209160 39360 209320 39520
rect 209160 39520 209320 39680
rect 209160 39680 209320 39840
rect 209160 39840 209320 40000
rect 209160 40000 209320 40160
rect 209160 40160 209320 40320
rect 209160 40320 209320 40480
rect 209160 40480 209320 40640
rect 209160 40640 209320 40800
rect 209160 40800 209320 40960
rect 209160 40960 209320 41120
rect 209160 41120 209320 41280
rect 209160 41280 209320 41440
rect 209160 41440 209320 41600
rect 209160 41600 209320 41760
rect 209160 41760 209320 41920
rect 209160 41920 209320 42080
rect 209160 42080 209320 42240
rect 209160 42240 209320 42400
rect 209160 42400 209320 42560
rect 209160 42560 209320 42720
rect 209160 42720 209320 42880
rect 209160 42880 209320 43040
rect 209160 43040 209320 43200
rect 209160 43200 209320 43360
rect 209160 43360 209320 43520
rect 209160 43520 209320 43680
rect 209160 43680 209320 43840
rect 209160 43840 209320 44000
rect 209160 44000 209320 44160
rect 209160 44160 209320 44320
rect 209160 44320 209320 44480
rect 209160 44480 209320 44640
rect 209160 44640 209320 44800
rect 209160 44800 209320 44960
rect 209160 44960 209320 45120
rect 209160 45120 209320 45280
rect 209160 45280 209320 45440
rect 209160 45440 209320 45600
rect 209160 45600 209320 45760
rect 209160 45760 209320 45920
rect 209160 46880 209320 47040
rect 209160 47040 209320 47200
rect 209160 47200 209320 47360
rect 209160 47360 209320 47520
rect 209160 47520 209320 47680
rect 209160 47680 209320 47840
rect 209160 47840 209320 48000
rect 209160 48000 209320 48160
rect 209160 48160 209320 48320
rect 209160 48320 209320 48480
rect 209160 48480 209320 48640
rect 209160 48640 209320 48800
rect 209160 48800 209320 48960
rect 209160 48960 209320 49120
rect 209160 49120 209320 49280
rect 209160 49280 209320 49440
rect 209160 51840 209320 52000
rect 209160 52000 209320 52160
rect 209160 52160 209320 52320
rect 209160 52320 209320 52480
rect 209160 52480 209320 52640
rect 209160 52640 209320 52800
rect 209160 52800 209320 52960
rect 209160 52960 209320 53120
rect 209160 53120 209320 53280
rect 209160 53280 209320 53440
rect 209160 53440 209320 53600
rect 209160 53600 209320 53760
rect 209160 53760 209320 53920
rect 209160 53920 209320 54080
rect 209160 54080 209320 54240
rect 209160 54240 209320 54400
rect 209160 54400 209320 54560
rect 209320 40160 209480 40320
rect 209320 40320 209480 40480
rect 209320 40480 209480 40640
rect 209320 40640 209480 40800
rect 209320 40800 209480 40960
rect 209320 40960 209480 41120
rect 209320 41120 209480 41280
rect 209320 41280 209480 41440
rect 209320 41440 209480 41600
rect 209320 41600 209480 41760
rect 209320 41760 209480 41920
rect 209320 41920 209480 42080
rect 209320 42080 209480 42240
rect 209320 42240 209480 42400
rect 209320 42400 209480 42560
rect 209320 42560 209480 42720
rect 209320 42720 209480 42880
rect 209320 42880 209480 43040
rect 209320 43040 209480 43200
rect 209320 43200 209480 43360
rect 209320 43360 209480 43520
rect 209320 43520 209480 43680
rect 209320 43680 209480 43840
rect 209320 43840 209480 44000
rect 209320 44000 209480 44160
rect 209320 44160 209480 44320
rect 209320 44320 209480 44480
rect 209320 44480 209480 44640
rect 209320 44640 209480 44800
rect 209320 44800 209480 44960
rect 209320 44960 209480 45120
rect 209320 45120 209480 45280
rect 209320 45280 209480 45440
rect 209320 45440 209480 45600
rect 209320 45600 209480 45760
rect 209320 45760 209480 45920
rect 209320 46880 209480 47040
rect 209320 47040 209480 47200
rect 209320 47200 209480 47360
rect 209320 47360 209480 47520
rect 209320 47520 209480 47680
rect 209320 47680 209480 47840
rect 209320 47840 209480 48000
rect 209320 48000 209480 48160
rect 209320 48160 209480 48320
rect 209320 48320 209480 48480
rect 209320 48480 209480 48640
rect 209320 48640 209480 48800
rect 209320 48800 209480 48960
rect 209320 48960 209480 49120
rect 209320 49120 209480 49280
rect 209320 49280 209480 49440
rect 209320 52000 209480 52160
rect 209320 52160 209480 52320
rect 209320 52320 209480 52480
rect 209320 52480 209480 52640
rect 209320 52640 209480 52800
rect 209320 52800 209480 52960
rect 209320 52960 209480 53120
rect 209320 53120 209480 53280
rect 209320 53280 209480 53440
rect 209320 53440 209480 53600
rect 209320 53600 209480 53760
rect 209320 53760 209480 53920
rect 209320 53920 209480 54080
rect 209320 54080 209480 54240
rect 209320 54240 209480 54400
rect 209320 54400 209480 54560
rect 209480 42560 209640 42720
rect 209480 42720 209640 42880
rect 209480 42880 209640 43040
rect 209480 43040 209640 43200
rect 209480 43200 209640 43360
rect 209480 43360 209640 43520
rect 209480 43520 209640 43680
rect 209480 43680 209640 43840
rect 209480 43840 209640 44000
rect 209480 44000 209640 44160
rect 209480 44160 209640 44320
rect 209480 44320 209640 44480
rect 209480 44480 209640 44640
rect 209480 44640 209640 44800
rect 209480 44800 209640 44960
rect 209480 44960 209640 45120
rect 209480 45120 209640 45280
rect 209480 45280 209640 45440
rect 209480 45440 209640 45600
rect 209480 45600 209640 45760
rect 209480 45760 209640 45920
rect 209480 46720 209640 46880
rect 209480 46880 209640 47040
rect 209480 47040 209640 47200
rect 209480 47200 209640 47360
rect 209480 47360 209640 47520
rect 209480 47520 209640 47680
rect 209480 47680 209640 47840
rect 209480 47840 209640 48000
rect 209480 48000 209640 48160
rect 209480 48160 209640 48320
rect 209480 48320 209640 48480
rect 209480 48480 209640 48640
rect 209480 48640 209640 48800
rect 209480 48800 209640 48960
rect 209480 48960 209640 49120
rect 209480 49120 209640 49280
rect 209480 49280 209640 49440
rect 209480 52000 209640 52160
rect 209480 52160 209640 52320
rect 209480 52320 209640 52480
rect 209480 52480 209640 52640
rect 209480 52640 209640 52800
rect 209480 52800 209640 52960
rect 209480 52960 209640 53120
rect 209480 53120 209640 53280
rect 209480 53280 209640 53440
rect 209480 53440 209640 53600
rect 209480 53600 209640 53760
rect 209480 53760 209640 53920
rect 209480 53920 209640 54080
rect 209480 54080 209640 54240
rect 209480 54240 209640 54400
rect 209480 54400 209640 54560
rect 209640 43200 209800 43360
rect 209640 43360 209800 43520
rect 209640 43520 209800 43680
rect 209640 43680 209800 43840
rect 209640 43840 209800 44000
rect 209640 44000 209800 44160
rect 209640 44160 209800 44320
rect 209640 44320 209800 44480
rect 209640 44480 209800 44640
rect 209640 44640 209800 44800
rect 209640 44800 209800 44960
rect 209640 44960 209800 45120
rect 209640 45120 209800 45280
rect 209640 45280 209800 45440
rect 209640 45440 209800 45600
rect 209640 45600 209800 45760
rect 209640 45760 209800 45920
rect 209640 46880 209800 47040
rect 209640 47040 209800 47200
rect 209640 47200 209800 47360
rect 209640 47360 209800 47520
rect 209640 47520 209800 47680
rect 209640 47680 209800 47840
rect 209640 47840 209800 48000
rect 209640 48000 209800 48160
rect 209640 48160 209800 48320
rect 209640 48320 209800 48480
rect 209640 48480 209800 48640
rect 209640 48640 209800 48800
rect 209640 48800 209800 48960
rect 209640 48960 209800 49120
rect 209640 49120 209800 49280
rect 209640 49280 209800 49440
rect 209640 52000 209800 52160
rect 209640 52160 209800 52320
rect 209640 52320 209800 52480
rect 209640 52480 209800 52640
rect 209640 52640 209800 52800
rect 209640 52800 209800 52960
rect 209640 52960 209800 53120
rect 209640 53120 209800 53280
rect 209640 53280 209800 53440
rect 209640 53440 209800 53600
rect 209640 53600 209800 53760
rect 209640 53760 209800 53920
rect 209640 53920 209800 54080
rect 209640 54080 209800 54240
rect 209640 54240 209800 54400
rect 209640 54400 209800 54560
rect 209800 43520 209960 43680
rect 209800 43680 209960 43840
rect 209800 43840 209960 44000
rect 209800 44000 209960 44160
rect 209800 44160 209960 44320
rect 209800 44320 209960 44480
rect 209800 44480 209960 44640
rect 209800 44640 209960 44800
rect 209800 44800 209960 44960
rect 209800 44960 209960 45120
rect 209800 45120 209960 45280
rect 209800 45280 209960 45440
rect 209800 45440 209960 45600
rect 209800 45600 209960 45760
rect 209800 45760 209960 45920
rect 209800 46720 209960 46880
rect 209800 46880 209960 47040
rect 209800 47040 209960 47200
rect 209800 47200 209960 47360
rect 209800 47360 209960 47520
rect 209800 47520 209960 47680
rect 209800 47680 209960 47840
rect 209800 47840 209960 48000
rect 209800 48000 209960 48160
rect 209800 48160 209960 48320
rect 209800 48320 209960 48480
rect 209800 48480 209960 48640
rect 209800 48640 209960 48800
rect 209800 48800 209960 48960
rect 209800 48960 209960 49120
rect 209800 49120 209960 49280
rect 209800 49280 209960 49440
rect 209800 52000 209960 52160
rect 209800 52160 209960 52320
rect 209800 52320 209960 52480
rect 209800 52480 209960 52640
rect 209800 52640 209960 52800
rect 209800 52800 209960 52960
rect 209800 52960 209960 53120
rect 209800 53120 209960 53280
rect 209800 53280 209960 53440
rect 209800 53440 209960 53600
rect 209800 53600 209960 53760
rect 209800 53760 209960 53920
rect 209800 53920 209960 54080
rect 209800 54080 209960 54240
rect 209800 54240 209960 54400
rect 209800 54400 209960 54560
rect 209960 43840 210120 44000
rect 209960 44000 210120 44160
rect 209960 44160 210120 44320
rect 209960 44320 210120 44480
rect 209960 44480 210120 44640
rect 209960 44640 210120 44800
rect 209960 44800 210120 44960
rect 209960 44960 210120 45120
rect 209960 45120 210120 45280
rect 209960 45280 210120 45440
rect 209960 45440 210120 45600
rect 209960 45600 210120 45760
rect 209960 45760 210120 45920
rect 209960 46720 210120 46880
rect 209960 46880 210120 47040
rect 209960 47040 210120 47200
rect 209960 47200 210120 47360
rect 209960 47360 210120 47520
rect 209960 47520 210120 47680
rect 209960 47680 210120 47840
rect 209960 47840 210120 48000
rect 209960 48000 210120 48160
rect 209960 48160 210120 48320
rect 209960 48320 210120 48480
rect 209960 48480 210120 48640
rect 209960 48640 210120 48800
rect 209960 48800 210120 48960
rect 209960 48960 210120 49120
rect 209960 49120 210120 49280
rect 209960 49280 210120 49440
rect 209960 49440 210120 49600
rect 209960 52000 210120 52160
rect 209960 52160 210120 52320
rect 209960 52320 210120 52480
rect 209960 52480 210120 52640
rect 209960 52640 210120 52800
rect 209960 52800 210120 52960
rect 209960 52960 210120 53120
rect 209960 53120 210120 53280
rect 209960 53280 210120 53440
rect 209960 53440 210120 53600
rect 209960 53600 210120 53760
rect 209960 53760 210120 53920
rect 209960 53920 210120 54080
rect 209960 54080 210120 54240
rect 209960 54240 210120 54400
rect 209960 54400 210120 54560
rect 210120 44320 210280 44480
rect 210120 44480 210280 44640
rect 210120 44640 210280 44800
rect 210120 44800 210280 44960
rect 210120 44960 210280 45120
rect 210120 45120 210280 45280
rect 210120 45280 210280 45440
rect 210120 45440 210280 45600
rect 210120 45600 210280 45760
rect 210120 45760 210280 45920
rect 210120 46720 210280 46880
rect 210120 46880 210280 47040
rect 210120 47040 210280 47200
rect 210120 47200 210280 47360
rect 210120 47360 210280 47520
rect 210120 47520 210280 47680
rect 210120 47680 210280 47840
rect 210120 47840 210280 48000
rect 210120 48000 210280 48160
rect 210120 48160 210280 48320
rect 210120 48320 210280 48480
rect 210120 48480 210280 48640
rect 210120 48640 210280 48800
rect 210120 48800 210280 48960
rect 210120 48960 210280 49120
rect 210120 49120 210280 49280
rect 210120 49280 210280 49440
rect 210120 49440 210280 49600
rect 210120 52000 210280 52160
rect 210120 52160 210280 52320
rect 210120 52320 210280 52480
rect 210120 52480 210280 52640
rect 210120 52640 210280 52800
rect 210120 52800 210280 52960
rect 210120 52960 210280 53120
rect 210120 53120 210280 53280
rect 210120 53280 210280 53440
rect 210120 53440 210280 53600
rect 210120 53600 210280 53760
rect 210120 53760 210280 53920
rect 210120 53920 210280 54080
rect 210120 54080 210280 54240
rect 210120 54240 210280 54400
rect 210120 54400 210280 54560
rect 210280 44800 210440 44960
rect 210280 44960 210440 45120
rect 210280 45120 210440 45280
rect 210280 45280 210440 45440
rect 210280 45440 210440 45600
rect 210280 45600 210440 45760
rect 210280 45760 210440 45920
rect 210280 46720 210440 46880
rect 210280 46880 210440 47040
rect 210280 47040 210440 47200
rect 210280 47200 210440 47360
rect 210280 47360 210440 47520
rect 210280 47520 210440 47680
rect 210280 47680 210440 47840
rect 210280 47840 210440 48000
rect 210280 48000 210440 48160
rect 210280 48160 210440 48320
rect 210280 48320 210440 48480
rect 210280 48480 210440 48640
rect 210280 48640 210440 48800
rect 210280 48800 210440 48960
rect 210280 48960 210440 49120
rect 210280 49120 210440 49280
rect 210280 49280 210440 49440
rect 210280 49440 210440 49600
rect 210280 49600 210440 49760
rect 210280 51840 210440 52000
rect 210280 52000 210440 52160
rect 210280 52160 210440 52320
rect 210280 52320 210440 52480
rect 210280 52480 210440 52640
rect 210280 52640 210440 52800
rect 210280 52800 210440 52960
rect 210280 52960 210440 53120
rect 210280 53120 210440 53280
rect 210280 53280 210440 53440
rect 210280 53440 210440 53600
rect 210280 53600 210440 53760
rect 210280 53760 210440 53920
rect 210280 53920 210440 54080
rect 210280 54080 210440 54240
rect 210280 54240 210440 54400
rect 210440 45440 210600 45600
rect 210440 45600 210600 45760
rect 210440 45760 210600 45920
rect 210440 46880 210600 47040
rect 210440 47040 210600 47200
rect 210440 47200 210600 47360
rect 210440 47360 210600 47520
rect 210440 47520 210600 47680
rect 210440 47680 210600 47840
rect 210440 47840 210600 48000
rect 210440 48000 210600 48160
rect 210440 48160 210600 48320
rect 210440 48320 210600 48480
rect 210440 48480 210600 48640
rect 210440 48640 210600 48800
rect 210440 48800 210600 48960
rect 210440 48960 210600 49120
rect 210440 49120 210600 49280
rect 210440 49280 210600 49440
rect 210440 49440 210600 49600
rect 210440 49600 210600 49760
rect 210440 49760 210600 49920
rect 210440 51680 210600 51840
rect 210440 51840 210600 52000
rect 210440 52000 210600 52160
rect 210440 52160 210600 52320
rect 210440 52320 210600 52480
rect 210440 52480 210600 52640
rect 210440 52640 210600 52800
rect 210440 52800 210600 52960
rect 210440 52960 210600 53120
rect 210440 53120 210600 53280
rect 210440 53280 210600 53440
rect 210440 53440 210600 53600
rect 210440 53600 210600 53760
rect 210440 53760 210600 53920
rect 210440 53920 210600 54080
rect 210440 54080 210600 54240
rect 210440 54240 210600 54400
rect 210600 46880 210760 47040
rect 210600 47040 210760 47200
rect 210600 47200 210760 47360
rect 210600 47360 210760 47520
rect 210600 47520 210760 47680
rect 210600 47680 210760 47840
rect 210600 47840 210760 48000
rect 210600 48000 210760 48160
rect 210600 48160 210760 48320
rect 210600 48320 210760 48480
rect 210600 48480 210760 48640
rect 210600 48640 210760 48800
rect 210600 48800 210760 48960
rect 210600 48960 210760 49120
rect 210600 49120 210760 49280
rect 210600 49280 210760 49440
rect 210600 49440 210760 49600
rect 210600 49600 210760 49760
rect 210600 49760 210760 49920
rect 210600 49920 210760 50080
rect 210600 51520 210760 51680
rect 210600 51680 210760 51840
rect 210600 51840 210760 52000
rect 210600 52000 210760 52160
rect 210600 52160 210760 52320
rect 210600 52320 210760 52480
rect 210600 52480 210760 52640
rect 210600 52640 210760 52800
rect 210600 52800 210760 52960
rect 210600 52960 210760 53120
rect 210600 53120 210760 53280
rect 210600 53280 210760 53440
rect 210600 53440 210760 53600
rect 210600 53600 210760 53760
rect 210600 53760 210760 53920
rect 210600 53920 210760 54080
rect 210600 54080 210760 54240
rect 210600 54240 210760 54400
rect 210760 46880 210920 47040
rect 210760 47040 210920 47200
rect 210760 47200 210920 47360
rect 210760 47360 210920 47520
rect 210760 47520 210920 47680
rect 210760 47680 210920 47840
rect 210760 47840 210920 48000
rect 210760 48000 210920 48160
rect 210760 48160 210920 48320
rect 210760 48320 210920 48480
rect 210760 48480 210920 48640
rect 210760 48640 210920 48800
rect 210760 48800 210920 48960
rect 210760 48960 210920 49120
rect 210760 49120 210920 49280
rect 210760 49280 210920 49440
rect 210760 49440 210920 49600
rect 210760 49600 210920 49760
rect 210760 49760 210920 49920
rect 210760 49920 210920 50080
rect 210760 50080 210920 50240
rect 210760 50240 210920 50400
rect 210760 51360 210920 51520
rect 210760 51520 210920 51680
rect 210760 51680 210920 51840
rect 210760 51840 210920 52000
rect 210760 52000 210920 52160
rect 210760 52160 210920 52320
rect 210760 52320 210920 52480
rect 210760 52480 210920 52640
rect 210760 52640 210920 52800
rect 210760 52800 210920 52960
rect 210760 52960 210920 53120
rect 210760 53120 210920 53280
rect 210760 53280 210920 53440
rect 210760 53440 210920 53600
rect 210760 53600 210920 53760
rect 210760 53760 210920 53920
rect 210760 53920 210920 54080
rect 210760 54080 210920 54240
rect 210920 46880 211080 47040
rect 210920 47040 211080 47200
rect 210920 47200 211080 47360
rect 210920 47360 211080 47520
rect 210920 47520 211080 47680
rect 210920 47680 211080 47840
rect 210920 47840 211080 48000
rect 210920 48000 211080 48160
rect 210920 48160 211080 48320
rect 210920 48320 211080 48480
rect 210920 48480 211080 48640
rect 210920 48640 211080 48800
rect 210920 48800 211080 48960
rect 210920 48960 211080 49120
rect 210920 49120 211080 49280
rect 210920 49280 211080 49440
rect 210920 49440 211080 49600
rect 210920 49600 211080 49760
rect 210920 49760 211080 49920
rect 210920 49920 211080 50080
rect 210920 50080 211080 50240
rect 210920 50240 211080 50400
rect 210920 50400 211080 50560
rect 210920 50560 211080 50720
rect 210920 50720 211080 50880
rect 210920 50880 211080 51040
rect 210920 51040 211080 51200
rect 210920 51200 211080 51360
rect 210920 51360 211080 51520
rect 210920 51520 211080 51680
rect 210920 51680 211080 51840
rect 210920 51840 211080 52000
rect 210920 52000 211080 52160
rect 210920 52160 211080 52320
rect 210920 52320 211080 52480
rect 210920 52480 211080 52640
rect 210920 52640 211080 52800
rect 210920 52800 211080 52960
rect 210920 52960 211080 53120
rect 210920 53120 211080 53280
rect 210920 53280 211080 53440
rect 210920 53440 211080 53600
rect 210920 53600 211080 53760
rect 210920 53760 211080 53920
rect 210920 53920 211080 54080
rect 210920 54080 211080 54240
rect 211080 46880 211240 47040
rect 211080 47040 211240 47200
rect 211080 47200 211240 47360
rect 211080 47360 211240 47520
rect 211080 47520 211240 47680
rect 211080 47680 211240 47840
rect 211080 47840 211240 48000
rect 211080 48000 211240 48160
rect 211080 48160 211240 48320
rect 211080 48320 211240 48480
rect 211080 48480 211240 48640
rect 211080 48640 211240 48800
rect 211080 48800 211240 48960
rect 211080 48960 211240 49120
rect 211080 49120 211240 49280
rect 211080 49280 211240 49440
rect 211080 49440 211240 49600
rect 211080 49600 211240 49760
rect 211080 49760 211240 49920
rect 211080 49920 211240 50080
rect 211080 50080 211240 50240
rect 211080 50240 211240 50400
rect 211080 50400 211240 50560
rect 211080 50560 211240 50720
rect 211080 50720 211240 50880
rect 211080 50880 211240 51040
rect 211080 51040 211240 51200
rect 211080 51200 211240 51360
rect 211080 51360 211240 51520
rect 211080 51520 211240 51680
rect 211080 51680 211240 51840
rect 211080 51840 211240 52000
rect 211080 52000 211240 52160
rect 211080 52160 211240 52320
rect 211080 52320 211240 52480
rect 211080 52480 211240 52640
rect 211080 52640 211240 52800
rect 211080 52800 211240 52960
rect 211080 52960 211240 53120
rect 211080 53120 211240 53280
rect 211080 53280 211240 53440
rect 211080 53440 211240 53600
rect 211080 53600 211240 53760
rect 211080 53760 211240 53920
rect 211080 53920 211240 54080
rect 211240 47040 211400 47200
rect 211240 47200 211400 47360
rect 211240 47360 211400 47520
rect 211240 47520 211400 47680
rect 211240 47680 211400 47840
rect 211240 47840 211400 48000
rect 211240 48000 211400 48160
rect 211240 48160 211400 48320
rect 211240 48320 211400 48480
rect 211240 48480 211400 48640
rect 211240 48640 211400 48800
rect 211240 48800 211400 48960
rect 211240 48960 211400 49120
rect 211240 49120 211400 49280
rect 211240 49280 211400 49440
rect 211240 49440 211400 49600
rect 211240 49600 211400 49760
rect 211240 49760 211400 49920
rect 211240 49920 211400 50080
rect 211240 50080 211400 50240
rect 211240 50240 211400 50400
rect 211240 50400 211400 50560
rect 211240 50560 211400 50720
rect 211240 50720 211400 50880
rect 211240 50880 211400 51040
rect 211240 51040 211400 51200
rect 211240 51200 211400 51360
rect 211240 51360 211400 51520
rect 211240 51520 211400 51680
rect 211240 51680 211400 51840
rect 211240 51840 211400 52000
rect 211240 52000 211400 52160
rect 211240 52160 211400 52320
rect 211240 52320 211400 52480
rect 211240 52480 211400 52640
rect 211240 52640 211400 52800
rect 211240 52800 211400 52960
rect 211240 52960 211400 53120
rect 211240 53120 211400 53280
rect 211240 53280 211400 53440
rect 211240 53440 211400 53600
rect 211240 53600 211400 53760
rect 211240 53760 211400 53920
rect 211240 53920 211400 54080
rect 211400 47040 211560 47200
rect 211400 47200 211560 47360
rect 211400 47360 211560 47520
rect 211400 47520 211560 47680
rect 211400 47680 211560 47840
rect 211400 47840 211560 48000
rect 211400 48000 211560 48160
rect 211400 48160 211560 48320
rect 211400 48320 211560 48480
rect 211400 48480 211560 48640
rect 211400 48640 211560 48800
rect 211400 48800 211560 48960
rect 211400 48960 211560 49120
rect 211400 49120 211560 49280
rect 211400 49280 211560 49440
rect 211400 49440 211560 49600
rect 211400 49600 211560 49760
rect 211400 49760 211560 49920
rect 211400 49920 211560 50080
rect 211400 50080 211560 50240
rect 211400 50240 211560 50400
rect 211400 50400 211560 50560
rect 211400 50560 211560 50720
rect 211400 50720 211560 50880
rect 211400 50880 211560 51040
rect 211400 51040 211560 51200
rect 211400 51200 211560 51360
rect 211400 51360 211560 51520
rect 211400 51520 211560 51680
rect 211400 51680 211560 51840
rect 211400 51840 211560 52000
rect 211400 52000 211560 52160
rect 211400 52160 211560 52320
rect 211400 52320 211560 52480
rect 211400 52480 211560 52640
rect 211400 52640 211560 52800
rect 211400 52800 211560 52960
rect 211400 52960 211560 53120
rect 211400 53120 211560 53280
rect 211400 53280 211560 53440
rect 211400 53440 211560 53600
rect 211400 53600 211560 53760
rect 211400 53760 211560 53920
rect 211560 47200 211720 47360
rect 211560 47360 211720 47520
rect 211560 47520 211720 47680
rect 211560 47680 211720 47840
rect 211560 47840 211720 48000
rect 211560 48000 211720 48160
rect 211560 48160 211720 48320
rect 211560 48320 211720 48480
rect 211560 48480 211720 48640
rect 211560 48640 211720 48800
rect 211560 48800 211720 48960
rect 211560 48960 211720 49120
rect 211560 49120 211720 49280
rect 211560 49280 211720 49440
rect 211560 49440 211720 49600
rect 211560 49600 211720 49760
rect 211560 49760 211720 49920
rect 211560 49920 211720 50080
rect 211560 50080 211720 50240
rect 211560 50240 211720 50400
rect 211560 50400 211720 50560
rect 211560 50560 211720 50720
rect 211560 50720 211720 50880
rect 211560 50880 211720 51040
rect 211560 51040 211720 51200
rect 211560 51200 211720 51360
rect 211560 51360 211720 51520
rect 211560 51520 211720 51680
rect 211560 51680 211720 51840
rect 211560 51840 211720 52000
rect 211560 52000 211720 52160
rect 211560 52160 211720 52320
rect 211560 52320 211720 52480
rect 211560 52480 211720 52640
rect 211560 52640 211720 52800
rect 211560 52800 211720 52960
rect 211560 52960 211720 53120
rect 211560 53120 211720 53280
rect 211560 53280 211720 53440
rect 211560 53440 211720 53600
rect 211560 53600 211720 53760
rect 211720 47200 211880 47360
rect 211720 47360 211880 47520
rect 211720 47520 211880 47680
rect 211720 47680 211880 47840
rect 211720 47840 211880 48000
rect 211720 48000 211880 48160
rect 211720 48160 211880 48320
rect 211720 48320 211880 48480
rect 211720 48480 211880 48640
rect 211720 48640 211880 48800
rect 211720 48800 211880 48960
rect 211720 48960 211880 49120
rect 211720 49120 211880 49280
rect 211720 49280 211880 49440
rect 211720 49440 211880 49600
rect 211720 49600 211880 49760
rect 211720 49760 211880 49920
rect 211720 49920 211880 50080
rect 211720 50080 211880 50240
rect 211720 50240 211880 50400
rect 211720 50400 211880 50560
rect 211720 50560 211880 50720
rect 211720 50720 211880 50880
rect 211720 50880 211880 51040
rect 211720 51040 211880 51200
rect 211720 51200 211880 51360
rect 211720 51360 211880 51520
rect 211720 51520 211880 51680
rect 211720 51680 211880 51840
rect 211720 51840 211880 52000
rect 211720 52000 211880 52160
rect 211720 52160 211880 52320
rect 211720 52320 211880 52480
rect 211720 52480 211880 52640
rect 211720 52640 211880 52800
rect 211720 52800 211880 52960
rect 211720 52960 211880 53120
rect 211720 53120 211880 53280
rect 211720 53280 211880 53440
rect 211720 53440 211880 53600
rect 211880 47360 212040 47520
rect 211880 47520 212040 47680
rect 211880 47680 212040 47840
rect 211880 47840 212040 48000
rect 211880 48000 212040 48160
rect 211880 48160 212040 48320
rect 211880 48320 212040 48480
rect 211880 48480 212040 48640
rect 211880 48640 212040 48800
rect 211880 48800 212040 48960
rect 211880 48960 212040 49120
rect 211880 49120 212040 49280
rect 211880 49280 212040 49440
rect 211880 49440 212040 49600
rect 211880 49600 212040 49760
rect 211880 49760 212040 49920
rect 211880 49920 212040 50080
rect 211880 50080 212040 50240
rect 211880 50240 212040 50400
rect 211880 50400 212040 50560
rect 211880 50560 212040 50720
rect 211880 50720 212040 50880
rect 211880 50880 212040 51040
rect 211880 51040 212040 51200
rect 211880 51200 212040 51360
rect 211880 51360 212040 51520
rect 211880 51520 212040 51680
rect 211880 51680 212040 51840
rect 211880 51840 212040 52000
rect 211880 52000 212040 52160
rect 211880 52160 212040 52320
rect 211880 52320 212040 52480
rect 211880 52480 212040 52640
rect 211880 52640 212040 52800
rect 211880 52800 212040 52960
rect 211880 52960 212040 53120
rect 211880 53120 212040 53280
rect 211880 53280 212040 53440
rect 211880 53440 212040 53600
rect 212040 47360 212200 47520
rect 212040 47520 212200 47680
rect 212040 47680 212200 47840
rect 212040 47840 212200 48000
rect 212040 48000 212200 48160
rect 212040 48160 212200 48320
rect 212040 48320 212200 48480
rect 212040 48480 212200 48640
rect 212040 48640 212200 48800
rect 212040 48800 212200 48960
rect 212040 48960 212200 49120
rect 212040 49120 212200 49280
rect 212040 49280 212200 49440
rect 212040 49440 212200 49600
rect 212040 49600 212200 49760
rect 212040 49760 212200 49920
rect 212040 49920 212200 50080
rect 212040 50080 212200 50240
rect 212040 50240 212200 50400
rect 212040 50400 212200 50560
rect 212040 50560 212200 50720
rect 212040 50720 212200 50880
rect 212040 50880 212200 51040
rect 212040 51040 212200 51200
rect 212040 51200 212200 51360
rect 212040 51360 212200 51520
rect 212040 51520 212200 51680
rect 212040 51680 212200 51840
rect 212040 51840 212200 52000
rect 212040 52000 212200 52160
rect 212040 52160 212200 52320
rect 212040 52320 212200 52480
rect 212040 52480 212200 52640
rect 212040 52640 212200 52800
rect 212040 52800 212200 52960
rect 212040 52960 212200 53120
rect 212040 53120 212200 53280
rect 212040 53280 212200 53440
rect 212200 47520 212360 47680
rect 212200 47680 212360 47840
rect 212200 47840 212360 48000
rect 212200 48000 212360 48160
rect 212200 48160 212360 48320
rect 212200 48320 212360 48480
rect 212200 48480 212360 48640
rect 212200 48640 212360 48800
rect 212200 48800 212360 48960
rect 212200 48960 212360 49120
rect 212200 49120 212360 49280
rect 212200 49280 212360 49440
rect 212200 49440 212360 49600
rect 212200 49600 212360 49760
rect 212200 49760 212360 49920
rect 212200 49920 212360 50080
rect 212200 50080 212360 50240
rect 212200 50240 212360 50400
rect 212200 50400 212360 50560
rect 212200 50560 212360 50720
rect 212200 50720 212360 50880
rect 212200 50880 212360 51040
rect 212200 51040 212360 51200
rect 212200 51200 212360 51360
rect 212200 51360 212360 51520
rect 212200 51520 212360 51680
rect 212200 51680 212360 51840
rect 212200 51840 212360 52000
rect 212200 52000 212360 52160
rect 212200 52160 212360 52320
rect 212200 52320 212360 52480
rect 212200 52480 212360 52640
rect 212200 52640 212360 52800
rect 212200 52800 212360 52960
rect 212200 52960 212360 53120
rect 212360 47680 212520 47840
rect 212360 47840 212520 48000
rect 212360 48000 212520 48160
rect 212360 48160 212520 48320
rect 212360 48320 212520 48480
rect 212360 48480 212520 48640
rect 212360 48640 212520 48800
rect 212360 48800 212520 48960
rect 212360 48960 212520 49120
rect 212360 49120 212520 49280
rect 212360 49280 212520 49440
rect 212360 49440 212520 49600
rect 212360 49600 212520 49760
rect 212360 49760 212520 49920
rect 212360 49920 212520 50080
rect 212360 50080 212520 50240
rect 212360 50240 212520 50400
rect 212360 50400 212520 50560
rect 212360 50560 212520 50720
rect 212360 50720 212520 50880
rect 212360 50880 212520 51040
rect 212360 51040 212520 51200
rect 212360 51200 212520 51360
rect 212360 51360 212520 51520
rect 212360 51520 212520 51680
rect 212360 51680 212520 51840
rect 212360 51840 212520 52000
rect 212360 52000 212520 52160
rect 212360 52160 212520 52320
rect 212360 52320 212520 52480
rect 212360 52480 212520 52640
rect 212360 52640 212520 52800
rect 212360 52800 212520 52960
rect 212520 47840 212680 48000
rect 212520 48000 212680 48160
rect 212520 48160 212680 48320
rect 212520 48320 212680 48480
rect 212520 48480 212680 48640
rect 212520 48640 212680 48800
rect 212520 48800 212680 48960
rect 212520 48960 212680 49120
rect 212520 49120 212680 49280
rect 212520 49280 212680 49440
rect 212520 49440 212680 49600
rect 212520 49600 212680 49760
rect 212520 49760 212680 49920
rect 212520 49920 212680 50080
rect 212520 50080 212680 50240
rect 212520 50240 212680 50400
rect 212520 50400 212680 50560
rect 212520 50560 212680 50720
rect 212520 50720 212680 50880
rect 212520 50880 212680 51040
rect 212520 51040 212680 51200
rect 212520 51200 212680 51360
rect 212520 51360 212680 51520
rect 212520 51520 212680 51680
rect 212520 51680 212680 51840
rect 212520 51840 212680 52000
rect 212520 52000 212680 52160
rect 212520 52160 212680 52320
rect 212520 52320 212680 52480
rect 212520 52480 212680 52640
rect 212520 52640 212680 52800
rect 212680 48000 212840 48160
rect 212680 48160 212840 48320
rect 212680 48320 212840 48480
rect 212680 48480 212840 48640
rect 212680 48640 212840 48800
rect 212680 48800 212840 48960
rect 212680 48960 212840 49120
rect 212680 49120 212840 49280
rect 212680 49280 212840 49440
rect 212680 49440 212840 49600
rect 212680 49600 212840 49760
rect 212680 49760 212840 49920
rect 212680 49920 212840 50080
rect 212680 50080 212840 50240
rect 212680 50240 212840 50400
rect 212680 50400 212840 50560
rect 212680 50560 212840 50720
rect 212680 50720 212840 50880
rect 212680 50880 212840 51040
rect 212680 51040 212840 51200
rect 212680 51200 212840 51360
rect 212680 51360 212840 51520
rect 212680 51520 212840 51680
rect 212680 51680 212840 51840
rect 212680 51840 212840 52000
rect 212680 52000 212840 52160
rect 212680 52160 212840 52320
rect 212680 52320 212840 52480
rect 212840 48320 213000 48480
rect 212840 48480 213000 48640
rect 212840 48640 213000 48800
rect 212840 48800 213000 48960
rect 212840 48960 213000 49120
rect 212840 49120 213000 49280
rect 212840 49280 213000 49440
rect 212840 49440 213000 49600
rect 212840 49600 213000 49760
rect 212840 49760 213000 49920
rect 212840 49920 213000 50080
rect 212840 50080 213000 50240
rect 212840 50240 213000 50400
rect 212840 50400 213000 50560
rect 212840 50560 213000 50720
rect 212840 50720 213000 50880
rect 212840 50880 213000 51040
rect 212840 51040 213000 51200
rect 212840 51200 213000 51360
rect 212840 51360 213000 51520
rect 212840 51520 213000 51680
rect 212840 51680 213000 51840
rect 212840 51840 213000 52000
rect 212840 52000 213000 52160
rect 213000 48640 213160 48800
rect 213000 48800 213160 48960
rect 213000 48960 213160 49120
rect 213000 49120 213160 49280
rect 213000 49280 213160 49440
rect 213000 49440 213160 49600
rect 213000 49600 213160 49760
rect 213000 49760 213160 49920
rect 213000 49920 213160 50080
rect 213000 50080 213160 50240
rect 213000 50240 213160 50400
rect 213000 50400 213160 50560
rect 213000 50560 213160 50720
rect 213000 50720 213160 50880
rect 213000 50880 213160 51040
rect 213000 51040 213160 51200
rect 213000 51200 213160 51360
rect 213000 51360 213160 51520
rect 213000 51520 213160 51680
rect 213000 51680 213160 51840
rect 213160 49120 213320 49280
rect 213160 49280 213320 49440
rect 213160 49440 213320 49600
rect 213160 49600 213320 49760
rect 213160 49760 213320 49920
rect 213160 49920 213320 50080
rect 213160 50080 213320 50240
rect 213160 50240 213320 50400
rect 213160 50400 213320 50560
rect 213160 50560 213320 50720
rect 213160 50720 213320 50880
rect 213160 50880 213320 51040
rect 213160 51040 213320 51200
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use skullfet_inverter  skullfet_inverter_0
timestamp 1640879321
transform 1 0 275500 0 1 336500
box 0 0 1070 1440
use skullfet_nand  skullfet_nand_0
timestamp 1641004779
transform 1 0 43808 0 1 324936
box 0 0 1620 1431
use skullfet_inverter_xl  skullfet_inverter_xl_0
timestamp 1641001583
transform 1 0 239740 0 1 288434
box 0 0 10700 14400
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
