magic
tech sky130A
timestamp 1640879321
<< metal1 >>
rect 47300 133000 68900 135700
rect 44600 130300 68900 133000
rect 39200 124900 74300 130300
rect 36500 114100 77000 124900
rect 36500 111400 44600 114100
rect 36500 108700 41900 111400
rect 39200 106000 41900 108700
rect 52700 106000 60800 114100
rect 68900 111400 77000 114100
rect 71600 108700 77000 111400
rect 71600 106000 74300 108700
rect 39200 103300 44600 106000
rect 50000 103300 63500 106000
rect 68900 103300 74300 106000
rect 39200 100600 55400 103300
rect 58100 100600 71600 103300
rect 44600 97900 52700 100600
rect 60800 97900 71600 100600
rect 47300 92500 66200 97900
rect 31100 89800 39200 92500
rect 47300 89800 50000 92500
rect 52700 89800 55400 92500
rect 58100 89800 60800 92500
rect 63500 89800 66200 92500
rect 74300 89800 82400 92500
rect 28400 84400 41900 89800
rect 71600 84400 85100 89800
rect 31100 81700 47300 84400
rect 66200 81700 82400 84400
rect 39200 79000 50000 81700
rect 63500 79000 74300 81700
rect 44600 76300 55400 79000
rect 58100 76300 68900 79000
rect 50000 70900 63500 76300
rect 44600 68200 55400 70900
rect 58100 68200 68900 70900
rect 31100 65500 50000 68200
rect 63500 65500 85100 68200
rect 28400 62800 44600 65500
rect 68900 62800 85100 65500
rect 28400 60100 39200 62800
rect 74300 60100 85100 62800
rect 28400 57400 36500 60100
rect 77000 57400 85100 60100
rect 31100 54700 33800 57400
rect 47300 54700 50000 57400
rect 52700 54700 55400 57400
rect 58100 54700 60800 57400
rect 63500 54700 66200 57400
rect 79700 54700 82400 57400
rect 47300 49300 66200 54700
rect 44600 46600 52700 49300
rect 60800 46600 71600 49300
rect 39200 43900 55400 46600
rect 58100 43900 71600 46600
rect 39200 41200 44600 43900
rect 50000 41200 63500 43900
rect 68900 41200 74300 43900
rect 39200 38500 41900 41200
rect 36500 35800 41900 38500
rect 36500 33100 44600 35800
rect 52700 33100 60800 41200
rect 71600 38500 74300 41200
rect 71600 35800 77000 38500
rect 68900 33100 77000 35800
rect 36500 22300 77000 33100
rect 39200 16900 74300 22300
rect 44600 14200 68900 16900
rect 47300 11500 68900 14200
<< metal2 >>
rect 47300 133000 68900 135700
rect 44600 130300 68900 133000
rect 39200 124900 74300 130300
rect 36500 114100 77000 124900
rect 36500 111400 44600 114100
rect 36500 108700 41900 111400
rect 39200 106000 41900 108700
rect 52700 106000 60800 114100
rect 68900 111400 77000 114100
rect 71600 108700 77000 111400
rect 71600 106000 74300 108700
rect 39200 103300 44600 106000
rect 50000 103300 63500 106000
rect 68900 103300 74300 106000
rect 39200 100600 55400 103300
rect 58100 100600 71600 103300
rect 44600 97900 52700 100600
rect 60800 97900 71600 100600
rect 47300 92500 66200 97900
rect 31100 89800 39200 92500
rect 47300 89800 50000 92500
rect 52700 89800 55400 92500
rect 58100 89800 60800 92500
rect 63500 89800 66200 92500
rect 74300 89800 82400 92500
rect 28400 84400 41900 89800
rect 71600 84400 85100 89800
rect 31100 81700 47300 84400
rect 66200 81700 82400 84400
rect 39200 79000 50000 81700
rect 63500 79000 74300 81700
rect 44600 76300 55400 79000
rect 58100 76300 68900 79000
rect 50000 70900 63500 76300
rect 44600 68200 55400 70900
rect 58100 68200 68900 70900
rect 31100 65500 50000 68200
rect 63500 65500 85100 68200
rect 28400 62800 44600 65500
rect 68900 62800 85100 65500
rect 28400 60100 39200 62800
rect 74300 60100 85100 62800
rect 28400 57400 36500 60100
rect 77000 57400 85100 60100
rect 31100 54700 33800 57400
rect 47300 54700 50000 57400
rect 52700 54700 55400 57400
rect 58100 54700 60800 57400
rect 63500 54700 66200 57400
rect 79700 54700 82400 57400
rect 47300 49300 66200 54700
rect 44600 46600 52700 49300
rect 60800 46600 71600 49300
rect 39200 43900 55400 46600
rect 58100 43900 71600 46600
rect 39200 41200 44600 43900
rect 50000 41200 63500 43900
rect 68900 41200 74300 43900
rect 39200 38500 41900 41200
rect 36500 35800 41900 38500
rect 36500 33100 44600 35800
rect 52700 33100 60800 41200
rect 71600 38500 74300 41200
rect 71600 35800 77000 38500
rect 68900 33100 77000 35800
rect 36500 22300 77000 33100
rect 39200 16900 74300 22300
rect 44600 14200 68900 16900
rect 47300 11500 68900 14200
<< metal3 >>
rect 47300 133000 68900 135700
rect 44600 130300 68900 133000
rect 39200 124900 74300 130300
rect 36500 114100 77000 124900
rect 36500 111400 44600 114100
rect 36500 108700 41900 111400
rect 39200 106000 41900 108700
rect 52700 106000 60800 114100
rect 68900 111400 77000 114100
rect 71600 108700 77000 111400
rect 71600 106000 74300 108700
rect 39200 103300 44600 106000
rect 50000 103300 63500 106000
rect 68900 103300 74300 106000
rect 39200 100600 55400 103300
rect 58100 100600 71600 103300
rect 44600 97900 52700 100600
rect 60800 97900 71600 100600
rect 47300 92500 66200 97900
rect 31100 89800 39200 92500
rect 47300 89800 50000 92500
rect 52700 89800 55400 92500
rect 58100 89800 60800 92500
rect 63500 89800 66200 92500
rect 74300 89800 82400 92500
rect 28400 84400 41900 89800
rect 71600 84400 85100 89800
rect 31100 81700 47300 84400
rect 66200 81700 82400 84400
rect 39200 79000 50000 81700
rect 63500 79000 74300 81700
rect 44600 76300 55400 79000
rect 58100 76300 68900 79000
rect 50000 70900 63500 76300
rect 44600 68200 55400 70900
rect 58100 68200 68900 70900
rect 31100 65500 50000 68200
rect 63500 65500 85100 68200
rect 28400 62800 44600 65500
rect 68900 62800 85100 65500
rect 28400 60100 39200 62800
rect 74300 60100 85100 62800
rect 28400 57400 36500 60100
rect 77000 57400 85100 60100
rect 31100 54700 33800 57400
rect 47300 54700 50000 57400
rect 52700 54700 55400 57400
rect 58100 54700 60800 57400
rect 63500 54700 66200 57400
rect 79700 54700 82400 57400
rect 47300 49300 66200 54700
rect 44600 46600 52700 49300
rect 60800 46600 71600 49300
rect 39200 43900 55400 46600
rect 58100 43900 71600 46600
rect 39200 41200 44600 43900
rect 50000 41200 63500 43900
rect 68900 41200 74300 43900
rect 39200 38500 41900 41200
rect 36500 35800 41900 38500
rect 36500 33100 44600 35800
rect 52700 33100 60800 41200
rect 71600 38500 74300 41200
rect 71600 35800 77000 38500
rect 68900 33100 77000 35800
rect 36500 22300 77000 33100
rect 39200 16900 74300 22300
rect 44600 14200 68900 16900
rect 47300 11500 68900 14200
<< metal4 >>
rect 47300 133000 68900 135700
rect 44600 130300 68900 133000
rect 39200 124900 74300 130300
rect 36500 114100 77000 124900
rect 36500 111400 44600 114100
rect 36500 108700 41900 111400
rect 39200 106000 41900 108700
rect 52700 106000 60800 114100
rect 68900 111400 77000 114100
rect 71600 108700 77000 111400
rect 71600 106000 74300 108700
rect 39200 103300 44600 106000
rect 50000 103300 63500 106000
rect 68900 103300 74300 106000
rect 39200 100600 55400 103300
rect 58100 100600 71600 103300
rect 44600 97900 52700 100600
rect 60800 97900 71600 100600
rect 47300 92500 66200 97900
rect 31100 89800 39200 92500
rect 47300 89800 50000 92500
rect 52700 89800 55400 92500
rect 58100 89800 60800 92500
rect 63500 89800 66200 92500
rect 74300 89800 82400 92500
rect 28400 84400 41900 89800
rect 71600 84400 85100 89800
rect 31100 81700 47300 84400
rect 66200 81700 82400 84400
rect 39200 79000 50000 81700
rect 63500 79000 74300 81700
rect 44600 76300 55400 79000
rect 58100 76300 68900 79000
rect 50000 70900 63500 76300
rect 44600 68200 55400 70900
rect 58100 68200 68900 70900
rect 31100 65500 50000 68200
rect 63500 65500 85100 68200
rect 28400 62800 44600 65500
rect 68900 62800 85100 65500
rect 28400 60100 39200 62800
rect 74300 60100 85100 62800
rect 28400 57400 36500 60100
rect 77000 57400 85100 60100
rect 31100 54700 33800 57400
rect 47300 54700 50000 57400
rect 52700 54700 55400 57400
rect 58100 54700 60800 57400
rect 63500 54700 66200 57400
rect 79700 54700 82400 57400
rect 47300 49300 66200 54700
rect 44600 46600 52700 49300
rect 60800 46600 71600 49300
rect 39200 43900 55400 46600
rect 58100 43900 71600 46600
rect 39200 41200 44600 43900
rect 50000 41200 63500 43900
rect 68900 41200 74300 43900
rect 39200 38500 41900 41200
rect 36500 35800 41900 38500
rect 36500 33100 44600 35800
rect 52700 33100 60800 41200
rect 71600 38500 74300 41200
rect 71600 35800 77000 38500
rect 68900 33100 77000 35800
rect 36500 22300 77000 33100
rect 39200 16900 74300 22300
rect 44600 14200 68900 16900
rect 47300 11500 68900 14200
<< metal5 >>
rect 47300 133000 68900 135700
rect 44600 130300 68900 133000
rect 39200 124900 74300 130300
rect 36500 114100 77000 124900
rect 36500 111400 44600 114100
rect 36500 108700 41900 111400
rect 39200 106000 41900 108700
rect 52700 106000 60800 114100
rect 68900 111400 77000 114100
rect 71600 108700 77000 111400
rect 71600 106000 74300 108700
rect 39200 103300 44600 106000
rect 50000 103300 63500 106000
rect 68900 103300 74300 106000
rect 39200 100600 55400 103300
rect 58100 100600 71600 103300
rect 44600 97900 52700 100600
rect 60800 97900 71600 100600
rect 47300 92500 66200 97900
rect 31100 89800 39200 92500
rect 47300 89800 50000 92500
rect 52700 89800 55400 92500
rect 58100 89800 60800 92500
rect 63500 89800 66200 92500
rect 74300 89800 82400 92500
rect 28400 84400 41900 89800
rect 71600 84400 85100 89800
rect 31100 81700 47300 84400
rect 66200 81700 82400 84400
rect 39200 79000 50000 81700
rect 63500 79000 74300 81700
rect 44600 76300 55400 79000
rect 58100 76300 68900 79000
rect 50000 70900 63500 76300
rect 44600 68200 55400 70900
rect 58100 68200 68900 70900
rect 31100 65500 50000 68200
rect 63500 65500 85100 68200
rect 28400 62800 44600 65500
rect 68900 62800 85100 65500
rect 28400 60100 39200 62800
rect 74300 60100 85100 62800
rect 28400 57400 36500 60100
rect 77000 57400 85100 60100
rect 31100 54700 33800 57400
rect 47300 54700 50000 57400
rect 52700 54700 55400 57400
rect 58100 54700 60800 57400
rect 63500 54700 66200 57400
rect 79700 54700 82400 57400
rect 47300 49300 66200 54700
rect 44600 46600 52700 49300
rect 60800 46600 71600 49300
rect 39200 43900 55400 46600
rect 58100 43900 71600 46600
rect 39200 41200 44600 43900
rect 50000 41200 63500 43900
rect 68900 41200 74300 43900
rect 39200 38500 41900 41200
rect 36500 35800 41900 38500
rect 36500 33100 44600 35800
rect 52700 33100 60800 41200
rect 71600 38500 74300 41200
rect 71600 35800 77000 38500
rect 68900 33100 77000 35800
rect 36500 22300 77000 33100
rect 39200 16900 74300 22300
rect 44600 14200 68900 16900
rect 47300 11500 68900 14200
<< end >>
