magic
tech sky130A
timestamp 1641003052
<< metal1 >>
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< metal2 >>
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< metal3 >>
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
rect 111182 255271 192182 260671
rect 111182 120271 116582 255271
rect 186782 120271 192182 255271
rect 111182 114871 192182 120271
<< metal4 >>
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< metal5 >>
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< end >>
