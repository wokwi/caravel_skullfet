magic
tech sky130A
timestamp 1641006614
<< locali >>
rect 44080 325330 44170 325340
rect 44080 325310 44090 325330
rect 44160 325310 44170 325330
rect 44080 325220 44170 325310
<< viali >>
rect 275750 337500 275780 337560
rect 276370 337280 276400 337320
rect 45110 326150 45140 326180
rect 45010 326030 45040 326060
rect 44090 325310 44160 325330
rect 242300 295600 242600 296200
rect 248400 295900 248700 296200
<< metal1 >>
rect 275270 338070 284400 338140
rect 284570 338070 284630 338140
rect 275270 338040 284630 338070
rect 275270 337580 275370 338040
rect 275270 337560 275790 337580
rect 275270 337500 275750 337560
rect 275780 337500 275790 337560
rect 275270 337480 275790 337500
rect 276360 337320 289100 337330
rect 276360 337280 276370 337320
rect 276400 337280 289100 337320
rect 276360 337230 289100 337280
rect 43290 326550 43510 326570
rect 43290 326460 43310 326550
rect 43470 326490 43510 326550
rect 43470 326460 45050 326490
rect 43290 326450 43510 326460
rect 45000 326060 45050 326460
rect 45100 326410 45150 326420
rect 45100 326340 45110 326410
rect 45140 326340 45150 326410
rect 45100 326180 45150 326340
rect 45100 326150 45110 326180
rect 45140 326150 45150 326180
rect 45100 326140 45150 326150
rect 45000 326030 45010 326060
rect 45040 326030 45050 326060
rect 45000 326020 45050 326030
rect 43700 325310 43710 325340
rect 43770 325330 44170 325340
rect 43770 325310 44090 325330
rect 44160 325310 44170 325330
rect 43700 325300 44170 325310
rect 248200 300400 249500 300500
rect 248200 300200 248300 300400
rect 248700 300200 249500 300400
rect 248200 300100 249500 300200
rect 249000 296300 249500 300100
rect 241400 296200 242700 296300
rect 241400 295600 241500 296200
rect 241900 295600 242300 296200
rect 242600 295600 242700 296200
rect 248300 296200 249500 296300
rect 248300 295900 248400 296200
rect 248700 295900 249500 296200
rect 248300 295800 249500 295900
rect 241400 295500 242700 295600
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< via1 >>
rect 284400 338070 284570 338140
rect 275520 337910 275590 337940
rect 275510 336500 275580 336530
rect 43310 326460 43470 326550
rect 45110 326340 45140 326410
rect 43710 325310 43770 325340
rect 45330 325120 45360 325180
rect 43910 325060 43940 325110
rect 249300 302500 250300 302700
rect 248300 300200 248700 300400
rect 241500 295600 241900 296200
rect 249200 288500 249800 288700
<< metal2 >>
rect 9350 351530 9750 351610
rect 207600 351600 208400 351700
rect 9350 351280 9450 351530
rect 9680 351280 9750 351530
rect 9350 329210 9750 351280
rect 35450 351550 35810 351600
rect 35450 351190 35490 351550
rect 35760 351190 35810 351550
rect 35450 335700 35810 351190
rect 61480 351460 61700 351500
rect 61480 351190 61500 351460
rect 61660 351190 61700 351460
rect 35430 335660 37330 335700
rect 35430 335530 43780 335660
rect 35430 335510 37330 335530
rect 9310 326570 9760 329210
rect 43680 329020 43780 335530
rect 9310 326550 43510 326570
rect 9310 326460 43310 326550
rect 43470 326460 43510 326550
rect 9310 326450 43510 326460
rect 43700 325340 43770 329020
rect 61480 326420 61700 351190
rect 45100 326410 61700 326420
rect 45100 326340 45110 326410
rect 45140 326340 61700 326410
rect 45100 326320 61700 326340
rect 207600 351300 207700 351600
rect 208300 351300 208400 351600
rect 43700 325310 43710 325340
rect 43700 325300 43770 325310
rect 45320 325180 45510 325190
rect 45320 325120 45330 325180
rect 45360 325120 45510 325180
rect 43600 325110 43950 325120
rect 43600 325060 43620 325110
rect 43730 325060 43910 325110
rect 43940 325060 43950 325110
rect 43600 325050 43950 325060
rect 45320 324240 45510 325120
rect 45320 324140 45360 324240
rect 45490 324140 45510 324240
rect 45320 323870 45510 324140
rect 207600 296300 208400 351300
rect 233500 351400 234200 351500
rect 233500 351200 233600 351400
rect 234100 351200 234200 351400
rect 233500 314400 234200 351200
rect 284360 349440 284630 349490
rect 284360 349220 284420 349440
rect 284560 349220 284630 349440
rect 284360 338140 284630 349220
rect 284360 338070 284400 338140
rect 284570 338070 284630 338140
rect 284360 338040 284630 338070
rect 288710 340370 289070 340420
rect 288710 340130 288760 340370
rect 289030 340130 289070 340370
rect 275500 338000 275600 338010
rect 275500 337950 275520 338000
rect 275580 337950 275600 338000
rect 275500 337940 275600 337950
rect 275500 337910 275520 337940
rect 275590 337910 275600 337940
rect 275500 337900 275600 337910
rect 288710 337220 289070 340130
rect 275500 336530 275590 336540
rect 275500 336500 275510 336530
rect 275580 336500 275590 336530
rect 275500 336490 275590 336500
rect 275500 336450 275520 336490
rect 275570 336450 275590 336490
rect 275500 336400 275590 336450
rect 248200 314400 248800 314500
rect 233500 313800 248800 314400
rect 248200 300400 248800 313800
rect 249200 303200 250400 303300
rect 249200 302900 249300 303200
rect 250300 302900 250400 303200
rect 249200 302700 250400 302900
rect 249200 302500 249300 302700
rect 250300 302500 250400 302700
rect 249200 302400 250400 302500
rect 248200 300200 248300 300400
rect 248700 300200 248800 300400
rect 248200 300100 248800 300200
rect 207600 296200 242000 296300
rect 207600 295600 241500 296200
rect 241900 295600 242000 296200
rect 207600 295500 242000 295600
rect 249000 288700 250000 288800
rect 249000 288500 249200 288700
rect 249800 288500 250000 288700
rect 249000 277000 250000 288500
rect 278000 277000 281000 278000
rect 249000 276000 279000 277000
rect 280000 276000 281000 277000
rect 278000 275003 281000 276000
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< via2 >>
rect 9450 351280 9680 351530
rect 35490 351190 35760 351550
rect 61500 351190 61660 351460
rect 207700 351300 208300 351600
rect 43620 325060 43730 325110
rect 45360 324140 45490 324240
rect 233600 351200 234100 351400
rect 284420 349220 284560 349440
rect 288760 340130 289030 340370
rect 275520 337950 275580 338000
rect 275520 336450 275570 336490
rect 249300 302900 250300 303200
rect 279000 276000 280000 277000
<< metal3 >>
rect 8097 351530 10597 352400
rect 8097 351280 9450 351530
rect 9680 351280 10597 351530
rect 8097 351150 10597 351280
rect 34097 351550 36597 352400
rect 34097 351190 35490 351550
rect 35760 351190 36597 351550
rect 34097 351150 36597 351190
rect 60097 351460 62597 352400
rect 60097 351190 61500 351460
rect 61660 351190 62597 351460
rect 60097 351150 62597 351190
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351600 209197 352400
rect 206697 351300 207700 351600
rect 208300 351300 209197 351600
rect 206697 351150 209197 351300
rect 232697 351400 235197 352400
rect 232697 351200 233600 351400
rect 234100 351200 235197 351400
rect 232697 351150 235197 351200
rect 255297 351500 257697 352400
rect 260297 351500 262697 352400
rect 255297 351170 257700 351500
rect 260297 351170 262700 351500
rect 255300 350407 257700 351170
rect 255275 349200 257700 350407
rect 260300 349200 262700 351170
rect 283297 351150 285797 352400
rect 255275 348040 262700 349200
rect 284300 349440 284700 351150
rect 284300 349220 284420 349440
rect 284560 349220 284700 349440
rect 284300 348800 284700 349220
rect 274710 348040 275610 348050
rect 255275 347500 275610 348040
rect -400 340121 850 342621
rect 43480 331950 43760 331960
rect 255275 331950 256842 347500
rect 260660 347490 275610 347500
rect 275460 338000 275610 347490
rect 291150 340400 292400 341492
rect 288600 340370 292400 340400
rect 288600 340130 288760 340370
rect 289030 340130 292400 340370
rect 288600 340100 292400 340130
rect 291150 338992 292400 340100
rect 275460 337950 275520 338000
rect 275580 337950 275610 338000
rect 275460 337930 275610 337950
rect 275300 336490 275900 336500
rect 275300 336450 275520 336490
rect 275570 336450 275900 336490
rect 43480 330700 256860 331950
rect 43480 330340 43760 330700
rect 43490 325110 43750 330340
rect 43490 325060 43620 325110
rect 43730 325060 43750 325110
rect 43490 325050 43750 325060
rect -400 321921 830 324321
rect 45300 324240 45970 324260
rect 45300 324140 45360 324240
rect 45490 324140 45970 324240
rect -400 316921 830 319321
rect 45300 284100 45970 324140
rect 255275 307400 256842 330700
rect 255300 307300 256842 307400
rect 249200 305900 256842 307300
rect 249200 303200 250400 305900
rect 249200 302900 249300 303200
rect 250300 302900 250400 303200
rect 249200 302600 250400 302900
rect 45260 284050 66400 284100
rect 275300 284050 275900 336450
rect 291170 319892 292400 322292
rect 291170 314892 292400 317292
rect 291760 294736 292400 294792
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 291760 292372 292400 292428
rect 291760 291781 292400 291837
rect 45260 282800 276000 284050
rect 45260 282780 66400 282800
rect -400 279721 830 282121
rect 275300 277800 275900 282800
rect 275300 277700 290300 277800
rect 275300 277681 291800 277700
rect -400 274721 830 277121
rect 275300 277000 292400 277681
rect 275300 276000 279000 277000
rect 280000 276000 292400 277000
rect 275300 275300 292400 276000
rect 275300 275200 290300 275300
rect 291170 275281 292400 275300
rect 287300 272700 288370 275200
rect 287300 272681 291800 272700
rect 287300 270300 292400 272681
rect 287300 270290 288370 270300
rect 291170 270281 292400 270300
rect -400 255765 240 255821
rect 111182 255271 192182 260671
rect -400 255174 240 255230
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect -400 234154 240 234210
rect -400 233563 240 233619
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect -400 212543 240 212599
rect -400 211952 240 212008
rect -400 211361 240 211417
rect -400 210770 240 210826
rect -400 210179 240 210235
rect -400 209588 240 209644
rect -400 190932 240 190988
rect -400 190341 240 190397
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect -400 169321 240 169377
rect -400 168730 240 168786
rect -400 168139 240 168195
rect -400 167548 240 167604
rect -400 166957 240 167013
rect -400 166366 240 166422
rect -400 147710 240 147766
rect -400 147119 240 147175
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect -400 126199 240 126255
rect -400 125608 240 125664
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect 111182 120271 116582 255271
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
rect 186782 120271 192182 255271
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect 291760 227814 292400 227870
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 291760 202648 292400 202704
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 291760 179437 292400 179493
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect 291760 137570 292400 137626
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect 111182 114871 192182 120271
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect -400 107444 830 109844
rect -400 102444 830 104844
rect 291170 95715 292400 98115
rect 291170 90715 292400 93115
rect -400 86444 830 88844
rect -400 81444 830 83844
rect 291170 73415 292400 75815
rect 291170 68415 292400 70815
rect -400 62388 240 62444
rect -400 61797 240 61853
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect -400 40777 240 40833
rect -400 40186 240 40242
rect -400 39595 240 39651
rect -400 39004 240 39060
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect -400 19166 240 19222
rect -400 18575 240 18631
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect -400 8455 240 8511
rect 291760 8455 292400 8511
rect -400 7864 240 7920
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< metal4 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 142282 247871 163882 250571
rect 139582 245171 163882 247871
rect 134182 239771 169282 245171
rect 131482 228971 171982 239771
rect 131482 226271 139582 228971
rect 131482 223571 136882 226271
rect 134182 220871 136882 223571
rect 147682 220871 155782 228971
rect 163882 226271 171982 228971
rect 166582 223571 171982 226271
rect 166582 220871 169282 223571
rect 134182 218171 139582 220871
rect 144982 218171 158482 220871
rect 163882 218171 169282 220871
rect 134182 215471 150382 218171
rect 153082 215471 166582 218171
rect 139582 212771 147682 215471
rect 155782 212771 166582 215471
rect 142282 207371 161182 212771
rect 126082 204671 134182 207371
rect 142282 204671 144982 207371
rect 147682 204671 150382 207371
rect 153082 204671 155782 207371
rect 158482 204671 161182 207371
rect 169282 204671 177382 207371
rect 123382 199271 136882 204671
rect 166582 199271 180082 204671
rect 126082 196571 142282 199271
rect 161182 196571 177382 199271
rect 134182 193871 144982 196571
rect 158482 193871 169282 196571
rect 139582 191171 150382 193871
rect 153082 191171 163882 193871
rect 144982 185771 158482 191171
rect 139582 183071 150382 185771
rect 153082 183071 163882 185771
rect 126082 180371 144982 183071
rect 158482 180371 180082 183071
rect 123382 177671 139582 180371
rect 163882 177671 180082 180371
rect 123382 174971 134182 177671
rect 169282 174971 180082 177671
rect 123382 172271 131482 174971
rect 171982 172271 180082 174971
rect 126082 169571 128782 172271
rect 142282 169571 144982 172271
rect 147682 169571 150382 172271
rect 153082 169571 155782 172271
rect 158482 169571 161182 172271
rect 174682 169571 177382 172271
rect 142282 164171 161182 169571
rect 139582 161471 147682 164171
rect 155782 161471 166582 164171
rect 134182 158771 150382 161471
rect 153082 158771 166582 161471
rect 134182 156071 139582 158771
rect 144982 156071 158482 158771
rect 163882 156071 169282 158771
rect 134182 153371 136882 156071
rect 131482 150671 136882 153371
rect 131482 147971 139582 150671
rect 147682 147971 155782 156071
rect 166582 153371 169282 156071
rect 166582 150671 171982 153371
rect 163882 147971 171982 150671
rect 131482 137171 171982 147971
rect 134182 131771 169282 137171
rect 139582 129071 163882 131771
rect 142282 126371 163882 129071
<< metal4 >>
rect 110800 35500 110900 35600
rect 110900 34800 111000 34900
rect 110900 34900 111000 35000
rect 110900 35000 111000 35100
rect 110900 35100 111000 35200
rect 110900 35200 111000 35300
rect 110900 35300 111000 35400
rect 110900 35400 111000 35500
rect 110900 35500 111000 35600
rect 110900 35600 111000 35700
rect 110900 35700 111000 35800
rect 110900 35800 111000 35900
rect 110900 35900 111000 36000
rect 110900 36000 111000 36100
rect 111000 34500 111100 34600
rect 111000 34600 111100 34700
rect 111000 34700 111100 34800
rect 111000 34800 111100 34900
rect 111000 34900 111100 35000
rect 111000 35000 111100 35100
rect 111000 35100 111100 35200
rect 111000 35200 111100 35300
rect 111000 35300 111100 35400
rect 111000 35400 111100 35500
rect 111000 35500 111100 35600
rect 111000 35600 111100 35700
rect 111000 35700 111100 35800
rect 111000 35800 111100 35900
rect 111000 35900 111100 36000
rect 111000 36000 111100 36100
rect 111000 36100 111100 36200
rect 111000 36200 111100 36300
rect 111000 36300 111100 36400
rect 111100 34300 111200 34400
rect 111100 34400 111200 34500
rect 111100 34500 111200 34600
rect 111100 34600 111200 34700
rect 111100 34700 111200 34800
rect 111100 34800 111200 34900
rect 111100 34900 111200 35000
rect 111100 35000 111200 35100
rect 111100 35100 111200 35200
rect 111100 35200 111200 35300
rect 111100 35300 111200 35400
rect 111100 35400 111200 35500
rect 111100 35500 111200 35600
rect 111100 35600 111200 35700
rect 111100 35700 111200 35800
rect 111100 35800 111200 35900
rect 111100 35900 111200 36000
rect 111100 36000 111200 36100
rect 111100 36100 111200 36200
rect 111100 36200 111200 36300
rect 111100 36300 111200 36400
rect 111100 36400 111200 36500
rect 111100 36500 111200 36600
rect 111200 34100 111300 34200
rect 111200 34200 111300 34300
rect 111200 34300 111300 34400
rect 111200 34400 111300 34500
rect 111200 34500 111300 34600
rect 111200 34600 111300 34700
rect 111200 34700 111300 34800
rect 111200 34800 111300 34900
rect 111200 34900 111300 35000
rect 111200 35000 111300 35100
rect 111200 35100 111300 35200
rect 111200 35200 111300 35300
rect 111200 35300 111300 35400
rect 111200 35400 111300 35500
rect 111200 35500 111300 35600
rect 111200 35600 111300 35700
rect 111200 35700 111300 35800
rect 111200 35800 111300 35900
rect 111200 35900 111300 36000
rect 111200 36000 111300 36100
rect 111200 36100 111300 36200
rect 111200 36200 111300 36300
rect 111200 36300 111300 36400
rect 111200 36400 111300 36500
rect 111200 36500 111300 36600
rect 111200 36600 111300 36700
rect 111300 34000 111400 34100
rect 111300 34100 111400 34200
rect 111300 34200 111400 34300
rect 111300 34300 111400 34400
rect 111300 34400 111400 34500
rect 111300 34500 111400 34600
rect 111300 34600 111400 34700
rect 111300 34700 111400 34800
rect 111300 34800 111400 34900
rect 111300 34900 111400 35000
rect 111300 35000 111400 35100
rect 111300 35100 111400 35200
rect 111300 35200 111400 35300
rect 111300 35300 111400 35400
rect 111300 35400 111400 35500
rect 111300 35500 111400 35600
rect 111300 35600 111400 35700
rect 111300 35700 111400 35800
rect 111300 35800 111400 35900
rect 111300 35900 111400 36000
rect 111300 36000 111400 36100
rect 111300 36100 111400 36200
rect 111300 36200 111400 36300
rect 111300 36300 111400 36400
rect 111300 36400 111400 36500
rect 111300 36500 111400 36600
rect 111300 36600 111400 36700
rect 111300 36700 111400 36800
rect 111300 36800 111400 36900
rect 111400 33900 111500 34000
rect 111400 34000 111500 34100
rect 111400 34100 111500 34200
rect 111400 34200 111500 34300
rect 111400 34300 111500 34400
rect 111400 34400 111500 34500
rect 111400 34500 111500 34600
rect 111400 34600 111500 34700
rect 111400 34700 111500 34800
rect 111400 34800 111500 34900
rect 111400 34900 111500 35000
rect 111400 35000 111500 35100
rect 111400 35100 111500 35200
rect 111400 35200 111500 35300
rect 111400 35300 111500 35400
rect 111400 35400 111500 35500
rect 111400 35500 111500 35600
rect 111400 35600 111500 35700
rect 111400 35700 111500 35800
rect 111400 35800 111500 35900
rect 111400 35900 111500 36000
rect 111400 36000 111500 36100
rect 111400 36100 111500 36200
rect 111400 36200 111500 36300
rect 111400 36300 111500 36400
rect 111400 36400 111500 36500
rect 111400 36500 111500 36600
rect 111400 36600 111500 36700
rect 111400 36700 111500 36800
rect 111400 36800 111500 36900
rect 111400 36900 111500 37000
rect 111500 33800 111600 33900
rect 111500 33900 111600 34000
rect 111500 34000 111600 34100
rect 111500 34100 111600 34200
rect 111500 34200 111600 34300
rect 111500 34300 111600 34400
rect 111500 34400 111600 34500
rect 111500 34500 111600 34600
rect 111500 34600 111600 34700
rect 111500 34700 111600 34800
rect 111500 34800 111600 34900
rect 111500 34900 111600 35000
rect 111500 35000 111600 35100
rect 111500 35100 111600 35200
rect 111500 35200 111600 35300
rect 111500 35300 111600 35400
rect 111500 35400 111600 35500
rect 111500 35500 111600 35600
rect 111500 35600 111600 35700
rect 111500 35700 111600 35800
rect 111500 35800 111600 35900
rect 111500 35900 111600 36000
rect 111500 36000 111600 36100
rect 111500 36100 111600 36200
rect 111500 36200 111600 36300
rect 111500 36300 111600 36400
rect 111500 36400 111600 36500
rect 111500 36500 111600 36600
rect 111500 36600 111600 36700
rect 111500 36700 111600 36800
rect 111500 36800 111600 36900
rect 111500 36900 111600 37000
rect 111500 37000 111600 37100
rect 111600 33600 111700 33700
rect 111600 33700 111700 33800
rect 111600 33800 111700 33900
rect 111600 33900 111700 34000
rect 111600 34000 111700 34100
rect 111600 34100 111700 34200
rect 111600 34200 111700 34300
rect 111600 34300 111700 34400
rect 111600 34400 111700 34500
rect 111600 34500 111700 34600
rect 111600 34600 111700 34700
rect 111600 34700 111700 34800
rect 111600 34800 111700 34900
rect 111600 34900 111700 35000
rect 111600 35000 111700 35100
rect 111600 35100 111700 35200
rect 111600 35200 111700 35300
rect 111600 35300 111700 35400
rect 111600 35400 111700 35500
rect 111600 35500 111700 35600
rect 111600 35600 111700 35700
rect 111600 35700 111700 35800
rect 111600 35800 111700 35900
rect 111600 35900 111700 36000
rect 111600 36000 111700 36100
rect 111600 36100 111700 36200
rect 111600 36200 111700 36300
rect 111600 36300 111700 36400
rect 111600 36400 111700 36500
rect 111600 36500 111700 36600
rect 111600 36600 111700 36700
rect 111600 36700 111700 36800
rect 111600 36800 111700 36900
rect 111600 36900 111700 37000
rect 111600 37000 111700 37100
rect 111600 37100 111700 37200
rect 111700 33600 111800 33700
rect 111700 33700 111800 33800
rect 111700 33800 111800 33900
rect 111700 33900 111800 34000
rect 111700 34000 111800 34100
rect 111700 34100 111800 34200
rect 111700 34200 111800 34300
rect 111700 34300 111800 34400
rect 111700 34400 111800 34500
rect 111700 34500 111800 34600
rect 111700 34600 111800 34700
rect 111700 34700 111800 34800
rect 111700 34800 111800 34900
rect 111700 34900 111800 35000
rect 111700 35000 111800 35100
rect 111700 35100 111800 35200
rect 111700 35200 111800 35300
rect 111700 35300 111800 35400
rect 111700 35400 111800 35500
rect 111700 35500 111800 35600
rect 111700 35600 111800 35700
rect 111700 35700 111800 35800
rect 111700 35800 111800 35900
rect 111700 35900 111800 36000
rect 111700 36000 111800 36100
rect 111700 36100 111800 36200
rect 111700 36200 111800 36300
rect 111700 36300 111800 36400
rect 111700 36400 111800 36500
rect 111700 36500 111800 36600
rect 111700 36600 111800 36700
rect 111700 36700 111800 36800
rect 111700 36800 111800 36900
rect 111700 36900 111800 37000
rect 111700 37000 111800 37100
rect 111700 37100 111800 37200
rect 111700 37200 111800 37300
rect 111800 33500 111900 33600
rect 111800 33600 111900 33700
rect 111800 33700 111900 33800
rect 111800 33800 111900 33900
rect 111800 33900 111900 34000
rect 111800 34000 111900 34100
rect 111800 34100 111900 34200
rect 111800 34200 111900 34300
rect 111800 34300 111900 34400
rect 111800 34400 111900 34500
rect 111800 34500 111900 34600
rect 111800 34600 111900 34700
rect 111800 34700 111900 34800
rect 111800 34800 111900 34900
rect 111800 34900 111900 35000
rect 111800 35000 111900 35100
rect 111800 35100 111900 35200
rect 111800 35200 111900 35300
rect 111800 35300 111900 35400
rect 111800 35400 111900 35500
rect 111800 35500 111900 35600
rect 111800 35600 111900 35700
rect 111800 35700 111900 35800
rect 111800 35800 111900 35900
rect 111800 35900 111900 36000
rect 111800 36000 111900 36100
rect 111800 36100 111900 36200
rect 111800 36200 111900 36300
rect 111800 36300 111900 36400
rect 111800 36400 111900 36500
rect 111800 36500 111900 36600
rect 111800 36600 111900 36700
rect 111800 36700 111900 36800
rect 111800 36800 111900 36900
rect 111800 36900 111900 37000
rect 111800 37000 111900 37100
rect 111800 37100 111900 37200
rect 111800 37200 111900 37300
rect 111900 33400 112000 33500
rect 111900 33500 112000 33600
rect 111900 33600 112000 33700
rect 111900 33700 112000 33800
rect 111900 33800 112000 33900
rect 111900 33900 112000 34000
rect 111900 34000 112000 34100
rect 111900 34100 112000 34200
rect 111900 34200 112000 34300
rect 111900 34300 112000 34400
rect 111900 34400 112000 34500
rect 111900 34500 112000 34600
rect 111900 34600 112000 34700
rect 111900 34700 112000 34800
rect 111900 34800 112000 34900
rect 111900 34900 112000 35000
rect 111900 35000 112000 35100
rect 111900 35100 112000 35200
rect 111900 35200 112000 35300
rect 111900 35300 112000 35400
rect 111900 35400 112000 35500
rect 111900 35500 112000 35600
rect 111900 35600 112000 35700
rect 111900 35700 112000 35800
rect 111900 35800 112000 35900
rect 111900 35900 112000 36000
rect 111900 36000 112000 36100
rect 111900 36100 112000 36200
rect 111900 36200 112000 36300
rect 111900 36300 112000 36400
rect 111900 36400 112000 36500
rect 111900 36500 112000 36600
rect 111900 36600 112000 36700
rect 111900 36700 112000 36800
rect 111900 36800 112000 36900
rect 111900 36900 112000 37000
rect 111900 37000 112000 37100
rect 111900 37100 112000 37200
rect 111900 37200 112000 37300
rect 111900 37300 112000 37400
rect 112000 33300 112100 33400
rect 112000 33400 112100 33500
rect 112000 33500 112100 33600
rect 112000 33600 112100 33700
rect 112000 33700 112100 33800
rect 112000 33800 112100 33900
rect 112000 33900 112100 34000
rect 112000 34000 112100 34100
rect 112000 34100 112100 34200
rect 112000 34200 112100 34300
rect 112000 34300 112100 34400
rect 112000 34400 112100 34500
rect 112000 34500 112100 34600
rect 112000 34600 112100 34700
rect 112000 34700 112100 34800
rect 112000 34800 112100 34900
rect 112000 34900 112100 35000
rect 112000 35000 112100 35100
rect 112000 35100 112100 35200
rect 112000 35200 112100 35300
rect 112000 35300 112100 35400
rect 112000 35400 112100 35500
rect 112000 35500 112100 35600
rect 112000 35600 112100 35700
rect 112000 35700 112100 35800
rect 112000 35800 112100 35900
rect 112000 35900 112100 36000
rect 112000 36000 112100 36100
rect 112000 36100 112100 36200
rect 112000 36200 112100 36300
rect 112000 36300 112100 36400
rect 112000 36400 112100 36500
rect 112000 36500 112100 36600
rect 112000 36600 112100 36700
rect 112000 36700 112100 36800
rect 112000 36800 112100 36900
rect 112000 36900 112100 37000
rect 112000 37000 112100 37100
rect 112000 37100 112100 37200
rect 112000 37200 112100 37300
rect 112000 37300 112100 37400
rect 112000 37400 112100 37500
rect 112100 33300 112200 33400
rect 112100 33400 112200 33500
rect 112100 33500 112200 33600
rect 112100 33600 112200 33700
rect 112100 33700 112200 33800
rect 112100 33800 112200 33900
rect 112100 33900 112200 34000
rect 112100 34000 112200 34100
rect 112100 34100 112200 34200
rect 112100 34200 112200 34300
rect 112100 34300 112200 34400
rect 112100 34400 112200 34500
rect 112100 34500 112200 34600
rect 112100 34600 112200 34700
rect 112100 34700 112200 34800
rect 112100 34800 112200 34900
rect 112100 34900 112200 35000
rect 112100 35000 112200 35100
rect 112100 35100 112200 35200
rect 112100 35200 112200 35300
rect 112100 35300 112200 35400
rect 112100 35400 112200 35500
rect 112100 35500 112200 35600
rect 112100 35600 112200 35700
rect 112100 35700 112200 35800
rect 112100 35800 112200 35900
rect 112100 35900 112200 36000
rect 112100 36000 112200 36100
rect 112100 36100 112200 36200
rect 112100 36200 112200 36300
rect 112100 36300 112200 36400
rect 112100 36400 112200 36500
rect 112100 36500 112200 36600
rect 112100 36600 112200 36700
rect 112100 36700 112200 36800
rect 112100 36800 112200 36900
rect 112100 36900 112200 37000
rect 112100 37000 112200 37100
rect 112100 37100 112200 37200
rect 112100 37200 112200 37300
rect 112100 37300 112200 37400
rect 112100 37400 112200 37500
rect 112200 33200 112300 33300
rect 112200 33300 112300 33400
rect 112200 33400 112300 33500
rect 112200 33500 112300 33600
rect 112200 33600 112300 33700
rect 112200 33700 112300 33800
rect 112200 33800 112300 33900
rect 112200 33900 112300 34000
rect 112200 34000 112300 34100
rect 112200 34100 112300 34200
rect 112200 34200 112300 34300
rect 112200 34300 112300 34400
rect 112200 34400 112300 34500
rect 112200 34500 112300 34600
rect 112200 34600 112300 34700
rect 112200 34700 112300 34800
rect 112200 34800 112300 34900
rect 112200 34900 112300 35000
rect 112200 35000 112300 35100
rect 112200 35100 112300 35200
rect 112200 35200 112300 35300
rect 112200 35300 112300 35400
rect 112200 35400 112300 35500
rect 112200 35500 112300 35600
rect 112200 35600 112300 35700
rect 112200 35700 112300 35800
rect 112200 35800 112300 35900
rect 112200 35900 112300 36000
rect 112200 36000 112300 36100
rect 112200 36100 112300 36200
rect 112200 36200 112300 36300
rect 112200 36300 112300 36400
rect 112200 36400 112300 36500
rect 112200 36500 112300 36600
rect 112200 36600 112300 36700
rect 112200 36700 112300 36800
rect 112200 36800 112300 36900
rect 112200 36900 112300 37000
rect 112200 37000 112300 37100
rect 112200 37100 112300 37200
rect 112200 37200 112300 37300
rect 112200 37300 112300 37400
rect 112200 37400 112300 37500
rect 112200 37500 112300 37600
rect 112300 33200 112400 33300
rect 112300 33300 112400 33400
rect 112300 33400 112400 33500
rect 112300 33500 112400 33600
rect 112300 33600 112400 33700
rect 112300 33700 112400 33800
rect 112300 33800 112400 33900
rect 112300 33900 112400 34000
rect 112300 34000 112400 34100
rect 112300 34100 112400 34200
rect 112300 34200 112400 34300
rect 112300 34300 112400 34400
rect 112300 34400 112400 34500
rect 112300 34500 112400 34600
rect 112300 34600 112400 34700
rect 112300 34700 112400 34800
rect 112300 34800 112400 34900
rect 112300 34900 112400 35000
rect 112300 35000 112400 35100
rect 112300 35100 112400 35200
rect 112300 35200 112400 35300
rect 112300 35300 112400 35400
rect 112300 35400 112400 35500
rect 112300 35500 112400 35600
rect 112300 35600 112400 35700
rect 112300 35700 112400 35800
rect 112300 35800 112400 35900
rect 112300 35900 112400 36000
rect 112300 36000 112400 36100
rect 112300 36100 112400 36200
rect 112300 36200 112400 36300
rect 112300 36300 112400 36400
rect 112300 36400 112400 36500
rect 112300 36500 112400 36600
rect 112300 36600 112400 36700
rect 112300 36700 112400 36800
rect 112300 36800 112400 36900
rect 112300 36900 112400 37000
rect 112300 37000 112400 37100
rect 112300 37100 112400 37200
rect 112300 37200 112400 37300
rect 112300 37300 112400 37400
rect 112300 37400 112400 37500
rect 112300 37500 112400 37600
rect 112400 33100 112500 33200
rect 112400 33200 112500 33300
rect 112400 33300 112500 33400
rect 112400 33400 112500 33500
rect 112400 33500 112500 33600
rect 112400 33600 112500 33700
rect 112400 33700 112500 33800
rect 112400 33800 112500 33900
rect 112400 33900 112500 34000
rect 112400 34000 112500 34100
rect 112400 34100 112500 34200
rect 112400 34200 112500 34300
rect 112400 34300 112500 34400
rect 112400 34400 112500 34500
rect 112400 34500 112500 34600
rect 112400 34600 112500 34700
rect 112400 34700 112500 34800
rect 112400 34800 112500 34900
rect 112400 34900 112500 35000
rect 112400 35000 112500 35100
rect 112400 35100 112500 35200
rect 112400 35200 112500 35300
rect 112400 35300 112500 35400
rect 112400 35400 112500 35500
rect 112400 35500 112500 35600
rect 112400 35600 112500 35700
rect 112400 35700 112500 35800
rect 112400 35800 112500 35900
rect 112400 35900 112500 36000
rect 112400 36000 112500 36100
rect 112400 36100 112500 36200
rect 112400 36200 112500 36300
rect 112400 36300 112500 36400
rect 112400 36400 112500 36500
rect 112400 36500 112500 36600
rect 112400 36600 112500 36700
rect 112400 36700 112500 36800
rect 112400 36800 112500 36900
rect 112400 36900 112500 37000
rect 112400 37000 112500 37100
rect 112400 37100 112500 37200
rect 112400 37200 112500 37300
rect 112400 37300 112500 37400
rect 112400 37400 112500 37500
rect 112400 37500 112500 37600
rect 112500 33000 112600 33100
rect 112500 33100 112600 33200
rect 112500 33200 112600 33300
rect 112500 33300 112600 33400
rect 112500 33400 112600 33500
rect 112500 33500 112600 33600
rect 112500 33600 112600 33700
rect 112500 33700 112600 33800
rect 112500 33800 112600 33900
rect 112500 33900 112600 34000
rect 112500 34000 112600 34100
rect 112500 34100 112600 34200
rect 112500 34200 112600 34300
rect 112500 34300 112600 34400
rect 112500 34400 112600 34500
rect 112500 34500 112600 34600
rect 112500 34600 112600 34700
rect 112500 34700 112600 34800
rect 112500 34800 112600 34900
rect 112500 34900 112600 35000
rect 112500 35000 112600 35100
rect 112500 35100 112600 35200
rect 112500 35200 112600 35300
rect 112500 35600 112600 35700
rect 112500 35700 112600 35800
rect 112500 35800 112600 35900
rect 112500 35900 112600 36000
rect 112500 36000 112600 36100
rect 112500 36100 112600 36200
rect 112500 36200 112600 36300
rect 112500 36300 112600 36400
rect 112500 36400 112600 36500
rect 112500 36500 112600 36600
rect 112500 36600 112600 36700
rect 112500 36700 112600 36800
rect 112500 36800 112600 36900
rect 112500 36900 112600 37000
rect 112500 37000 112600 37100
rect 112500 37100 112600 37200
rect 112500 37200 112600 37300
rect 112500 37300 112600 37400
rect 112500 37400 112600 37500
rect 112500 37500 112600 37600
rect 112500 37600 112600 37700
rect 112600 33000 112700 33100
rect 112600 33100 112700 33200
rect 112600 33200 112700 33300
rect 112600 33300 112700 33400
rect 112600 33400 112700 33500
rect 112600 33500 112700 33600
rect 112600 33600 112700 33700
rect 112600 33700 112700 33800
rect 112600 33800 112700 33900
rect 112600 33900 112700 34000
rect 112600 34000 112700 34100
rect 112600 34100 112700 34200
rect 112600 34200 112700 34300
rect 112600 34300 112700 34400
rect 112600 34400 112700 34500
rect 112600 34500 112700 34600
rect 112600 34600 112700 34700
rect 112600 34700 112700 34800
rect 112600 34800 112700 34900
rect 112600 34900 112700 35000
rect 112600 35000 112700 35100
rect 112600 35800 112700 35900
rect 112600 35900 112700 36000
rect 112600 36000 112700 36100
rect 112600 36100 112700 36200
rect 112600 36200 112700 36300
rect 112600 36300 112700 36400
rect 112600 36400 112700 36500
rect 112600 36500 112700 36600
rect 112600 36600 112700 36700
rect 112600 36700 112700 36800
rect 112600 36800 112700 36900
rect 112600 36900 112700 37000
rect 112600 37000 112700 37100
rect 112600 37100 112700 37200
rect 112600 37200 112700 37300
rect 112600 37300 112700 37400
rect 112600 37400 112700 37500
rect 112600 37500 112700 37600
rect 112600 37600 112700 37700
rect 112700 32900 112800 33000
rect 112700 33000 112800 33100
rect 112700 33100 112800 33200
rect 112700 33200 112800 33300
rect 112700 33300 112800 33400
rect 112700 33400 112800 33500
rect 112700 33500 112800 33600
rect 112700 33600 112800 33700
rect 112700 33700 112800 33800
rect 112700 33800 112800 33900
rect 112700 33900 112800 34000
rect 112700 34000 112800 34100
rect 112700 34100 112800 34200
rect 112700 34200 112800 34300
rect 112700 34300 112800 34400
rect 112700 34400 112800 34500
rect 112700 34500 112800 34600
rect 112700 34600 112800 34700
rect 112700 34700 112800 34800
rect 112700 34800 112800 34900
rect 112700 34900 112800 35000
rect 112700 35900 112800 36000
rect 112700 36000 112800 36100
rect 112700 36100 112800 36200
rect 112700 36200 112800 36300
rect 112700 36300 112800 36400
rect 112700 36400 112800 36500
rect 112700 36500 112800 36600
rect 112700 36600 112800 36700
rect 112700 36700 112800 36800
rect 112700 36800 112800 36900
rect 112700 36900 112800 37000
rect 112700 37000 112800 37100
rect 112700 37100 112800 37200
rect 112700 37200 112800 37300
rect 112700 37300 112800 37400
rect 112700 37400 112800 37500
rect 112700 37500 112800 37600
rect 112700 37600 112800 37700
rect 112800 32900 112900 33000
rect 112800 33000 112900 33100
rect 112800 33100 112900 33200
rect 112800 33200 112900 33300
rect 112800 33300 112900 33400
rect 112800 33400 112900 33500
rect 112800 33500 112900 33600
rect 112800 33600 112900 33700
rect 112800 33700 112900 33800
rect 112800 33800 112900 33900
rect 112800 33900 112900 34000
rect 112800 34000 112900 34100
rect 112800 34100 112900 34200
rect 112800 34200 112900 34300
rect 112800 34300 112900 34400
rect 112800 34400 112900 34500
rect 112800 34500 112900 34600
rect 112800 34600 112900 34700
rect 112800 34700 112900 34800
rect 112800 34800 112900 34900
rect 112800 36000 112900 36100
rect 112800 36100 112900 36200
rect 112800 36200 112900 36300
rect 112800 36300 112900 36400
rect 112800 36400 112900 36500
rect 112800 36500 112900 36600
rect 112800 36600 112900 36700
rect 112800 36700 112900 36800
rect 112800 36800 112900 36900
rect 112800 36900 112900 37000
rect 112800 37000 112900 37100
rect 112800 37100 112900 37200
rect 112800 37200 112900 37300
rect 112800 37300 112900 37400
rect 112800 37400 112900 37500
rect 112800 37500 112900 37600
rect 112800 37600 112900 37700
rect 112900 32800 113000 32900
rect 112900 32900 113000 33000
rect 112900 33000 113000 33100
rect 112900 33100 113000 33200
rect 112900 33200 113000 33300
rect 112900 33300 113000 33400
rect 112900 33400 113000 33500
rect 112900 33500 113000 33600
rect 112900 33600 113000 33700
rect 112900 33700 113000 33800
rect 112900 33800 113000 33900
rect 112900 33900 113000 34000
rect 112900 34000 113000 34100
rect 112900 34100 113000 34200
rect 112900 34200 113000 34300
rect 112900 34300 113000 34400
rect 112900 34400 113000 34500
rect 112900 34500 113000 34600
rect 112900 34600 113000 34700
rect 112900 34700 113000 34800
rect 112900 34800 113000 34900
rect 112900 36100 113000 36200
rect 112900 36200 113000 36300
rect 112900 36300 113000 36400
rect 112900 36400 113000 36500
rect 112900 36500 113000 36600
rect 112900 36600 113000 36700
rect 112900 36700 113000 36800
rect 112900 36800 113000 36900
rect 112900 36900 113000 37000
rect 112900 37000 113000 37100
rect 112900 37100 113000 37200
rect 112900 37200 113000 37300
rect 112900 37300 113000 37400
rect 112900 37400 113000 37500
rect 112900 37500 113000 37600
rect 112900 37600 113000 37700
rect 112900 37700 113000 37800
rect 113000 32700 113100 32800
rect 113000 32800 113100 32900
rect 113000 32900 113100 33000
rect 113000 33000 113100 33100
rect 113000 33100 113100 33200
rect 113000 33200 113100 33300
rect 113000 33300 113100 33400
rect 113000 33400 113100 33500
rect 113000 33500 113100 33600
rect 113000 33600 113100 33700
rect 113000 33700 113100 33800
rect 113000 33800 113100 33900
rect 113000 33900 113100 34000
rect 113000 34000 113100 34100
rect 113000 34100 113100 34200
rect 113000 34200 113100 34300
rect 113000 34300 113100 34400
rect 113000 34400 113100 34500
rect 113000 34500 113100 34600
rect 113000 34600 113100 34700
rect 113000 34700 113100 34800
rect 113000 36100 113100 36200
rect 113000 36200 113100 36300
rect 113000 36300 113100 36400
rect 113000 36400 113100 36500
rect 113000 36500 113100 36600
rect 113000 36600 113100 36700
rect 113000 36700 113100 36800
rect 113000 36800 113100 36900
rect 113000 36900 113100 37000
rect 113000 37000 113100 37100
rect 113000 37100 113100 37200
rect 113000 37200 113100 37300
rect 113000 37300 113100 37400
rect 113000 37400 113100 37500
rect 113000 37500 113100 37600
rect 113000 37600 113100 37700
rect 113000 37700 113100 37800
rect 113100 32600 113200 32700
rect 113100 32700 113200 32800
rect 113100 32800 113200 32900
rect 113100 32900 113200 33000
rect 113100 33000 113200 33100
rect 113100 33100 113200 33200
rect 113100 33200 113200 33300
rect 113100 33300 113200 33400
rect 113100 33400 113200 33500
rect 113100 33500 113200 33600
rect 113100 33600 113200 33700
rect 113100 33700 113200 33800
rect 113100 33800 113200 33900
rect 113100 33900 113200 34000
rect 113100 34000 113200 34100
rect 113100 34100 113200 34200
rect 113100 34200 113200 34300
rect 113100 34300 113200 34400
rect 113100 34400 113200 34500
rect 113100 34500 113200 34600
rect 113100 34600 113200 34700
rect 113100 34700 113200 34800
rect 113100 36200 113200 36300
rect 113100 36300 113200 36400
rect 113100 36400 113200 36500
rect 113100 36500 113200 36600
rect 113100 36600 113200 36700
rect 113100 36700 113200 36800
rect 113100 36800 113200 36900
rect 113100 36900 113200 37000
rect 113100 37000 113200 37100
rect 113100 37100 113200 37200
rect 113100 37200 113200 37300
rect 113100 37300 113200 37400
rect 113100 37400 113200 37500
rect 113100 37500 113200 37600
rect 113100 37600 113200 37700
rect 113100 37700 113200 37800
rect 113200 32500 113300 32600
rect 113200 32600 113300 32700
rect 113200 32700 113300 32800
rect 113200 32800 113300 32900
rect 113200 32900 113300 33000
rect 113200 33000 113300 33100
rect 113200 33100 113300 33200
rect 113200 33200 113300 33300
rect 113200 33300 113300 33400
rect 113200 33400 113300 33500
rect 113200 33500 113300 33600
rect 113200 33600 113300 33700
rect 113200 33700 113300 33800
rect 113200 33800 113300 33900
rect 113200 33900 113300 34000
rect 113200 34000 113300 34100
rect 113200 34100 113300 34200
rect 113200 34200 113300 34300
rect 113200 34300 113300 34400
rect 113200 34400 113300 34500
rect 113200 34500 113300 34600
rect 113200 34600 113300 34700
rect 113200 36200 113300 36300
rect 113200 36300 113300 36400
rect 113200 36400 113300 36500
rect 113200 36500 113300 36600
rect 113200 36600 113300 36700
rect 113200 36700 113300 36800
rect 113200 36800 113300 36900
rect 113200 36900 113300 37000
rect 113200 37000 113300 37100
rect 113200 37100 113300 37200
rect 113200 37200 113300 37300
rect 113200 37300 113300 37400
rect 113200 37400 113300 37500
rect 113200 37500 113300 37600
rect 113200 37600 113300 37700
rect 113200 37700 113300 37800
rect 113300 32300 113400 32400
rect 113300 32400 113400 32500
rect 113300 32500 113400 32600
rect 113300 32600 113400 32700
rect 113300 32700 113400 32800
rect 113300 32800 113400 32900
rect 113300 32900 113400 33000
rect 113300 33000 113400 33100
rect 113300 33100 113400 33200
rect 113300 33200 113400 33300
rect 113300 33300 113400 33400
rect 113300 33400 113400 33500
rect 113300 33500 113400 33600
rect 113300 33600 113400 33700
rect 113300 33700 113400 33800
rect 113300 33800 113400 33900
rect 113300 33900 113400 34000
rect 113300 34000 113400 34100
rect 113300 34100 113400 34200
rect 113300 34200 113400 34300
rect 113300 34300 113400 34400
rect 113300 34400 113400 34500
rect 113300 34500 113400 34600
rect 113300 34600 113400 34700
rect 113300 36200 113400 36300
rect 113300 36300 113400 36400
rect 113300 36400 113400 36500
rect 113300 36500 113400 36600
rect 113300 36600 113400 36700
rect 113300 36700 113400 36800
rect 113300 36800 113400 36900
rect 113300 36900 113400 37000
rect 113300 37000 113400 37100
rect 113300 37100 113400 37200
rect 113300 37200 113400 37300
rect 113300 37300 113400 37400
rect 113300 37400 113400 37500
rect 113300 37500 113400 37600
rect 113300 37600 113400 37700
rect 113300 37700 113400 37800
rect 113400 32100 113500 32200
rect 113400 32200 113500 32300
rect 113400 32300 113500 32400
rect 113400 32400 113500 32500
rect 113400 32500 113500 32600
rect 113400 32600 113500 32700
rect 113400 32700 113500 32800
rect 113400 32800 113500 32900
rect 113400 32900 113500 33000
rect 113400 33000 113500 33100
rect 113400 33100 113500 33200
rect 113400 33200 113500 33300
rect 113400 33300 113500 33400
rect 113400 33400 113500 33500
rect 113400 33500 113500 33600
rect 113400 33600 113500 33700
rect 113400 33700 113500 33800
rect 113400 33800 113500 33900
rect 113400 33900 113500 34000
rect 113400 34000 113500 34100
rect 113400 34100 113500 34200
rect 113400 34200 113500 34300
rect 113400 34300 113500 34400
rect 113400 34400 113500 34500
rect 113400 34500 113500 34600
rect 113400 34600 113500 34700
rect 113400 36200 113500 36300
rect 113400 36300 113500 36400
rect 113400 36400 113500 36500
rect 113400 36500 113500 36600
rect 113400 36600 113500 36700
rect 113400 36700 113500 36800
rect 113400 36800 113500 36900
rect 113400 36900 113500 37000
rect 113400 37000 113500 37100
rect 113400 37100 113500 37200
rect 113400 37200 113500 37300
rect 113400 37300 113500 37400
rect 113400 37400 113500 37500
rect 113400 37500 113500 37600
rect 113400 37600 113500 37700
rect 113400 37700 113500 37800
rect 113500 32000 113600 32100
rect 113500 32100 113600 32200
rect 113500 32200 113600 32300
rect 113500 32300 113600 32400
rect 113500 32400 113600 32500
rect 113500 32500 113600 32600
rect 113500 32600 113600 32700
rect 113500 32700 113600 32800
rect 113500 32800 113600 32900
rect 113500 32900 113600 33000
rect 113500 33000 113600 33100
rect 113500 33100 113600 33200
rect 113500 33200 113600 33300
rect 113500 33300 113600 33400
rect 113500 33400 113600 33500
rect 113500 33500 113600 33600
rect 113500 33600 113600 33700
rect 113500 33700 113600 33800
rect 113500 33800 113600 33900
rect 113500 33900 113600 34000
rect 113500 34000 113600 34100
rect 113500 34100 113600 34200
rect 113500 34200 113600 34300
rect 113500 34300 113600 34400
rect 113500 34400 113600 34500
rect 113500 34500 113600 34600
rect 113500 34600 113600 34700
rect 113500 36200 113600 36300
rect 113500 36300 113600 36400
rect 113500 36400 113600 36500
rect 113500 36500 113600 36600
rect 113500 36600 113600 36700
rect 113500 36700 113600 36800
rect 113500 36800 113600 36900
rect 113500 36900 113600 37000
rect 113500 37000 113600 37100
rect 113500 37100 113600 37200
rect 113500 37200 113600 37300
rect 113500 37300 113600 37400
rect 113500 37400 113600 37500
rect 113500 37500 113600 37600
rect 113500 37600 113600 37700
rect 113500 37700 113600 37800
rect 113600 31700 113700 31800
rect 113600 31800 113700 31900
rect 113600 31900 113700 32000
rect 113600 32000 113700 32100
rect 113600 32100 113700 32200
rect 113600 32200 113700 32300
rect 113600 32300 113700 32400
rect 113600 32400 113700 32500
rect 113600 32500 113700 32600
rect 113600 32600 113700 32700
rect 113600 32700 113700 32800
rect 113600 32800 113700 32900
rect 113600 32900 113700 33000
rect 113600 33000 113700 33100
rect 113600 33100 113700 33200
rect 113600 33200 113700 33300
rect 113600 33300 113700 33400
rect 113600 33400 113700 33500
rect 113600 33500 113700 33600
rect 113600 33600 113700 33700
rect 113600 33700 113700 33800
rect 113600 33800 113700 33900
rect 113600 33900 113700 34000
rect 113600 34000 113700 34100
rect 113600 34100 113700 34200
rect 113600 34200 113700 34300
rect 113600 34300 113700 34400
rect 113600 34400 113700 34500
rect 113600 34500 113700 34600
rect 113600 34600 113700 34700
rect 113600 36200 113700 36300
rect 113600 36300 113700 36400
rect 113600 36400 113700 36500
rect 113600 36500 113700 36600
rect 113600 36600 113700 36700
rect 113600 36700 113700 36800
rect 113600 36800 113700 36900
rect 113600 36900 113700 37000
rect 113600 37000 113700 37100
rect 113600 37100 113700 37200
rect 113600 37200 113700 37300
rect 113600 37300 113700 37400
rect 113600 37400 113700 37500
rect 113600 37500 113700 37600
rect 113600 37600 113700 37700
rect 113600 37700 113700 37800
rect 113700 31500 113800 31600
rect 113700 31600 113800 31700
rect 113700 31700 113800 31800
rect 113700 31800 113800 31900
rect 113700 31900 113800 32000
rect 113700 32000 113800 32100
rect 113700 32100 113800 32200
rect 113700 32200 113800 32300
rect 113700 32300 113800 32400
rect 113700 32400 113800 32500
rect 113700 32500 113800 32600
rect 113700 32600 113800 32700
rect 113700 32700 113800 32800
rect 113700 32800 113800 32900
rect 113700 32900 113800 33000
rect 113700 33000 113800 33100
rect 113700 33100 113800 33200
rect 113700 33200 113800 33300
rect 113700 33300 113800 33400
rect 113700 33400 113800 33500
rect 113700 33500 113800 33600
rect 113700 33600 113800 33700
rect 113700 33700 113800 33800
rect 113700 33800 113800 33900
rect 113700 33900 113800 34000
rect 113700 34000 113800 34100
rect 113700 34100 113800 34200
rect 113700 34200 113800 34300
rect 113700 34300 113800 34400
rect 113700 34400 113800 34500
rect 113700 34500 113800 34600
rect 113700 34600 113800 34700
rect 113700 36100 113800 36200
rect 113700 36200 113800 36300
rect 113700 36300 113800 36400
rect 113700 36400 113800 36500
rect 113700 36500 113800 36600
rect 113700 36600 113800 36700
rect 113700 36700 113800 36800
rect 113700 36800 113800 36900
rect 113700 36900 113800 37000
rect 113700 37000 113800 37100
rect 113700 37100 113800 37200
rect 113700 37200 113800 37300
rect 113700 37300 113800 37400
rect 113700 37400 113800 37500
rect 113700 37500 113800 37600
rect 113700 37600 113800 37700
rect 113700 37700 113800 37800
rect 113800 31300 113900 31400
rect 113800 31400 113900 31500
rect 113800 31500 113900 31600
rect 113800 31600 113900 31700
rect 113800 31700 113900 31800
rect 113800 31800 113900 31900
rect 113800 31900 113900 32000
rect 113800 32000 113900 32100
rect 113800 32100 113900 32200
rect 113800 32200 113900 32300
rect 113800 32300 113900 32400
rect 113800 32400 113900 32500
rect 113800 32500 113900 32600
rect 113800 32600 113900 32700
rect 113800 32700 113900 32800
rect 113800 32800 113900 32900
rect 113800 32900 113900 33000
rect 113800 33000 113900 33100
rect 113800 33100 113900 33200
rect 113800 33200 113900 33300
rect 113800 33300 113900 33400
rect 113800 33400 113900 33500
rect 113800 33500 113900 33600
rect 113800 33600 113900 33700
rect 113800 33700 113900 33800
rect 113800 33800 113900 33900
rect 113800 33900 113900 34000
rect 113800 34000 113900 34100
rect 113800 34100 113900 34200
rect 113800 34200 113900 34300
rect 113800 34300 113900 34400
rect 113800 34400 113900 34500
rect 113800 34500 113900 34600
rect 113800 34600 113900 34700
rect 113800 36000 113900 36100
rect 113800 36100 113900 36200
rect 113800 36200 113900 36300
rect 113800 36300 113900 36400
rect 113800 36400 113900 36500
rect 113800 36500 113900 36600
rect 113800 36600 113900 36700
rect 113800 36700 113900 36800
rect 113800 36800 113900 36900
rect 113800 36900 113900 37000
rect 113800 37000 113900 37100
rect 113800 37100 113900 37200
rect 113800 37200 113900 37300
rect 113800 37300 113900 37400
rect 113800 37400 113900 37500
rect 113800 37500 113900 37600
rect 113800 37600 113900 37700
rect 113800 37700 113900 37800
rect 113900 31000 114000 31100
rect 113900 31100 114000 31200
rect 113900 31200 114000 31300
rect 113900 31300 114000 31400
rect 113900 31400 114000 31500
rect 113900 31500 114000 31600
rect 113900 31600 114000 31700
rect 113900 31700 114000 31800
rect 113900 31800 114000 31900
rect 113900 31900 114000 32000
rect 113900 32000 114000 32100
rect 113900 32100 114000 32200
rect 113900 32200 114000 32300
rect 113900 32300 114000 32400
rect 113900 32400 114000 32500
rect 113900 32500 114000 32600
rect 113900 32600 114000 32700
rect 113900 32700 114000 32800
rect 113900 32800 114000 32900
rect 113900 32900 114000 33000
rect 113900 33000 114000 33100
rect 113900 33100 114000 33200
rect 113900 33200 114000 33300
rect 113900 33300 114000 33400
rect 113900 33400 114000 33500
rect 113900 33500 114000 33600
rect 113900 33600 114000 33700
rect 113900 33700 114000 33800
rect 113900 33800 114000 33900
rect 113900 33900 114000 34000
rect 113900 34000 114000 34100
rect 113900 34100 114000 34200
rect 113900 34200 114000 34300
rect 113900 34300 114000 34400
rect 113900 34400 114000 34500
rect 113900 34500 114000 34600
rect 113900 34600 114000 34700
rect 113900 34700 114000 34800
rect 113900 35800 114000 35900
rect 113900 35900 114000 36000
rect 113900 36000 114000 36100
rect 113900 36100 114000 36200
rect 113900 36200 114000 36300
rect 113900 36300 114000 36400
rect 113900 36400 114000 36500
rect 113900 36500 114000 36600
rect 113900 36600 114000 36700
rect 113900 36700 114000 36800
rect 113900 36800 114000 36900
rect 113900 36900 114000 37000
rect 113900 37000 114000 37100
rect 113900 37100 114000 37200
rect 113900 37200 114000 37300
rect 113900 37300 114000 37400
rect 113900 37400 114000 37500
rect 113900 37500 114000 37600
rect 113900 37600 114000 37700
rect 114000 30800 114100 30900
rect 114000 30900 114100 31000
rect 114000 31000 114100 31100
rect 114000 31100 114100 31200
rect 114000 31200 114100 31300
rect 114000 31300 114100 31400
rect 114000 31400 114100 31500
rect 114000 31500 114100 31600
rect 114000 31600 114100 31700
rect 114000 31700 114100 31800
rect 114000 31800 114100 31900
rect 114000 31900 114100 32000
rect 114000 32000 114100 32100
rect 114000 32100 114100 32200
rect 114000 32200 114100 32300
rect 114000 32300 114100 32400
rect 114000 32400 114100 32500
rect 114000 32500 114100 32600
rect 114000 32600 114100 32700
rect 114000 32700 114100 32800
rect 114000 32800 114100 32900
rect 114000 32900 114100 33000
rect 114000 33000 114100 33100
rect 114000 33100 114100 33200
rect 114000 33200 114100 33300
rect 114000 33300 114100 33400
rect 114000 33400 114100 33500
rect 114000 33500 114100 33600
rect 114000 33600 114100 33700
rect 114000 33700 114100 33800
rect 114000 33800 114100 33900
rect 114000 33900 114100 34000
rect 114000 34000 114100 34100
rect 114000 34100 114100 34200
rect 114000 34200 114100 34300
rect 114000 34300 114100 34400
rect 114000 34400 114100 34500
rect 114000 34500 114100 34600
rect 114000 34600 114100 34700
rect 114000 34700 114100 34800
rect 114000 34800 114100 34900
rect 114000 34900 114100 35000
rect 114000 35000 114100 35100
rect 114000 35300 114100 35400
rect 114000 35500 114100 35600
rect 114000 35600 114100 35700
rect 114000 35700 114100 35800
rect 114000 35800 114100 35900
rect 114000 35900 114100 36000
rect 114000 36000 114100 36100
rect 114000 36100 114100 36200
rect 114000 36200 114100 36300
rect 114000 36300 114100 36400
rect 114000 36400 114100 36500
rect 114000 36500 114100 36600
rect 114000 36600 114100 36700
rect 114000 36700 114100 36800
rect 114000 36800 114100 36900
rect 114000 36900 114100 37000
rect 114000 37000 114100 37100
rect 114000 37100 114100 37200
rect 114000 37200 114100 37300
rect 114000 37300 114100 37400
rect 114000 37400 114100 37500
rect 114000 37500 114100 37600
rect 114000 37600 114100 37700
rect 114100 30500 114200 30600
rect 114100 30600 114200 30700
rect 114100 30700 114200 30800
rect 114100 30800 114200 30900
rect 114100 30900 114200 31000
rect 114100 31000 114200 31100
rect 114100 31100 114200 31200
rect 114100 31200 114200 31300
rect 114100 31300 114200 31400
rect 114100 31400 114200 31500
rect 114100 31500 114200 31600
rect 114100 31600 114200 31700
rect 114100 31700 114200 31800
rect 114100 31800 114200 31900
rect 114100 31900 114200 32000
rect 114100 32000 114200 32100
rect 114100 32100 114200 32200
rect 114100 32200 114200 32300
rect 114100 32300 114200 32400
rect 114100 32400 114200 32500
rect 114100 32500 114200 32600
rect 114100 32600 114200 32700
rect 114100 32700 114200 32800
rect 114100 32800 114200 32900
rect 114100 32900 114200 33000
rect 114100 33000 114200 33100
rect 114100 33100 114200 33200
rect 114100 33200 114200 33300
rect 114100 33300 114200 33400
rect 114100 33400 114200 33500
rect 114100 33500 114200 33600
rect 114100 33600 114200 33700
rect 114100 33700 114200 33800
rect 114100 33800 114200 33900
rect 114100 33900 114200 34000
rect 114100 34000 114200 34100
rect 114100 34100 114200 34200
rect 114100 34200 114200 34300
rect 114100 34300 114200 34400
rect 114100 34400 114200 34500
rect 114100 34500 114200 34600
rect 114100 34600 114200 34700
rect 114100 34700 114200 34800
rect 114100 34800 114200 34900
rect 114100 34900 114200 35000
rect 114100 35000 114200 35100
rect 114100 35100 114200 35200
rect 114100 35200 114200 35300
rect 114100 35300 114200 35400
rect 114100 35400 114200 35500
rect 114100 35500 114200 35600
rect 114100 35600 114200 35700
rect 114100 35700 114200 35800
rect 114100 35800 114200 35900
rect 114100 35900 114200 36000
rect 114100 36000 114200 36100
rect 114100 36100 114200 36200
rect 114100 36200 114200 36300
rect 114100 36300 114200 36400
rect 114100 36400 114200 36500
rect 114100 36500 114200 36600
rect 114100 36600 114200 36700
rect 114100 36700 114200 36800
rect 114100 36800 114200 36900
rect 114100 36900 114200 37000
rect 114100 37000 114200 37100
rect 114100 37100 114200 37200
rect 114100 37200 114200 37300
rect 114100 37300 114200 37400
rect 114100 37400 114200 37500
rect 114100 37500 114200 37600
rect 114100 37600 114200 37700
rect 114200 30200 114300 30300
rect 114200 30300 114300 30400
rect 114200 30400 114300 30500
rect 114200 30500 114300 30600
rect 114200 30600 114300 30700
rect 114200 30700 114300 30800
rect 114200 30800 114300 30900
rect 114200 30900 114300 31000
rect 114200 31000 114300 31100
rect 114200 31100 114300 31200
rect 114200 31200 114300 31300
rect 114200 31300 114300 31400
rect 114200 31400 114300 31500
rect 114200 31500 114300 31600
rect 114200 31600 114300 31700
rect 114200 31700 114300 31800
rect 114200 31800 114300 31900
rect 114200 31900 114300 32000
rect 114200 32000 114300 32100
rect 114200 32100 114300 32200
rect 114200 32200 114300 32300
rect 114200 32300 114300 32400
rect 114200 32400 114300 32500
rect 114200 32500 114300 32600
rect 114200 32600 114300 32700
rect 114200 32700 114300 32800
rect 114200 32800 114300 32900
rect 114200 32900 114300 33000
rect 114200 33000 114300 33100
rect 114200 33100 114300 33200
rect 114200 33200 114300 33300
rect 114200 33300 114300 33400
rect 114200 33400 114300 33500
rect 114200 33500 114300 33600
rect 114200 33600 114300 33700
rect 114200 33700 114300 33800
rect 114200 33800 114300 33900
rect 114200 33900 114300 34000
rect 114200 34000 114300 34100
rect 114200 34100 114300 34200
rect 114200 34200 114300 34300
rect 114200 34300 114300 34400
rect 114200 34400 114300 34500
rect 114200 34500 114300 34600
rect 114200 34600 114300 34700
rect 114200 34700 114300 34800
rect 114200 34800 114300 34900
rect 114200 34900 114300 35000
rect 114200 35000 114300 35100
rect 114200 35100 114300 35200
rect 114200 35200 114300 35300
rect 114200 35300 114300 35400
rect 114200 35400 114300 35500
rect 114200 35500 114300 35600
rect 114200 35600 114300 35700
rect 114200 35700 114300 35800
rect 114200 35800 114300 35900
rect 114200 35900 114300 36000
rect 114200 36000 114300 36100
rect 114200 36100 114300 36200
rect 114200 36200 114300 36300
rect 114200 36300 114300 36400
rect 114200 36400 114300 36500
rect 114200 36500 114300 36600
rect 114200 36600 114300 36700
rect 114200 36700 114300 36800
rect 114200 36800 114300 36900
rect 114200 36900 114300 37000
rect 114200 37000 114300 37100
rect 114200 37100 114300 37200
rect 114200 37200 114300 37300
rect 114200 37300 114300 37400
rect 114200 37400 114300 37500
rect 114200 37500 114300 37600
rect 114300 29900 114400 30000
rect 114300 30000 114400 30100
rect 114300 30100 114400 30200
rect 114300 30200 114400 30300
rect 114300 30300 114400 30400
rect 114300 30400 114400 30500
rect 114300 30500 114400 30600
rect 114300 30600 114400 30700
rect 114300 30700 114400 30800
rect 114300 30800 114400 30900
rect 114300 30900 114400 31000
rect 114300 31000 114400 31100
rect 114300 31100 114400 31200
rect 114300 31200 114400 31300
rect 114300 31300 114400 31400
rect 114300 31400 114400 31500
rect 114300 31500 114400 31600
rect 114300 31600 114400 31700
rect 114300 31700 114400 31800
rect 114300 31800 114400 31900
rect 114300 31900 114400 32000
rect 114300 32000 114400 32100
rect 114300 32100 114400 32200
rect 114300 32200 114400 32300
rect 114300 32300 114400 32400
rect 114300 32400 114400 32500
rect 114300 32500 114400 32600
rect 114300 32600 114400 32700
rect 114300 32700 114400 32800
rect 114300 32800 114400 32900
rect 114300 32900 114400 33000
rect 114300 33000 114400 33100
rect 114300 33100 114400 33200
rect 114300 33200 114400 33300
rect 114300 33300 114400 33400
rect 114300 33400 114400 33500
rect 114300 33500 114400 33600
rect 114300 33600 114400 33700
rect 114300 33700 114400 33800
rect 114300 33800 114400 33900
rect 114300 33900 114400 34000
rect 114300 34000 114400 34100
rect 114300 34100 114400 34200
rect 114300 34200 114400 34300
rect 114300 34300 114400 34400
rect 114300 34400 114400 34500
rect 114300 34500 114400 34600
rect 114300 34600 114400 34700
rect 114300 34700 114400 34800
rect 114300 34800 114400 34900
rect 114300 34900 114400 35000
rect 114300 35000 114400 35100
rect 114300 35100 114400 35200
rect 114300 35200 114400 35300
rect 114300 35300 114400 35400
rect 114300 35400 114400 35500
rect 114300 35500 114400 35600
rect 114300 35600 114400 35700
rect 114300 35700 114400 35800
rect 114300 35800 114400 35900
rect 114300 35900 114400 36000
rect 114300 36000 114400 36100
rect 114300 36100 114400 36200
rect 114300 36200 114400 36300
rect 114300 36300 114400 36400
rect 114300 36400 114400 36500
rect 114300 36500 114400 36600
rect 114300 36600 114400 36700
rect 114300 36700 114400 36800
rect 114300 36800 114400 36900
rect 114300 36900 114400 37000
rect 114300 37000 114400 37100
rect 114300 37100 114400 37200
rect 114300 37200 114400 37300
rect 114300 37300 114400 37400
rect 114300 37400 114400 37500
rect 114300 37500 114400 37600
rect 114400 29600 114500 29700
rect 114400 29700 114500 29800
rect 114400 29800 114500 29900
rect 114400 29900 114500 30000
rect 114400 30000 114500 30100
rect 114400 30100 114500 30200
rect 114400 30200 114500 30300
rect 114400 30300 114500 30400
rect 114400 30400 114500 30500
rect 114400 30500 114500 30600
rect 114400 30600 114500 30700
rect 114400 30700 114500 30800
rect 114400 30800 114500 30900
rect 114400 30900 114500 31000
rect 114400 31000 114500 31100
rect 114400 31100 114500 31200
rect 114400 31200 114500 31300
rect 114400 31300 114500 31400
rect 114400 31400 114500 31500
rect 114400 31500 114500 31600
rect 114400 31600 114500 31700
rect 114400 31700 114500 31800
rect 114400 31800 114500 31900
rect 114400 31900 114500 32000
rect 114400 32000 114500 32100
rect 114400 32100 114500 32200
rect 114400 32200 114500 32300
rect 114400 32300 114500 32400
rect 114400 32400 114500 32500
rect 114400 32500 114500 32600
rect 114400 32600 114500 32700
rect 114400 32700 114500 32800
rect 114400 32800 114500 32900
rect 114400 32900 114500 33000
rect 114400 33000 114500 33100
rect 114400 33100 114500 33200
rect 114400 33200 114500 33300
rect 114400 33300 114500 33400
rect 114400 33400 114500 33500
rect 114400 33500 114500 33600
rect 114400 33600 114500 33700
rect 114400 33700 114500 33800
rect 114400 33800 114500 33900
rect 114400 33900 114500 34000
rect 114400 34000 114500 34100
rect 114400 34100 114500 34200
rect 114400 34200 114500 34300
rect 114400 34300 114500 34400
rect 114400 34400 114500 34500
rect 114400 34500 114500 34600
rect 114400 34600 114500 34700
rect 114400 34700 114500 34800
rect 114400 34800 114500 34900
rect 114400 34900 114500 35000
rect 114400 35000 114500 35100
rect 114400 35100 114500 35200
rect 114400 35200 114500 35300
rect 114400 35300 114500 35400
rect 114400 35400 114500 35500
rect 114400 35500 114500 35600
rect 114400 35600 114500 35700
rect 114400 35700 114500 35800
rect 114400 35800 114500 35900
rect 114400 35900 114500 36000
rect 114400 36000 114500 36100
rect 114400 36100 114500 36200
rect 114400 36200 114500 36300
rect 114400 36300 114500 36400
rect 114400 36400 114500 36500
rect 114400 36500 114500 36600
rect 114400 36600 114500 36700
rect 114400 36700 114500 36800
rect 114400 36800 114500 36900
rect 114400 36900 114500 37000
rect 114400 37000 114500 37100
rect 114400 37100 114500 37200
rect 114400 37200 114500 37300
rect 114400 37300 114500 37400
rect 114400 37400 114500 37500
rect 114400 37500 114500 37600
rect 114500 29300 114600 29400
rect 114500 29400 114600 29500
rect 114500 29500 114600 29600
rect 114500 29600 114600 29700
rect 114500 29700 114600 29800
rect 114500 29800 114600 29900
rect 114500 29900 114600 30000
rect 114500 30000 114600 30100
rect 114500 30100 114600 30200
rect 114500 30200 114600 30300
rect 114500 30300 114600 30400
rect 114500 30400 114600 30500
rect 114500 30500 114600 30600
rect 114500 30600 114600 30700
rect 114500 30700 114600 30800
rect 114500 30800 114600 30900
rect 114500 30900 114600 31000
rect 114500 31000 114600 31100
rect 114500 31100 114600 31200
rect 114500 31200 114600 31300
rect 114500 31300 114600 31400
rect 114500 31400 114600 31500
rect 114500 31500 114600 31600
rect 114500 31600 114600 31700
rect 114500 31700 114600 31800
rect 114500 31800 114600 31900
rect 114500 31900 114600 32000
rect 114500 32000 114600 32100
rect 114500 32100 114600 32200
rect 114500 32200 114600 32300
rect 114500 32300 114600 32400
rect 114500 32400 114600 32500
rect 114500 32500 114600 32600
rect 114500 32600 114600 32700
rect 114500 32700 114600 32800
rect 114500 32800 114600 32900
rect 114500 32900 114600 33000
rect 114500 33000 114600 33100
rect 114500 33100 114600 33200
rect 114500 33200 114600 33300
rect 114500 33300 114600 33400
rect 114500 33400 114600 33500
rect 114500 33500 114600 33600
rect 114500 33600 114600 33700
rect 114500 33700 114600 33800
rect 114500 33800 114600 33900
rect 114500 33900 114600 34000
rect 114500 34000 114600 34100
rect 114500 34100 114600 34200
rect 114500 34200 114600 34300
rect 114500 34300 114600 34400
rect 114500 34400 114600 34500
rect 114500 34500 114600 34600
rect 114500 34600 114600 34700
rect 114500 34700 114600 34800
rect 114500 34800 114600 34900
rect 114500 34900 114600 35000
rect 114500 35000 114600 35100
rect 114500 35100 114600 35200
rect 114500 35200 114600 35300
rect 114500 35300 114600 35400
rect 114500 35400 114600 35500
rect 114500 35500 114600 35600
rect 114500 35600 114600 35700
rect 114500 35700 114600 35800
rect 114500 35800 114600 35900
rect 114500 35900 114600 36000
rect 114500 36000 114600 36100
rect 114500 36100 114600 36200
rect 114500 36200 114600 36300
rect 114500 36300 114600 36400
rect 114500 36400 114600 36500
rect 114500 36500 114600 36600
rect 114500 36600 114600 36700
rect 114500 36700 114600 36800
rect 114500 36800 114600 36900
rect 114500 36900 114600 37000
rect 114500 37000 114600 37100
rect 114500 37100 114600 37200
rect 114500 37200 114600 37300
rect 114500 37300 114600 37400
rect 114500 37400 114600 37500
rect 114600 29100 114700 29200
rect 114600 29200 114700 29300
rect 114600 29300 114700 29400
rect 114600 29400 114700 29500
rect 114600 29500 114700 29600
rect 114600 29600 114700 29700
rect 114600 29700 114700 29800
rect 114600 29800 114700 29900
rect 114600 29900 114700 30000
rect 114600 30000 114700 30100
rect 114600 30100 114700 30200
rect 114600 30200 114700 30300
rect 114600 30300 114700 30400
rect 114600 30400 114700 30500
rect 114600 30500 114700 30600
rect 114600 30600 114700 30700
rect 114600 30700 114700 30800
rect 114600 30800 114700 30900
rect 114600 30900 114700 31000
rect 114600 31000 114700 31100
rect 114600 31100 114700 31200
rect 114600 31200 114700 31300
rect 114600 31300 114700 31400
rect 114600 31400 114700 31500
rect 114600 31500 114700 31600
rect 114600 31600 114700 31700
rect 114600 31700 114700 31800
rect 114600 31800 114700 31900
rect 114600 31900 114700 32000
rect 114600 32000 114700 32100
rect 114600 32100 114700 32200
rect 114600 32200 114700 32300
rect 114600 32300 114700 32400
rect 114600 32400 114700 32500
rect 114600 32500 114700 32600
rect 114600 32600 114700 32700
rect 114600 32700 114700 32800
rect 114600 32800 114700 32900
rect 114600 32900 114700 33000
rect 114600 33000 114700 33100
rect 114600 33100 114700 33200
rect 114600 33200 114700 33300
rect 114600 33300 114700 33400
rect 114600 33400 114700 33500
rect 114600 33500 114700 33600
rect 114600 33600 114700 33700
rect 114600 33700 114700 33800
rect 114600 33800 114700 33900
rect 114600 33900 114700 34000
rect 114600 34000 114700 34100
rect 114600 34100 114700 34200
rect 114600 34200 114700 34300
rect 114600 34300 114700 34400
rect 114600 34400 114700 34500
rect 114600 34500 114700 34600
rect 114600 34600 114700 34700
rect 114600 34700 114700 34800
rect 114600 34800 114700 34900
rect 114600 34900 114700 35000
rect 114600 35000 114700 35100
rect 114600 35100 114700 35200
rect 114600 35200 114700 35300
rect 114600 35300 114700 35400
rect 114600 35400 114700 35500
rect 114600 35500 114700 35600
rect 114600 35600 114700 35700
rect 114600 35700 114700 35800
rect 114600 35800 114700 35900
rect 114600 35900 114700 36000
rect 114600 36000 114700 36100
rect 114600 36100 114700 36200
rect 114600 36200 114700 36300
rect 114600 36300 114700 36400
rect 114600 36400 114700 36500
rect 114600 36500 114700 36600
rect 114600 36600 114700 36700
rect 114600 36700 114700 36800
rect 114600 36800 114700 36900
rect 114600 36900 114700 37000
rect 114600 37000 114700 37100
rect 114600 37100 114700 37200
rect 114600 37200 114700 37300
rect 114600 37300 114700 37400
rect 114700 22700 114800 22800
rect 114700 22800 114800 22900
rect 114700 22900 114800 23000
rect 114700 23000 114800 23100
rect 114700 23100 114800 23200
rect 114700 23200 114800 23300
rect 114700 23300 114800 23400
rect 114700 23400 114800 23500
rect 114700 23500 114800 23600
rect 114700 23600 114800 23700
rect 114700 23700 114800 23800
rect 114700 28800 114800 28900
rect 114700 28900 114800 29000
rect 114700 29000 114800 29100
rect 114700 29100 114800 29200
rect 114700 29200 114800 29300
rect 114700 29300 114800 29400
rect 114700 29400 114800 29500
rect 114700 29500 114800 29600
rect 114700 29600 114800 29700
rect 114700 29700 114800 29800
rect 114700 29800 114800 29900
rect 114700 29900 114800 30000
rect 114700 30000 114800 30100
rect 114700 30100 114800 30200
rect 114700 30200 114800 30300
rect 114700 30300 114800 30400
rect 114700 30400 114800 30500
rect 114700 30500 114800 30600
rect 114700 30600 114800 30700
rect 114700 30700 114800 30800
rect 114700 30800 114800 30900
rect 114700 30900 114800 31000
rect 114700 31000 114800 31100
rect 114700 31100 114800 31200
rect 114700 31200 114800 31300
rect 114700 31300 114800 31400
rect 114700 31400 114800 31500
rect 114700 31500 114800 31600
rect 114700 31600 114800 31700
rect 114700 31700 114800 31800
rect 114700 31800 114800 31900
rect 114700 31900 114800 32000
rect 114700 32000 114800 32100
rect 114700 32100 114800 32200
rect 114700 32200 114800 32300
rect 114700 32300 114800 32400
rect 114700 32400 114800 32500
rect 114700 32500 114800 32600
rect 114700 32600 114800 32700
rect 114700 32700 114800 32800
rect 114700 32800 114800 32900
rect 114700 32900 114800 33000
rect 114700 33000 114800 33100
rect 114700 33100 114800 33200
rect 114700 33200 114800 33300
rect 114700 33300 114800 33400
rect 114700 33400 114800 33500
rect 114700 33500 114800 33600
rect 114700 33600 114800 33700
rect 114700 33700 114800 33800
rect 114700 33800 114800 33900
rect 114700 33900 114800 34000
rect 114700 34000 114800 34100
rect 114700 34100 114800 34200
rect 114700 34200 114800 34300
rect 114700 34300 114800 34400
rect 114700 34400 114800 34500
rect 114700 34500 114800 34600
rect 114700 34600 114800 34700
rect 114700 34700 114800 34800
rect 114700 34800 114800 34900
rect 114700 34900 114800 35000
rect 114700 35000 114800 35100
rect 114700 35100 114800 35200
rect 114700 35200 114800 35300
rect 114700 35300 114800 35400
rect 114700 35400 114800 35500
rect 114700 35500 114800 35600
rect 114700 35600 114800 35700
rect 114700 35700 114800 35800
rect 114700 35800 114800 35900
rect 114700 35900 114800 36000
rect 114700 36000 114800 36100
rect 114700 36100 114800 36200
rect 114700 36200 114800 36300
rect 114700 36300 114800 36400
rect 114700 36400 114800 36500
rect 114700 36500 114800 36600
rect 114700 36600 114800 36700
rect 114700 36700 114800 36800
rect 114700 36800 114800 36900
rect 114700 36900 114800 37000
rect 114700 37000 114800 37100
rect 114700 37100 114800 37200
rect 114700 37200 114800 37300
rect 114700 37300 114800 37400
rect 114800 22300 114900 22400
rect 114800 22400 114900 22500
rect 114800 22500 114900 22600
rect 114800 22600 114900 22700
rect 114800 22700 114900 22800
rect 114800 22800 114900 22900
rect 114800 22900 114900 23000
rect 114800 23000 114900 23100
rect 114800 23100 114900 23200
rect 114800 23200 114900 23300
rect 114800 23300 114900 23400
rect 114800 23400 114900 23500
rect 114800 23500 114900 23600
rect 114800 23600 114900 23700
rect 114800 23700 114900 23800
rect 114800 23800 114900 23900
rect 114800 23900 114900 24000
rect 114800 24000 114900 24100
rect 114800 28500 114900 28600
rect 114800 28600 114900 28700
rect 114800 28700 114900 28800
rect 114800 28800 114900 28900
rect 114800 28900 114900 29000
rect 114800 29000 114900 29100
rect 114800 29100 114900 29200
rect 114800 29200 114900 29300
rect 114800 29300 114900 29400
rect 114800 29400 114900 29500
rect 114800 29500 114900 29600
rect 114800 29600 114900 29700
rect 114800 29700 114900 29800
rect 114800 29800 114900 29900
rect 114800 29900 114900 30000
rect 114800 30000 114900 30100
rect 114800 30100 114900 30200
rect 114800 30200 114900 30300
rect 114800 30300 114900 30400
rect 114800 30400 114900 30500
rect 114800 30500 114900 30600
rect 114800 30600 114900 30700
rect 114800 30700 114900 30800
rect 114800 30800 114900 30900
rect 114800 30900 114900 31000
rect 114800 31000 114900 31100
rect 114800 31100 114900 31200
rect 114800 31200 114900 31300
rect 114800 31300 114900 31400
rect 114800 31400 114900 31500
rect 114800 31500 114900 31600
rect 114800 31600 114900 31700
rect 114800 31700 114900 31800
rect 114800 31800 114900 31900
rect 114800 31900 114900 32000
rect 114800 32000 114900 32100
rect 114800 32100 114900 32200
rect 114800 32200 114900 32300
rect 114800 32300 114900 32400
rect 114800 32400 114900 32500
rect 114800 32500 114900 32600
rect 114800 32600 114900 32700
rect 114800 32700 114900 32800
rect 114800 32800 114900 32900
rect 114800 32900 114900 33000
rect 114800 33000 114900 33100
rect 114800 33100 114900 33200
rect 114800 33200 114900 33300
rect 114800 33300 114900 33400
rect 114800 33400 114900 33500
rect 114800 33500 114900 33600
rect 114800 33600 114900 33700
rect 114800 33700 114900 33800
rect 114800 33800 114900 33900
rect 114800 33900 114900 34000
rect 114800 34000 114900 34100
rect 114800 34100 114900 34200
rect 114800 34200 114900 34300
rect 114800 34300 114900 34400
rect 114800 34400 114900 34500
rect 114800 34500 114900 34600
rect 114800 34600 114900 34700
rect 114800 34700 114900 34800
rect 114800 34800 114900 34900
rect 114800 34900 114900 35000
rect 114800 35000 114900 35100
rect 114800 35100 114900 35200
rect 114800 35200 114900 35300
rect 114800 35300 114900 35400
rect 114800 35400 114900 35500
rect 114800 35500 114900 35600
rect 114800 35600 114900 35700
rect 114800 35700 114900 35800
rect 114800 35800 114900 35900
rect 114800 35900 114900 36000
rect 114800 36000 114900 36100
rect 114800 36100 114900 36200
rect 114800 36200 114900 36300
rect 114800 36300 114900 36400
rect 114800 36400 114900 36500
rect 114800 36500 114900 36600
rect 114800 36600 114900 36700
rect 114800 36700 114900 36800
rect 114800 36800 114900 36900
rect 114800 36900 114900 37000
rect 114800 37000 114900 37100
rect 114800 37100 114900 37200
rect 114800 37200 114900 37300
rect 114900 22100 115000 22200
rect 114900 22200 115000 22300
rect 114900 22300 115000 22400
rect 114900 22400 115000 22500
rect 114900 22500 115000 22600
rect 114900 22600 115000 22700
rect 114900 22700 115000 22800
rect 114900 22800 115000 22900
rect 114900 22900 115000 23000
rect 114900 23000 115000 23100
rect 114900 23100 115000 23200
rect 114900 23200 115000 23300
rect 114900 23300 115000 23400
rect 114900 23400 115000 23500
rect 114900 23500 115000 23600
rect 114900 23600 115000 23700
rect 114900 23700 115000 23800
rect 114900 23800 115000 23900
rect 114900 23900 115000 24000
rect 114900 24000 115000 24100
rect 114900 24100 115000 24200
rect 114900 24200 115000 24300
rect 114900 24300 115000 24400
rect 114900 28200 115000 28300
rect 114900 28300 115000 28400
rect 114900 28400 115000 28500
rect 114900 28500 115000 28600
rect 114900 28600 115000 28700
rect 114900 28700 115000 28800
rect 114900 28800 115000 28900
rect 114900 28900 115000 29000
rect 114900 29000 115000 29100
rect 114900 29100 115000 29200
rect 114900 29200 115000 29300
rect 114900 29300 115000 29400
rect 114900 29400 115000 29500
rect 114900 29500 115000 29600
rect 114900 29600 115000 29700
rect 114900 29700 115000 29800
rect 114900 29800 115000 29900
rect 114900 29900 115000 30000
rect 114900 30000 115000 30100
rect 114900 30100 115000 30200
rect 114900 30200 115000 30300
rect 114900 30300 115000 30400
rect 114900 30400 115000 30500
rect 114900 30500 115000 30600
rect 114900 30600 115000 30700
rect 114900 30700 115000 30800
rect 114900 30800 115000 30900
rect 114900 30900 115000 31000
rect 114900 31000 115000 31100
rect 114900 31100 115000 31200
rect 114900 31200 115000 31300
rect 114900 31300 115000 31400
rect 114900 31400 115000 31500
rect 114900 31500 115000 31600
rect 114900 31600 115000 31700
rect 114900 31700 115000 31800
rect 114900 31800 115000 31900
rect 114900 31900 115000 32000
rect 114900 32000 115000 32100
rect 114900 32100 115000 32200
rect 114900 32200 115000 32300
rect 114900 32300 115000 32400
rect 114900 32400 115000 32500
rect 114900 32500 115000 32600
rect 114900 32600 115000 32700
rect 114900 32700 115000 32800
rect 114900 32800 115000 32900
rect 114900 32900 115000 33000
rect 114900 33000 115000 33100
rect 114900 33100 115000 33200
rect 114900 33200 115000 33300
rect 114900 33300 115000 33400
rect 114900 33400 115000 33500
rect 114900 33500 115000 33600
rect 114900 33600 115000 33700
rect 114900 33700 115000 33800
rect 114900 33800 115000 33900
rect 114900 33900 115000 34000
rect 114900 34000 115000 34100
rect 114900 34100 115000 34200
rect 114900 34200 115000 34300
rect 114900 34300 115000 34400
rect 114900 34400 115000 34500
rect 114900 34500 115000 34600
rect 114900 34600 115000 34700
rect 114900 34700 115000 34800
rect 114900 34800 115000 34900
rect 114900 34900 115000 35000
rect 114900 35000 115000 35100
rect 114900 35100 115000 35200
rect 114900 35200 115000 35300
rect 114900 35300 115000 35400
rect 114900 35400 115000 35500
rect 114900 35500 115000 35600
rect 114900 35600 115000 35700
rect 114900 35700 115000 35800
rect 114900 35800 115000 35900
rect 114900 35900 115000 36000
rect 114900 36000 115000 36100
rect 114900 36100 115000 36200
rect 114900 36200 115000 36300
rect 114900 36300 115000 36400
rect 114900 36400 115000 36500
rect 114900 36500 115000 36600
rect 114900 36600 115000 36700
rect 114900 36700 115000 36800
rect 114900 36800 115000 36900
rect 114900 36900 115000 37000
rect 114900 37000 115000 37100
rect 114900 37100 115000 37200
rect 115000 21900 115100 22000
rect 115000 22000 115100 22100
rect 115000 22100 115100 22200
rect 115000 22200 115100 22300
rect 115000 22300 115100 22400
rect 115000 22400 115100 22500
rect 115000 22500 115100 22600
rect 115000 22600 115100 22700
rect 115000 22700 115100 22800
rect 115000 22800 115100 22900
rect 115000 22900 115100 23000
rect 115000 23000 115100 23100
rect 115000 23100 115100 23200
rect 115000 23200 115100 23300
rect 115000 23300 115100 23400
rect 115000 23400 115100 23500
rect 115000 23500 115100 23600
rect 115000 23600 115100 23700
rect 115000 23700 115100 23800
rect 115000 23800 115100 23900
rect 115000 23900 115100 24000
rect 115000 24000 115100 24100
rect 115000 24100 115100 24200
rect 115000 24200 115100 24300
rect 115000 24300 115100 24400
rect 115000 24400 115100 24500
rect 115000 24500 115100 24600
rect 115000 27900 115100 28000
rect 115000 28000 115100 28100
rect 115000 28100 115100 28200
rect 115000 28200 115100 28300
rect 115000 28300 115100 28400
rect 115000 28400 115100 28500
rect 115000 28500 115100 28600
rect 115000 28600 115100 28700
rect 115000 28700 115100 28800
rect 115000 28800 115100 28900
rect 115000 28900 115100 29000
rect 115000 29000 115100 29100
rect 115000 29100 115100 29200
rect 115000 29200 115100 29300
rect 115000 29300 115100 29400
rect 115000 29400 115100 29500
rect 115000 29500 115100 29600
rect 115000 29600 115100 29700
rect 115000 29700 115100 29800
rect 115000 29800 115100 29900
rect 115000 29900 115100 30000
rect 115000 30000 115100 30100
rect 115000 30100 115100 30200
rect 115000 30200 115100 30300
rect 115000 30300 115100 30400
rect 115000 30400 115100 30500
rect 115000 30500 115100 30600
rect 115000 30600 115100 30700
rect 115000 30700 115100 30800
rect 115000 30800 115100 30900
rect 115000 30900 115100 31000
rect 115000 31000 115100 31100
rect 115000 31100 115100 31200
rect 115000 31200 115100 31300
rect 115000 31300 115100 31400
rect 115000 31400 115100 31500
rect 115000 31500 115100 31600
rect 115000 31600 115100 31700
rect 115000 31700 115100 31800
rect 115000 31800 115100 31900
rect 115000 31900 115100 32000
rect 115000 32000 115100 32100
rect 115000 32100 115100 32200
rect 115000 32200 115100 32300
rect 115000 32300 115100 32400
rect 115000 32400 115100 32500
rect 115000 32500 115100 32600
rect 115000 32600 115100 32700
rect 115000 32700 115100 32800
rect 115000 32800 115100 32900
rect 115000 32900 115100 33000
rect 115000 33000 115100 33100
rect 115000 33100 115100 33200
rect 115000 33200 115100 33300
rect 115000 33300 115100 33400
rect 115000 33400 115100 33500
rect 115000 33500 115100 33600
rect 115000 33600 115100 33700
rect 115000 33700 115100 33800
rect 115000 33800 115100 33900
rect 115000 33900 115100 34000
rect 115000 34000 115100 34100
rect 115000 34100 115100 34200
rect 115000 34200 115100 34300
rect 115000 34300 115100 34400
rect 115000 34400 115100 34500
rect 115000 34500 115100 34600
rect 115000 34600 115100 34700
rect 115000 34700 115100 34800
rect 115000 34800 115100 34900
rect 115000 34900 115100 35000
rect 115000 35000 115100 35100
rect 115000 35100 115100 35200
rect 115000 35200 115100 35300
rect 115000 35300 115100 35400
rect 115000 35400 115100 35500
rect 115000 35500 115100 35600
rect 115000 35600 115100 35700
rect 115000 35700 115100 35800
rect 115000 35800 115100 35900
rect 115000 35900 115100 36000
rect 115000 36000 115100 36100
rect 115000 36100 115100 36200
rect 115000 36200 115100 36300
rect 115000 36300 115100 36400
rect 115000 36400 115100 36500
rect 115000 36500 115100 36600
rect 115000 36600 115100 36700
rect 115000 36700 115100 36800
rect 115000 36800 115100 36900
rect 115000 36900 115100 37000
rect 115000 37000 115100 37100
rect 115100 21800 115200 21900
rect 115100 21900 115200 22000
rect 115100 22000 115200 22100
rect 115100 22100 115200 22200
rect 115100 22200 115200 22300
rect 115100 22300 115200 22400
rect 115100 22400 115200 22500
rect 115100 22500 115200 22600
rect 115100 22600 115200 22700
rect 115100 22700 115200 22800
rect 115100 22800 115200 22900
rect 115100 22900 115200 23000
rect 115100 23000 115200 23100
rect 115100 23100 115200 23200
rect 115100 23200 115200 23300
rect 115100 23300 115200 23400
rect 115100 23400 115200 23500
rect 115100 23500 115200 23600
rect 115100 23600 115200 23700
rect 115100 23700 115200 23800
rect 115100 23800 115200 23900
rect 115100 23900 115200 24000
rect 115100 24000 115200 24100
rect 115100 24100 115200 24200
rect 115100 24200 115200 24300
rect 115100 24300 115200 24400
rect 115100 24400 115200 24500
rect 115100 24500 115200 24600
rect 115100 24600 115200 24700
rect 115100 27500 115200 27600
rect 115100 27600 115200 27700
rect 115100 27700 115200 27800
rect 115100 27800 115200 27900
rect 115100 27900 115200 28000
rect 115100 28000 115200 28100
rect 115100 28100 115200 28200
rect 115100 28200 115200 28300
rect 115100 28300 115200 28400
rect 115100 28400 115200 28500
rect 115100 28500 115200 28600
rect 115100 28600 115200 28700
rect 115100 28700 115200 28800
rect 115100 28800 115200 28900
rect 115100 28900 115200 29000
rect 115100 29000 115200 29100
rect 115100 29100 115200 29200
rect 115100 29200 115200 29300
rect 115100 29300 115200 29400
rect 115100 29400 115200 29500
rect 115100 29500 115200 29600
rect 115100 29600 115200 29700
rect 115100 29700 115200 29800
rect 115100 29800 115200 29900
rect 115100 29900 115200 30000
rect 115100 30000 115200 30100
rect 115100 30100 115200 30200
rect 115100 30200 115200 30300
rect 115100 30300 115200 30400
rect 115100 30400 115200 30500
rect 115100 30500 115200 30600
rect 115100 30600 115200 30700
rect 115100 30700 115200 30800
rect 115100 30800 115200 30900
rect 115100 30900 115200 31000
rect 115100 31000 115200 31100
rect 115100 31100 115200 31200
rect 115100 31200 115200 31300
rect 115100 31300 115200 31400
rect 115100 31400 115200 31500
rect 115100 31500 115200 31600
rect 115100 31600 115200 31700
rect 115100 31700 115200 31800
rect 115100 31800 115200 31900
rect 115100 31900 115200 32000
rect 115100 32000 115200 32100
rect 115100 32100 115200 32200
rect 115100 32200 115200 32300
rect 115100 32300 115200 32400
rect 115100 32400 115200 32500
rect 115100 32500 115200 32600
rect 115100 32600 115200 32700
rect 115100 32700 115200 32800
rect 115100 32800 115200 32900
rect 115100 32900 115200 33000
rect 115100 33000 115200 33100
rect 115100 33100 115200 33200
rect 115100 33200 115200 33300
rect 115100 33300 115200 33400
rect 115100 33400 115200 33500
rect 115100 33500 115200 33600
rect 115100 33600 115200 33700
rect 115100 33700 115200 33800
rect 115100 33800 115200 33900
rect 115100 33900 115200 34000
rect 115100 34000 115200 34100
rect 115100 34100 115200 34200
rect 115100 34200 115200 34300
rect 115100 34300 115200 34400
rect 115100 34400 115200 34500
rect 115100 34500 115200 34600
rect 115100 34600 115200 34700
rect 115100 34700 115200 34800
rect 115100 34800 115200 34900
rect 115100 34900 115200 35000
rect 115100 35000 115200 35100
rect 115100 35100 115200 35200
rect 115100 35200 115200 35300
rect 115100 35300 115200 35400
rect 115100 35400 115200 35500
rect 115100 35500 115200 35600
rect 115100 35600 115200 35700
rect 115100 35700 115200 35800
rect 115100 35800 115200 35900
rect 115100 35900 115200 36000
rect 115100 36000 115200 36100
rect 115100 36100 115200 36200
rect 115100 36200 115200 36300
rect 115100 36300 115200 36400
rect 115100 36400 115200 36500
rect 115100 36500 115200 36600
rect 115100 36600 115200 36700
rect 115100 36700 115200 36800
rect 115100 36800 115200 36900
rect 115100 36900 115200 37000
rect 115200 21600 115300 21700
rect 115200 21700 115300 21800
rect 115200 21800 115300 21900
rect 115200 21900 115300 22000
rect 115200 22000 115300 22100
rect 115200 22100 115300 22200
rect 115200 22200 115300 22300
rect 115200 22300 115300 22400
rect 115200 22400 115300 22500
rect 115200 22500 115300 22600
rect 115200 22600 115300 22700
rect 115200 22700 115300 22800
rect 115200 22800 115300 22900
rect 115200 22900 115300 23000
rect 115200 23000 115300 23100
rect 115200 23100 115300 23200
rect 115200 23200 115300 23300
rect 115200 23300 115300 23400
rect 115200 23400 115300 23500
rect 115200 23500 115300 23600
rect 115200 23600 115300 23700
rect 115200 23700 115300 23800
rect 115200 23800 115300 23900
rect 115200 23900 115300 24000
rect 115200 24000 115300 24100
rect 115200 24100 115300 24200
rect 115200 24200 115300 24300
rect 115200 24300 115300 24400
rect 115200 24400 115300 24500
rect 115200 24500 115300 24600
rect 115200 24600 115300 24700
rect 115200 24700 115300 24800
rect 115200 27200 115300 27300
rect 115200 27300 115300 27400
rect 115200 27400 115300 27500
rect 115200 27500 115300 27600
rect 115200 27600 115300 27700
rect 115200 27700 115300 27800
rect 115200 27800 115300 27900
rect 115200 27900 115300 28000
rect 115200 28000 115300 28100
rect 115200 28100 115300 28200
rect 115200 28200 115300 28300
rect 115200 28300 115300 28400
rect 115200 28400 115300 28500
rect 115200 28500 115300 28600
rect 115200 28600 115300 28700
rect 115200 28700 115300 28800
rect 115200 28800 115300 28900
rect 115200 28900 115300 29000
rect 115200 29000 115300 29100
rect 115200 29100 115300 29200
rect 115200 29200 115300 29300
rect 115200 29300 115300 29400
rect 115200 29400 115300 29500
rect 115200 29500 115300 29600
rect 115200 29600 115300 29700
rect 115200 29700 115300 29800
rect 115200 29800 115300 29900
rect 115200 29900 115300 30000
rect 115200 30000 115300 30100
rect 115200 30100 115300 30200
rect 115200 30200 115300 30300
rect 115200 30300 115300 30400
rect 115200 30400 115300 30500
rect 115200 30500 115300 30600
rect 115200 30600 115300 30700
rect 115200 30700 115300 30800
rect 115200 30800 115300 30900
rect 115200 30900 115300 31000
rect 115200 31000 115300 31100
rect 115200 31100 115300 31200
rect 115200 31200 115300 31300
rect 115200 31300 115300 31400
rect 115200 31400 115300 31500
rect 115200 31500 115300 31600
rect 115200 31600 115300 31700
rect 115200 31700 115300 31800
rect 115200 31800 115300 31900
rect 115200 31900 115300 32000
rect 115200 32000 115300 32100
rect 115200 32100 115300 32200
rect 115200 32200 115300 32300
rect 115200 32300 115300 32400
rect 115200 32400 115300 32500
rect 115200 33700 115300 33800
rect 115200 33800 115300 33900
rect 115200 33900 115300 34000
rect 115200 34000 115300 34100
rect 115200 34100 115300 34200
rect 115200 34200 115300 34300
rect 115200 34300 115300 34400
rect 115200 34400 115300 34500
rect 115200 34500 115300 34600
rect 115200 34600 115300 34700
rect 115200 34700 115300 34800
rect 115200 34800 115300 34900
rect 115200 34900 115300 35000
rect 115200 35000 115300 35100
rect 115200 35100 115300 35200
rect 115200 35200 115300 35300
rect 115200 35300 115300 35400
rect 115200 35400 115300 35500
rect 115200 35500 115300 35600
rect 115200 35600 115300 35700
rect 115200 35700 115300 35800
rect 115200 35800 115300 35900
rect 115200 35900 115300 36000
rect 115200 36000 115300 36100
rect 115200 36100 115300 36200
rect 115200 36200 115300 36300
rect 115200 36300 115300 36400
rect 115200 36400 115300 36500
rect 115200 36500 115300 36600
rect 115200 36600 115300 36700
rect 115200 36700 115300 36800
rect 115200 36800 115300 36900
rect 115300 21500 115400 21600
rect 115300 21600 115400 21700
rect 115300 21700 115400 21800
rect 115300 21800 115400 21900
rect 115300 21900 115400 22000
rect 115300 22000 115400 22100
rect 115300 22100 115400 22200
rect 115300 22200 115400 22300
rect 115300 22300 115400 22400
rect 115300 22400 115400 22500
rect 115300 22500 115400 22600
rect 115300 22600 115400 22700
rect 115300 22700 115400 22800
rect 115300 22800 115400 22900
rect 115300 22900 115400 23000
rect 115300 23000 115400 23100
rect 115300 23100 115400 23200
rect 115300 23200 115400 23300
rect 115300 23300 115400 23400
rect 115300 23400 115400 23500
rect 115300 23500 115400 23600
rect 115300 23600 115400 23700
rect 115300 23700 115400 23800
rect 115300 23800 115400 23900
rect 115300 23900 115400 24000
rect 115300 24000 115400 24100
rect 115300 24100 115400 24200
rect 115300 24200 115400 24300
rect 115300 24300 115400 24400
rect 115300 24400 115400 24500
rect 115300 24500 115400 24600
rect 115300 24600 115400 24700
rect 115300 24700 115400 24800
rect 115300 24800 115400 24900
rect 115300 24900 115400 25000
rect 115300 26900 115400 27000
rect 115300 27000 115400 27100
rect 115300 27100 115400 27200
rect 115300 27200 115400 27300
rect 115300 27300 115400 27400
rect 115300 27400 115400 27500
rect 115300 27500 115400 27600
rect 115300 27600 115400 27700
rect 115300 27700 115400 27800
rect 115300 27800 115400 27900
rect 115300 27900 115400 28000
rect 115300 28000 115400 28100
rect 115300 28100 115400 28200
rect 115300 28200 115400 28300
rect 115300 28300 115400 28400
rect 115300 28400 115400 28500
rect 115300 28500 115400 28600
rect 115300 28600 115400 28700
rect 115300 28700 115400 28800
rect 115300 28800 115400 28900
rect 115300 28900 115400 29000
rect 115300 29000 115400 29100
rect 115300 29100 115400 29200
rect 115300 29200 115400 29300
rect 115300 29300 115400 29400
rect 115300 29400 115400 29500
rect 115300 29500 115400 29600
rect 115300 29600 115400 29700
rect 115300 29700 115400 29800
rect 115300 29800 115400 29900
rect 115300 29900 115400 30000
rect 115300 30000 115400 30100
rect 115300 30100 115400 30200
rect 115300 30200 115400 30300
rect 115300 30300 115400 30400
rect 115300 30400 115400 30500
rect 115300 30500 115400 30600
rect 115300 30600 115400 30700
rect 115300 30700 115400 30800
rect 115300 30800 115400 30900
rect 115300 30900 115400 31000
rect 115300 31000 115400 31100
rect 115300 31100 115400 31200
rect 115300 31200 115400 31300
rect 115300 31300 115400 31400
rect 115300 31400 115400 31500
rect 115300 31500 115400 31600
rect 115300 31600 115400 31700
rect 115300 31700 115400 31800
rect 115300 31800 115400 31900
rect 115300 31900 115400 32000
rect 115300 32000 115400 32100
rect 115300 34000 115400 34100
rect 115300 34100 115400 34200
rect 115300 34200 115400 34300
rect 115300 34300 115400 34400
rect 115300 34400 115400 34500
rect 115300 34500 115400 34600
rect 115300 34600 115400 34700
rect 115300 34700 115400 34800
rect 115300 34800 115400 34900
rect 115300 34900 115400 35000
rect 115300 35000 115400 35100
rect 115300 35100 115400 35200
rect 115300 35200 115400 35300
rect 115300 35300 115400 35400
rect 115300 35400 115400 35500
rect 115300 35500 115400 35600
rect 115300 35600 115400 35700
rect 115300 35700 115400 35800
rect 115300 35800 115400 35900
rect 115300 35900 115400 36000
rect 115300 36000 115400 36100
rect 115300 36100 115400 36200
rect 115300 36200 115400 36300
rect 115300 36300 115400 36400
rect 115300 36400 115400 36500
rect 115300 36500 115400 36600
rect 115300 36600 115400 36700
rect 115300 36700 115400 36800
rect 115400 21400 115500 21500
rect 115400 21500 115500 21600
rect 115400 21600 115500 21700
rect 115400 21700 115500 21800
rect 115400 21800 115500 21900
rect 115400 21900 115500 22000
rect 115400 22000 115500 22100
rect 115400 22100 115500 22200
rect 115400 22200 115500 22300
rect 115400 22300 115500 22400
rect 115400 22400 115500 22500
rect 115400 22500 115500 22600
rect 115400 22600 115500 22700
rect 115400 22700 115500 22800
rect 115400 22800 115500 22900
rect 115400 22900 115500 23000
rect 115400 23000 115500 23100
rect 115400 23100 115500 23200
rect 115400 23200 115500 23300
rect 115400 23300 115500 23400
rect 115400 23400 115500 23500
rect 115400 23500 115500 23600
rect 115400 23600 115500 23700
rect 115400 23700 115500 23800
rect 115400 23800 115500 23900
rect 115400 23900 115500 24000
rect 115400 24000 115500 24100
rect 115400 24100 115500 24200
rect 115400 24200 115500 24300
rect 115400 24300 115500 24400
rect 115400 24400 115500 24500
rect 115400 24500 115500 24600
rect 115400 24600 115500 24700
rect 115400 24700 115500 24800
rect 115400 24800 115500 24900
rect 115400 24900 115500 25000
rect 115400 25000 115500 25100
rect 115400 25100 115500 25200
rect 115400 26400 115500 26500
rect 115400 26500 115500 26600
rect 115400 26600 115500 26700
rect 115400 26700 115500 26800
rect 115400 26800 115500 26900
rect 115400 26900 115500 27000
rect 115400 27000 115500 27100
rect 115400 27100 115500 27200
rect 115400 27200 115500 27300
rect 115400 27300 115500 27400
rect 115400 27400 115500 27500
rect 115400 27500 115500 27600
rect 115400 27600 115500 27700
rect 115400 27700 115500 27800
rect 115400 27800 115500 27900
rect 115400 27900 115500 28000
rect 115400 28000 115500 28100
rect 115400 28100 115500 28200
rect 115400 28200 115500 28300
rect 115400 28300 115500 28400
rect 115400 28400 115500 28500
rect 115400 28500 115500 28600
rect 115400 28600 115500 28700
rect 115400 28700 115500 28800
rect 115400 28800 115500 28900
rect 115400 28900 115500 29000
rect 115400 29000 115500 29100
rect 115400 29100 115500 29200
rect 115400 29200 115500 29300
rect 115400 29300 115500 29400
rect 115400 29400 115500 29500
rect 115400 29500 115500 29600
rect 115400 29600 115500 29700
rect 115400 29700 115500 29800
rect 115400 29800 115500 29900
rect 115400 29900 115500 30000
rect 115400 30000 115500 30100
rect 115400 30100 115500 30200
rect 115400 30200 115500 30300
rect 115400 30300 115500 30400
rect 115400 30400 115500 30500
rect 115400 30500 115500 30600
rect 115400 30600 115500 30700
rect 115400 30700 115500 30800
rect 115400 30800 115500 30900
rect 115400 30900 115500 31000
rect 115400 31000 115500 31100
rect 115400 31100 115500 31200
rect 115400 31200 115500 31300
rect 115400 31300 115500 31400
rect 115400 31400 115500 31500
rect 115400 31500 115500 31600
rect 115400 31600 115500 31700
rect 115400 31700 115500 31800
rect 115400 34200 115500 34300
rect 115400 34300 115500 34400
rect 115400 34400 115500 34500
rect 115400 34500 115500 34600
rect 115400 34600 115500 34700
rect 115400 34700 115500 34800
rect 115400 34800 115500 34900
rect 115400 34900 115500 35000
rect 115400 35000 115500 35100
rect 115400 35100 115500 35200
rect 115400 35200 115500 35300
rect 115400 35300 115500 35400
rect 115400 35400 115500 35500
rect 115400 35500 115500 35600
rect 115400 35600 115500 35700
rect 115400 35700 115500 35800
rect 115400 35800 115500 35900
rect 115400 35900 115500 36000
rect 115400 36000 115500 36100
rect 115400 36100 115500 36200
rect 115400 36200 115500 36300
rect 115400 36300 115500 36400
rect 115400 36400 115500 36500
rect 115400 36500 115500 36600
rect 115500 21300 115600 21400
rect 115500 21400 115600 21500
rect 115500 21500 115600 21600
rect 115500 21600 115600 21700
rect 115500 21700 115600 21800
rect 115500 21800 115600 21900
rect 115500 21900 115600 22000
rect 115500 22000 115600 22100
rect 115500 22100 115600 22200
rect 115500 22200 115600 22300
rect 115500 22300 115600 22400
rect 115500 22400 115600 22500
rect 115500 22500 115600 22600
rect 115500 22600 115600 22700
rect 115500 22700 115600 22800
rect 115500 22800 115600 22900
rect 115500 22900 115600 23000
rect 115500 23000 115600 23100
rect 115500 23100 115600 23200
rect 115500 23200 115600 23300
rect 115500 23300 115600 23400
rect 115500 23400 115600 23500
rect 115500 23500 115600 23600
rect 115500 23600 115600 23700
rect 115500 23700 115600 23800
rect 115500 23800 115600 23900
rect 115500 23900 115600 24000
rect 115500 24000 115600 24100
rect 115500 24100 115600 24200
rect 115500 24200 115600 24300
rect 115500 24300 115600 24400
rect 115500 24400 115600 24500
rect 115500 24500 115600 24600
rect 115500 24600 115600 24700
rect 115500 24700 115600 24800
rect 115500 24800 115600 24900
rect 115500 24900 115600 25000
rect 115500 25000 115600 25100
rect 115500 25100 115600 25200
rect 115500 25200 115600 25300
rect 115500 25300 115600 25400
rect 115500 25400 115600 25500
rect 115500 25500 115600 25600
rect 115500 25600 115600 25700
rect 115500 25700 115600 25800
rect 115500 25800 115600 25900
rect 115500 25900 115600 26000
rect 115500 26000 115600 26100
rect 115500 26100 115600 26200
rect 115500 26200 115600 26300
rect 115500 26300 115600 26400
rect 115500 26400 115600 26500
rect 115500 26500 115600 26600
rect 115500 26600 115600 26700
rect 115500 26700 115600 26800
rect 115500 26800 115600 26900
rect 115500 26900 115600 27000
rect 115500 27000 115600 27100
rect 115500 27100 115600 27200
rect 115500 27200 115600 27300
rect 115500 27300 115600 27400
rect 115500 27400 115600 27500
rect 115500 27500 115600 27600
rect 115500 27600 115600 27700
rect 115500 27700 115600 27800
rect 115500 27800 115600 27900
rect 115500 27900 115600 28000
rect 115500 28000 115600 28100
rect 115500 28100 115600 28200
rect 115500 28200 115600 28300
rect 115500 28300 115600 28400
rect 115500 28400 115600 28500
rect 115500 28500 115600 28600
rect 115500 28600 115600 28700
rect 115500 28700 115600 28800
rect 115500 28800 115600 28900
rect 115500 28900 115600 29000
rect 115500 29000 115600 29100
rect 115500 29100 115600 29200
rect 115500 29200 115600 29300
rect 115500 29300 115600 29400
rect 115500 29400 115600 29500
rect 115500 29500 115600 29600
rect 115500 29600 115600 29700
rect 115500 29700 115600 29800
rect 115500 29800 115600 29900
rect 115500 29900 115600 30000
rect 115500 30000 115600 30100
rect 115500 30100 115600 30200
rect 115500 30200 115600 30300
rect 115500 30300 115600 30400
rect 115500 30400 115600 30500
rect 115500 30500 115600 30600
rect 115500 30600 115600 30700
rect 115500 30700 115600 30800
rect 115500 30800 115600 30900
rect 115500 30900 115600 31000
rect 115500 31000 115600 31100
rect 115500 31100 115600 31200
rect 115500 31200 115600 31300
rect 115500 31300 115600 31400
rect 115500 34400 115600 34500
rect 115500 34500 115600 34600
rect 115500 34600 115600 34700
rect 115500 34700 115600 34800
rect 115500 34800 115600 34900
rect 115500 34900 115600 35000
rect 115500 35000 115600 35100
rect 115500 35100 115600 35200
rect 115500 35200 115600 35300
rect 115500 35300 115600 35400
rect 115500 35400 115600 35500
rect 115500 35500 115600 35600
rect 115500 35600 115600 35700
rect 115500 35700 115600 35800
rect 115500 35800 115600 35900
rect 115500 35900 115600 36000
rect 115500 36000 115600 36100
rect 115500 36100 115600 36200
rect 115500 36200 115600 36300
rect 115500 36300 115600 36400
rect 115600 21200 115700 21300
rect 115600 21300 115700 21400
rect 115600 21400 115700 21500
rect 115600 21500 115700 21600
rect 115600 21600 115700 21700
rect 115600 21700 115700 21800
rect 115600 21800 115700 21900
rect 115600 21900 115700 22000
rect 115600 22000 115700 22100
rect 115600 22100 115700 22200
rect 115600 22200 115700 22300
rect 115600 22300 115700 22400
rect 115600 22400 115700 22500
rect 115600 22500 115700 22600
rect 115600 22600 115700 22700
rect 115600 22700 115700 22800
rect 115600 22800 115700 22900
rect 115600 22900 115700 23000
rect 115600 23000 115700 23100
rect 115600 23100 115700 23200
rect 115600 23200 115700 23300
rect 115600 23300 115700 23400
rect 115600 23400 115700 23500
rect 115600 23500 115700 23600
rect 115600 23600 115700 23700
rect 115600 23700 115700 23800
rect 115600 23800 115700 23900
rect 115600 23900 115700 24000
rect 115600 24000 115700 24100
rect 115600 24100 115700 24200
rect 115600 24200 115700 24300
rect 115600 24300 115700 24400
rect 115600 24400 115700 24500
rect 115600 24500 115700 24600
rect 115600 24600 115700 24700
rect 115600 24700 115700 24800
rect 115600 24800 115700 24900
rect 115600 24900 115700 25000
rect 115600 25000 115700 25100
rect 115600 25100 115700 25200
rect 115600 25200 115700 25300
rect 115600 25300 115700 25400
rect 115600 25400 115700 25500
rect 115600 25500 115700 25600
rect 115600 25600 115700 25700
rect 115600 25700 115700 25800
rect 115600 25800 115700 25900
rect 115600 25900 115700 26000
rect 115600 26000 115700 26100
rect 115600 26100 115700 26200
rect 115600 26200 115700 26300
rect 115600 26300 115700 26400
rect 115600 26400 115700 26500
rect 115600 26500 115700 26600
rect 115600 26600 115700 26700
rect 115600 26700 115700 26800
rect 115600 26800 115700 26900
rect 115600 26900 115700 27000
rect 115600 27000 115700 27100
rect 115600 27100 115700 27200
rect 115600 27200 115700 27300
rect 115600 27300 115700 27400
rect 115600 27400 115700 27500
rect 115600 27500 115700 27600
rect 115600 27600 115700 27700
rect 115600 27700 115700 27800
rect 115600 27800 115700 27900
rect 115600 27900 115700 28000
rect 115600 28000 115700 28100
rect 115600 28100 115700 28200
rect 115600 28200 115700 28300
rect 115600 28300 115700 28400
rect 115600 28400 115700 28500
rect 115600 28500 115700 28600
rect 115600 28600 115700 28700
rect 115600 28700 115700 28800
rect 115600 28800 115700 28900
rect 115600 28900 115700 29000
rect 115600 29000 115700 29100
rect 115600 29100 115700 29200
rect 115600 29200 115700 29300
rect 115600 29300 115700 29400
rect 115600 29400 115700 29500
rect 115600 29500 115700 29600
rect 115600 29600 115700 29700
rect 115600 29700 115700 29800
rect 115600 29800 115700 29900
rect 115600 29900 115700 30000
rect 115600 30000 115700 30100
rect 115600 30100 115700 30200
rect 115600 30200 115700 30300
rect 115600 30300 115700 30400
rect 115600 30400 115700 30500
rect 115600 30500 115700 30600
rect 115600 30600 115700 30700
rect 115600 30700 115700 30800
rect 115600 30800 115700 30900
rect 115600 30900 115700 31000
rect 115600 31000 115700 31100
rect 115600 34600 115700 34700
rect 115600 34700 115700 34800
rect 115600 34800 115700 34900
rect 115600 34900 115700 35000
rect 115600 35000 115700 35100
rect 115600 35100 115700 35200
rect 115600 35200 115700 35300
rect 115600 35300 115700 35400
rect 115600 35400 115700 35500
rect 115600 35500 115700 35600
rect 115600 35600 115700 35700
rect 115600 35700 115700 35800
rect 115600 35800 115700 35900
rect 115600 35900 115700 36000
rect 115600 36000 115700 36100
rect 115600 36100 115700 36200
rect 115700 21100 115800 21200
rect 115700 21200 115800 21300
rect 115700 21300 115800 21400
rect 115700 21400 115800 21500
rect 115700 21500 115800 21600
rect 115700 21600 115800 21700
rect 115700 21700 115800 21800
rect 115700 21800 115800 21900
rect 115700 21900 115800 22000
rect 115700 22000 115800 22100
rect 115700 22100 115800 22200
rect 115700 22200 115800 22300
rect 115700 22300 115800 22400
rect 115700 22400 115800 22500
rect 115700 22500 115800 22600
rect 115700 22600 115800 22700
rect 115700 22700 115800 22800
rect 115700 22800 115800 22900
rect 115700 22900 115800 23000
rect 115700 23000 115800 23100
rect 115700 23100 115800 23200
rect 115700 23200 115800 23300
rect 115700 23300 115800 23400
rect 115700 23400 115800 23500
rect 115700 23500 115800 23600
rect 115700 23600 115800 23700
rect 115700 23700 115800 23800
rect 115700 23800 115800 23900
rect 115700 23900 115800 24000
rect 115700 24000 115800 24100
rect 115700 24100 115800 24200
rect 115700 24200 115800 24300
rect 115700 24300 115800 24400
rect 115700 24400 115800 24500
rect 115700 24500 115800 24600
rect 115700 24600 115800 24700
rect 115700 24700 115800 24800
rect 115700 24800 115800 24900
rect 115700 24900 115800 25000
rect 115700 25000 115800 25100
rect 115700 25100 115800 25200
rect 115700 25200 115800 25300
rect 115700 25300 115800 25400
rect 115700 25400 115800 25500
rect 115700 25500 115800 25600
rect 115700 25600 115800 25700
rect 115700 25700 115800 25800
rect 115700 25800 115800 25900
rect 115700 25900 115800 26000
rect 115700 26000 115800 26100
rect 115700 26100 115800 26200
rect 115700 26200 115800 26300
rect 115700 26300 115800 26400
rect 115700 26400 115800 26500
rect 115700 26500 115800 26600
rect 115700 26600 115800 26700
rect 115700 26700 115800 26800
rect 115700 26800 115800 26900
rect 115700 26900 115800 27000
rect 115700 27000 115800 27100
rect 115700 27100 115800 27200
rect 115700 27200 115800 27300
rect 115700 27300 115800 27400
rect 115700 27400 115800 27500
rect 115700 27500 115800 27600
rect 115700 27600 115800 27700
rect 115700 27700 115800 27800
rect 115700 27800 115800 27900
rect 115700 27900 115800 28000
rect 115700 28000 115800 28100
rect 115700 28100 115800 28200
rect 115700 28200 115800 28300
rect 115700 28300 115800 28400
rect 115700 28400 115800 28500
rect 115700 28500 115800 28600
rect 115700 28600 115800 28700
rect 115700 28700 115800 28800
rect 115700 28800 115800 28900
rect 115700 28900 115800 29000
rect 115700 29000 115800 29100
rect 115700 29100 115800 29200
rect 115700 29200 115800 29300
rect 115700 29300 115800 29400
rect 115700 29400 115800 29500
rect 115700 29500 115800 29600
rect 115700 29600 115800 29700
rect 115700 29700 115800 29800
rect 115700 29800 115800 29900
rect 115700 29900 115800 30000
rect 115700 30000 115800 30100
rect 115700 30100 115800 30200
rect 115700 30200 115800 30300
rect 115700 30300 115800 30400
rect 115700 30400 115800 30500
rect 115700 30500 115800 30600
rect 115700 30600 115800 30700
rect 115700 30700 115800 30800
rect 115700 35100 115800 35200
rect 115700 35200 115800 35300
rect 115700 35300 115800 35400
rect 115700 35400 115800 35500
rect 115700 35500 115800 35600
rect 115700 35600 115800 35700
rect 115700 35700 115800 35800
rect 115800 21100 115900 21200
rect 115800 21200 115900 21300
rect 115800 21300 115900 21400
rect 115800 21400 115900 21500
rect 115800 21500 115900 21600
rect 115800 21600 115900 21700
rect 115800 21700 115900 21800
rect 115800 21800 115900 21900
rect 115800 21900 115900 22000
rect 115800 22000 115900 22100
rect 115800 22100 115900 22200
rect 115800 22200 115900 22300
rect 115800 22300 115900 22400
rect 115800 22400 115900 22500
rect 115800 22500 115900 22600
rect 115800 22600 115900 22700
rect 115800 22700 115900 22800
rect 115800 22800 115900 22900
rect 115800 22900 115900 23000
rect 115800 23000 115900 23100
rect 115800 23100 115900 23200
rect 115800 23200 115900 23300
rect 115800 23300 115900 23400
rect 115800 23400 115900 23500
rect 115800 23500 115900 23600
rect 115800 23600 115900 23700
rect 115800 23700 115900 23800
rect 115800 23800 115900 23900
rect 115800 23900 115900 24000
rect 115800 24000 115900 24100
rect 115800 24100 115900 24200
rect 115800 24200 115900 24300
rect 115800 24300 115900 24400
rect 115800 24400 115900 24500
rect 115800 24500 115900 24600
rect 115800 24600 115900 24700
rect 115800 24700 115900 24800
rect 115800 24800 115900 24900
rect 115800 24900 115900 25000
rect 115800 25000 115900 25100
rect 115800 25100 115900 25200
rect 115800 25200 115900 25300
rect 115800 25300 115900 25400
rect 115800 25400 115900 25500
rect 115800 25500 115900 25600
rect 115800 25600 115900 25700
rect 115800 25700 115900 25800
rect 115800 25800 115900 25900
rect 115800 25900 115900 26000
rect 115800 26000 115900 26100
rect 115800 26100 115900 26200
rect 115800 26200 115900 26300
rect 115800 26300 115900 26400
rect 115800 26400 115900 26500
rect 115800 26500 115900 26600
rect 115800 26600 115900 26700
rect 115800 26700 115900 26800
rect 115800 26800 115900 26900
rect 115800 26900 115900 27000
rect 115800 27000 115900 27100
rect 115800 27100 115900 27200
rect 115800 27200 115900 27300
rect 115800 27300 115900 27400
rect 115800 27400 115900 27500
rect 115800 27500 115900 27600
rect 115800 27600 115900 27700
rect 115800 27700 115900 27800
rect 115800 27800 115900 27900
rect 115800 27900 115900 28000
rect 115800 28000 115900 28100
rect 115800 28100 115900 28200
rect 115800 28200 115900 28300
rect 115800 28300 115900 28400
rect 115800 28400 115900 28500
rect 115800 28500 115900 28600
rect 115800 28600 115900 28700
rect 115800 28700 115900 28800
rect 115800 28800 115900 28900
rect 115800 28900 115900 29000
rect 115800 29000 115900 29100
rect 115800 29100 115900 29200
rect 115800 29200 115900 29300
rect 115800 29300 115900 29400
rect 115800 29400 115900 29500
rect 115800 29500 115900 29600
rect 115800 29600 115900 29700
rect 115800 29700 115900 29800
rect 115800 29800 115900 29900
rect 115800 29900 115900 30000
rect 115800 30000 115900 30100
rect 115800 30100 115900 30200
rect 115800 30200 115900 30300
rect 115800 30300 115900 30400
rect 115800 30400 115900 30500
rect 115900 21000 116000 21100
rect 115900 21100 116000 21200
rect 115900 21200 116000 21300
rect 115900 21300 116000 21400
rect 115900 21400 116000 21500
rect 115900 21500 116000 21600
rect 115900 21600 116000 21700
rect 115900 21700 116000 21800
rect 115900 21800 116000 21900
rect 115900 21900 116000 22000
rect 115900 22000 116000 22100
rect 115900 22100 116000 22200
rect 115900 22200 116000 22300
rect 115900 22300 116000 22400
rect 115900 22400 116000 22500
rect 115900 22500 116000 22600
rect 115900 22600 116000 22700
rect 115900 22700 116000 22800
rect 115900 22800 116000 22900
rect 115900 22900 116000 23000
rect 115900 23000 116000 23100
rect 115900 23100 116000 23200
rect 115900 23200 116000 23300
rect 115900 23300 116000 23400
rect 115900 23400 116000 23500
rect 115900 23500 116000 23600
rect 115900 23600 116000 23700
rect 115900 23700 116000 23800
rect 115900 23800 116000 23900
rect 115900 23900 116000 24000
rect 115900 24000 116000 24100
rect 115900 24100 116000 24200
rect 115900 24200 116000 24300
rect 115900 24300 116000 24400
rect 115900 24400 116000 24500
rect 115900 24500 116000 24600
rect 115900 24600 116000 24700
rect 115900 24700 116000 24800
rect 115900 24800 116000 24900
rect 115900 24900 116000 25000
rect 115900 25000 116000 25100
rect 115900 25100 116000 25200
rect 115900 25200 116000 25300
rect 115900 25300 116000 25400
rect 115900 25400 116000 25500
rect 115900 25500 116000 25600
rect 115900 25600 116000 25700
rect 115900 25700 116000 25800
rect 115900 25800 116000 25900
rect 115900 25900 116000 26000
rect 115900 26000 116000 26100
rect 115900 26100 116000 26200
rect 115900 26200 116000 26300
rect 115900 26300 116000 26400
rect 115900 26400 116000 26500
rect 115900 26500 116000 26600
rect 115900 26600 116000 26700
rect 115900 26700 116000 26800
rect 115900 26800 116000 26900
rect 115900 26900 116000 27000
rect 115900 27000 116000 27100
rect 115900 27100 116000 27200
rect 115900 27200 116000 27300
rect 115900 27300 116000 27400
rect 115900 27400 116000 27500
rect 115900 27500 116000 27600
rect 115900 27600 116000 27700
rect 115900 27700 116000 27800
rect 115900 27800 116000 27900
rect 115900 27900 116000 28000
rect 115900 28000 116000 28100
rect 115900 28100 116000 28200
rect 115900 28200 116000 28300
rect 115900 28300 116000 28400
rect 115900 28400 116000 28500
rect 115900 28500 116000 28600
rect 115900 28600 116000 28700
rect 115900 28700 116000 28800
rect 115900 28800 116000 28900
rect 115900 28900 116000 29000
rect 115900 29000 116000 29100
rect 115900 29100 116000 29200
rect 115900 29200 116000 29300
rect 115900 29300 116000 29400
rect 115900 29400 116000 29500
rect 115900 29500 116000 29600
rect 115900 29600 116000 29700
rect 115900 29700 116000 29800
rect 115900 29800 116000 29900
rect 115900 29900 116000 30000
rect 115900 30000 116000 30100
rect 115900 30100 116000 30200
rect 116000 20900 116100 21000
rect 116000 21000 116100 21100
rect 116000 21100 116100 21200
rect 116000 21200 116100 21300
rect 116000 21300 116100 21400
rect 116000 21400 116100 21500
rect 116000 21500 116100 21600
rect 116000 21600 116100 21700
rect 116000 21700 116100 21800
rect 116000 21800 116100 21900
rect 116000 21900 116100 22000
rect 116000 22000 116100 22100
rect 116000 22100 116100 22200
rect 116000 22200 116100 22300
rect 116000 22300 116100 22400
rect 116000 22400 116100 22500
rect 116000 22500 116100 22600
rect 116000 22600 116100 22700
rect 116000 22700 116100 22800
rect 116000 22800 116100 22900
rect 116000 22900 116100 23000
rect 116000 23000 116100 23100
rect 116000 23100 116100 23200
rect 116000 23200 116100 23300
rect 116000 23300 116100 23400
rect 116000 23400 116100 23500
rect 116000 23500 116100 23600
rect 116000 23600 116100 23700
rect 116000 23700 116100 23800
rect 116000 23800 116100 23900
rect 116000 23900 116100 24000
rect 116000 24000 116100 24100
rect 116000 24100 116100 24200
rect 116000 24200 116100 24300
rect 116000 24300 116100 24400
rect 116000 24400 116100 24500
rect 116000 24500 116100 24600
rect 116000 24600 116100 24700
rect 116000 24700 116100 24800
rect 116000 24800 116100 24900
rect 116000 24900 116100 25000
rect 116000 25000 116100 25100
rect 116000 25100 116100 25200
rect 116000 25200 116100 25300
rect 116000 25300 116100 25400
rect 116000 25400 116100 25500
rect 116000 25500 116100 25600
rect 116000 25600 116100 25700
rect 116000 25700 116100 25800
rect 116000 25800 116100 25900
rect 116000 25900 116100 26000
rect 116000 26000 116100 26100
rect 116000 26100 116100 26200
rect 116000 26200 116100 26300
rect 116000 26300 116100 26400
rect 116000 26400 116100 26500
rect 116000 26500 116100 26600
rect 116000 26600 116100 26700
rect 116000 26700 116100 26800
rect 116000 26800 116100 26900
rect 116000 26900 116100 27000
rect 116000 27000 116100 27100
rect 116000 27100 116100 27200
rect 116000 27200 116100 27300
rect 116000 27300 116100 27400
rect 116000 27400 116100 27500
rect 116000 27500 116100 27600
rect 116000 27600 116100 27700
rect 116000 27700 116100 27800
rect 116000 27800 116100 27900
rect 116000 27900 116100 28000
rect 116000 28000 116100 28100
rect 116000 28100 116100 28200
rect 116000 28200 116100 28300
rect 116000 28300 116100 28400
rect 116000 28400 116100 28500
rect 116000 28500 116100 28600
rect 116000 28600 116100 28700
rect 116000 28700 116100 28800
rect 116000 28800 116100 28900
rect 116000 28900 116100 29000
rect 116000 29000 116100 29100
rect 116000 29100 116100 29200
rect 116000 29200 116100 29300
rect 116000 29300 116100 29400
rect 116000 29400 116100 29500
rect 116000 29500 116100 29600
rect 116000 29600 116100 29700
rect 116000 29700 116100 29800
rect 116000 29800 116100 29900
rect 116000 29900 116100 30000
rect 116100 20900 116200 21000
rect 116100 21000 116200 21100
rect 116100 21100 116200 21200
rect 116100 21200 116200 21300
rect 116100 21300 116200 21400
rect 116100 21400 116200 21500
rect 116100 21500 116200 21600
rect 116100 21600 116200 21700
rect 116100 21700 116200 21800
rect 116100 21800 116200 21900
rect 116100 21900 116200 22000
rect 116100 22000 116200 22100
rect 116100 22100 116200 22200
rect 116100 22200 116200 22300
rect 116100 22300 116200 22400
rect 116100 22400 116200 22500
rect 116100 22500 116200 22600
rect 116100 22600 116200 22700
rect 116100 22700 116200 22800
rect 116100 22800 116200 22900
rect 116100 22900 116200 23000
rect 116100 23000 116200 23100
rect 116100 23100 116200 23200
rect 116100 23200 116200 23300
rect 116100 23300 116200 23400
rect 116100 23400 116200 23500
rect 116100 23500 116200 23600
rect 116100 23600 116200 23700
rect 116100 23700 116200 23800
rect 116100 23800 116200 23900
rect 116100 23900 116200 24000
rect 116100 24000 116200 24100
rect 116100 24100 116200 24200
rect 116100 24200 116200 24300
rect 116100 24300 116200 24400
rect 116100 24400 116200 24500
rect 116100 24500 116200 24600
rect 116100 24600 116200 24700
rect 116100 24700 116200 24800
rect 116100 24800 116200 24900
rect 116100 24900 116200 25000
rect 116100 25000 116200 25100
rect 116100 25100 116200 25200
rect 116100 25200 116200 25300
rect 116100 25300 116200 25400
rect 116100 25400 116200 25500
rect 116100 25500 116200 25600
rect 116100 25600 116200 25700
rect 116100 25700 116200 25800
rect 116100 25800 116200 25900
rect 116100 25900 116200 26000
rect 116100 26000 116200 26100
rect 116100 26100 116200 26200
rect 116100 26200 116200 26300
rect 116100 26300 116200 26400
rect 116100 26400 116200 26500
rect 116100 26500 116200 26600
rect 116100 26600 116200 26700
rect 116100 26700 116200 26800
rect 116100 26800 116200 26900
rect 116100 26900 116200 27000
rect 116100 27000 116200 27100
rect 116100 27100 116200 27200
rect 116100 27200 116200 27300
rect 116100 27300 116200 27400
rect 116100 27400 116200 27500
rect 116100 27500 116200 27600
rect 116100 27600 116200 27700
rect 116100 27700 116200 27800
rect 116100 27800 116200 27900
rect 116100 27900 116200 28000
rect 116100 28000 116200 28100
rect 116100 28100 116200 28200
rect 116100 28200 116200 28300
rect 116100 28300 116200 28400
rect 116100 28400 116200 28500
rect 116100 28500 116200 28600
rect 116100 28600 116200 28700
rect 116100 28700 116200 28800
rect 116100 28800 116200 28900
rect 116100 28900 116200 29000
rect 116100 29000 116200 29100
rect 116100 29100 116200 29200
rect 116100 29200 116200 29300
rect 116100 29300 116200 29400
rect 116100 29400 116200 29500
rect 116100 29500 116200 29600
rect 116100 29600 116200 29700
rect 116200 20800 116300 20900
rect 116200 20900 116300 21000
rect 116200 21000 116300 21100
rect 116200 21100 116300 21200
rect 116200 21200 116300 21300
rect 116200 21300 116300 21400
rect 116200 21400 116300 21500
rect 116200 21500 116300 21600
rect 116200 21600 116300 21700
rect 116200 21700 116300 21800
rect 116200 21800 116300 21900
rect 116200 21900 116300 22000
rect 116200 22000 116300 22100
rect 116200 22100 116300 22200
rect 116200 22200 116300 22300
rect 116200 22300 116300 22400
rect 116200 22400 116300 22500
rect 116200 22500 116300 22600
rect 116200 22600 116300 22700
rect 116200 22700 116300 22800
rect 116200 22800 116300 22900
rect 116200 22900 116300 23000
rect 116200 23000 116300 23100
rect 116200 23100 116300 23200
rect 116200 23200 116300 23300
rect 116200 23300 116300 23400
rect 116200 23400 116300 23500
rect 116200 23500 116300 23600
rect 116200 23600 116300 23700
rect 116200 23700 116300 23800
rect 116200 23800 116300 23900
rect 116200 23900 116300 24000
rect 116200 24000 116300 24100
rect 116200 24100 116300 24200
rect 116200 24200 116300 24300
rect 116200 24300 116300 24400
rect 116200 24400 116300 24500
rect 116200 24500 116300 24600
rect 116200 24600 116300 24700
rect 116200 24700 116300 24800
rect 116200 24800 116300 24900
rect 116200 24900 116300 25000
rect 116200 25000 116300 25100
rect 116200 25100 116300 25200
rect 116200 25200 116300 25300
rect 116200 25300 116300 25400
rect 116200 25400 116300 25500
rect 116200 25500 116300 25600
rect 116200 25600 116300 25700
rect 116200 25700 116300 25800
rect 116200 25800 116300 25900
rect 116200 25900 116300 26000
rect 116200 26000 116300 26100
rect 116200 26100 116300 26200
rect 116200 26200 116300 26300
rect 116200 26300 116300 26400
rect 116200 26400 116300 26500
rect 116200 26500 116300 26600
rect 116200 26600 116300 26700
rect 116200 26700 116300 26800
rect 116200 26800 116300 26900
rect 116200 26900 116300 27000
rect 116200 27000 116300 27100
rect 116200 27100 116300 27200
rect 116200 27200 116300 27300
rect 116200 27300 116300 27400
rect 116200 27400 116300 27500
rect 116200 27500 116300 27600
rect 116200 27600 116300 27700
rect 116200 27700 116300 27800
rect 116200 27800 116300 27900
rect 116200 27900 116300 28000
rect 116200 28000 116300 28100
rect 116200 28100 116300 28200
rect 116200 28200 116300 28300
rect 116200 28300 116300 28400
rect 116200 28400 116300 28500
rect 116200 28500 116300 28600
rect 116200 28600 116300 28700
rect 116200 28700 116300 28800
rect 116200 28800 116300 28900
rect 116200 28900 116300 29000
rect 116200 29000 116300 29100
rect 116200 29100 116300 29200
rect 116200 29200 116300 29300
rect 116200 29300 116300 29400
rect 116300 20800 116400 20900
rect 116300 20900 116400 21000
rect 116300 21000 116400 21100
rect 116300 21100 116400 21200
rect 116300 21200 116400 21300
rect 116300 21300 116400 21400
rect 116300 21400 116400 21500
rect 116300 21500 116400 21600
rect 116300 21600 116400 21700
rect 116300 21700 116400 21800
rect 116300 21800 116400 21900
rect 116300 21900 116400 22000
rect 116300 22000 116400 22100
rect 116300 22100 116400 22200
rect 116300 22200 116400 22300
rect 116300 22300 116400 22400
rect 116300 22400 116400 22500
rect 116300 22500 116400 22600
rect 116300 22600 116400 22700
rect 116300 22700 116400 22800
rect 116300 22800 116400 22900
rect 116300 22900 116400 23000
rect 116300 23000 116400 23100
rect 116300 23100 116400 23200
rect 116300 23200 116400 23300
rect 116300 23300 116400 23400
rect 116300 23400 116400 23500
rect 116300 23500 116400 23600
rect 116300 23600 116400 23700
rect 116300 23700 116400 23800
rect 116300 23800 116400 23900
rect 116300 23900 116400 24000
rect 116300 24000 116400 24100
rect 116300 24100 116400 24200
rect 116300 24200 116400 24300
rect 116300 24300 116400 24400
rect 116300 24400 116400 24500
rect 116300 24500 116400 24600
rect 116300 24600 116400 24700
rect 116300 24700 116400 24800
rect 116300 24800 116400 24900
rect 116300 24900 116400 25000
rect 116300 25000 116400 25100
rect 116300 25100 116400 25200
rect 116300 25200 116400 25300
rect 116300 25300 116400 25400
rect 116300 25400 116400 25500
rect 116300 25500 116400 25600
rect 116300 25600 116400 25700
rect 116300 25700 116400 25800
rect 116300 25800 116400 25900
rect 116300 25900 116400 26000
rect 116300 26000 116400 26100
rect 116300 26100 116400 26200
rect 116300 26200 116400 26300
rect 116300 26300 116400 26400
rect 116300 26400 116400 26500
rect 116300 26500 116400 26600
rect 116300 26600 116400 26700
rect 116300 26700 116400 26800
rect 116300 26800 116400 26900
rect 116300 26900 116400 27000
rect 116300 27000 116400 27100
rect 116300 27100 116400 27200
rect 116300 27200 116400 27300
rect 116300 27300 116400 27400
rect 116300 27400 116400 27500
rect 116300 27500 116400 27600
rect 116300 27600 116400 27700
rect 116300 27700 116400 27800
rect 116300 27800 116400 27900
rect 116300 27900 116400 28000
rect 116300 28000 116400 28100
rect 116300 28100 116400 28200
rect 116300 28200 116400 28300
rect 116300 28300 116400 28400
rect 116300 28400 116400 28500
rect 116300 28500 116400 28600
rect 116300 28600 116400 28700
rect 116300 28700 116400 28800
rect 116300 28800 116400 28900
rect 116300 28900 116400 29000
rect 116300 29000 116400 29100
rect 116400 20800 116500 20900
rect 116400 20900 116500 21000
rect 116400 21000 116500 21100
rect 116400 21100 116500 21200
rect 116400 21200 116500 21300
rect 116400 21300 116500 21400
rect 116400 21400 116500 21500
rect 116400 21500 116500 21600
rect 116400 21600 116500 21700
rect 116400 21700 116500 21800
rect 116400 21800 116500 21900
rect 116400 21900 116500 22000
rect 116400 22000 116500 22100
rect 116400 22100 116500 22200
rect 116400 22200 116500 22300
rect 116400 22300 116500 22400
rect 116400 22400 116500 22500
rect 116400 22500 116500 22600
rect 116400 22600 116500 22700
rect 116400 22700 116500 22800
rect 116400 22800 116500 22900
rect 116400 22900 116500 23000
rect 116400 23000 116500 23100
rect 116400 23100 116500 23200
rect 116400 23200 116500 23300
rect 116400 23300 116500 23400
rect 116400 23400 116500 23500
rect 116400 23500 116500 23600
rect 116400 23600 116500 23700
rect 116400 23700 116500 23800
rect 116400 23800 116500 23900
rect 116400 23900 116500 24000
rect 116400 24000 116500 24100
rect 116400 24100 116500 24200
rect 116400 24200 116500 24300
rect 116400 24300 116500 24400
rect 116400 24400 116500 24500
rect 116400 24500 116500 24600
rect 116400 24600 116500 24700
rect 116400 24700 116500 24800
rect 116400 24800 116500 24900
rect 116400 24900 116500 25000
rect 116400 25000 116500 25100
rect 116400 25100 116500 25200
rect 116400 25200 116500 25300
rect 116400 25300 116500 25400
rect 116400 25400 116500 25500
rect 116400 25500 116500 25600
rect 116400 25600 116500 25700
rect 116400 25700 116500 25800
rect 116400 25800 116500 25900
rect 116400 25900 116500 26000
rect 116400 26000 116500 26100
rect 116400 26100 116500 26200
rect 116400 26200 116500 26300
rect 116400 26300 116500 26400
rect 116400 26400 116500 26500
rect 116400 26500 116500 26600
rect 116400 26600 116500 26700
rect 116400 26700 116500 26800
rect 116400 26800 116500 26900
rect 116400 26900 116500 27000
rect 116400 27000 116500 27100
rect 116400 27100 116500 27200
rect 116400 27200 116500 27300
rect 116400 27300 116500 27400
rect 116400 27400 116500 27500
rect 116400 27500 116500 27600
rect 116400 27600 116500 27700
rect 116400 27700 116500 27800
rect 116400 27800 116500 27900
rect 116400 27900 116500 28000
rect 116400 28000 116500 28100
rect 116400 28100 116500 28200
rect 116400 28200 116500 28300
rect 116400 28300 116500 28400
rect 116400 28400 116500 28500
rect 116400 28500 116500 28600
rect 116400 28600 116500 28700
rect 116400 28700 116500 28800
rect 116500 20800 116600 20900
rect 116500 20900 116600 21000
rect 116500 21000 116600 21100
rect 116500 21100 116600 21200
rect 116500 21200 116600 21300
rect 116500 21300 116600 21400
rect 116500 21400 116600 21500
rect 116500 21500 116600 21600
rect 116500 21600 116600 21700
rect 116500 21700 116600 21800
rect 116500 21800 116600 21900
rect 116500 21900 116600 22000
rect 116500 22000 116600 22100
rect 116500 22100 116600 22200
rect 116500 22200 116600 22300
rect 116500 22300 116600 22400
rect 116500 22400 116600 22500
rect 116500 22500 116600 22600
rect 116500 22600 116600 22700
rect 116500 22700 116600 22800
rect 116500 22800 116600 22900
rect 116500 22900 116600 23000
rect 116500 23000 116600 23100
rect 116500 23100 116600 23200
rect 116500 23200 116600 23300
rect 116500 23300 116600 23400
rect 116500 23400 116600 23500
rect 116500 23500 116600 23600
rect 116500 23600 116600 23700
rect 116500 23700 116600 23800
rect 116500 23800 116600 23900
rect 116500 23900 116600 24000
rect 116500 24000 116600 24100
rect 116500 24100 116600 24200
rect 116500 24200 116600 24300
rect 116500 24300 116600 24400
rect 116500 24400 116600 24500
rect 116500 24500 116600 24600
rect 116500 24600 116600 24700
rect 116500 24700 116600 24800
rect 116500 24800 116600 24900
rect 116500 24900 116600 25000
rect 116500 25000 116600 25100
rect 116500 25100 116600 25200
rect 116500 25200 116600 25300
rect 116500 25300 116600 25400
rect 116500 25400 116600 25500
rect 116500 25500 116600 25600
rect 116500 25600 116600 25700
rect 116500 25700 116600 25800
rect 116500 25800 116600 25900
rect 116500 25900 116600 26000
rect 116500 26000 116600 26100
rect 116500 26100 116600 26200
rect 116500 26200 116600 26300
rect 116500 26300 116600 26400
rect 116500 26400 116600 26500
rect 116500 26500 116600 26600
rect 116500 26600 116600 26700
rect 116500 26700 116600 26800
rect 116500 26800 116600 26900
rect 116500 26900 116600 27000
rect 116500 27000 116600 27100
rect 116500 27100 116600 27200
rect 116500 27200 116600 27300
rect 116500 27300 116600 27400
rect 116500 27400 116600 27500
rect 116500 27500 116600 27600
rect 116500 27600 116600 27700
rect 116500 27700 116600 27800
rect 116500 27800 116600 27900
rect 116500 27900 116600 28000
rect 116500 28000 116600 28100
rect 116500 28100 116600 28200
rect 116500 28200 116600 28300
rect 116500 28300 116600 28400
rect 116500 28400 116600 28500
rect 116600 20700 116700 20800
rect 116600 20800 116700 20900
rect 116600 20900 116700 21000
rect 116600 21000 116700 21100
rect 116600 21100 116700 21200
rect 116600 21200 116700 21300
rect 116600 21300 116700 21400
rect 116600 21400 116700 21500
rect 116600 21500 116700 21600
rect 116600 21600 116700 21700
rect 116600 21700 116700 21800
rect 116600 21800 116700 21900
rect 116600 21900 116700 22000
rect 116600 22000 116700 22100
rect 116600 22100 116700 22200
rect 116600 22200 116700 22300
rect 116600 22300 116700 22400
rect 116600 22400 116700 22500
rect 116600 22500 116700 22600
rect 116600 22600 116700 22700
rect 116600 22700 116700 22800
rect 116600 22800 116700 22900
rect 116600 22900 116700 23000
rect 116600 23000 116700 23100
rect 116600 23100 116700 23200
rect 116600 23800 116700 23900
rect 116600 23900 116700 24000
rect 116600 24000 116700 24100
rect 116600 24100 116700 24200
rect 116600 24200 116700 24300
rect 116600 24300 116700 24400
rect 116600 24400 116700 24500
rect 116600 24500 116700 24600
rect 116600 24600 116700 24700
rect 116600 24700 116700 24800
rect 116600 24800 116700 24900
rect 116600 24900 116700 25000
rect 116600 25000 116700 25100
rect 116600 25100 116700 25200
rect 116600 25200 116700 25300
rect 116600 25300 116700 25400
rect 116600 25400 116700 25500
rect 116600 25500 116700 25600
rect 116600 25600 116700 25700
rect 116600 25700 116700 25800
rect 116600 25800 116700 25900
rect 116600 25900 116700 26000
rect 116600 26000 116700 26100
rect 116600 26100 116700 26200
rect 116600 26200 116700 26300
rect 116600 26300 116700 26400
rect 116600 26400 116700 26500
rect 116600 26500 116700 26600
rect 116600 26600 116700 26700
rect 116600 26700 116700 26800
rect 116600 26800 116700 26900
rect 116600 26900 116700 27000
rect 116600 27000 116700 27100
rect 116600 27100 116700 27200
rect 116600 27200 116700 27300
rect 116600 27300 116700 27400
rect 116600 27400 116700 27500
rect 116600 27500 116700 27600
rect 116600 27600 116700 27700
rect 116600 27700 116700 27800
rect 116600 27800 116700 27900
rect 116600 27900 116700 28000
rect 116600 28000 116700 28100
rect 116600 28100 116700 28200
rect 116600 28200 116700 28300
rect 116700 20700 116800 20800
rect 116700 20800 116800 20900
rect 116700 20900 116800 21000
rect 116700 21000 116800 21100
rect 116700 21100 116800 21200
rect 116700 21200 116800 21300
rect 116700 21300 116800 21400
rect 116700 21400 116800 21500
rect 116700 21500 116800 21600
rect 116700 21600 116800 21700
rect 116700 21700 116800 21800
rect 116700 21800 116800 21900
rect 116700 21900 116800 22000
rect 116700 22000 116800 22100
rect 116700 22100 116800 22200
rect 116700 22200 116800 22300
rect 116700 22300 116800 22400
rect 116700 22400 116800 22500
rect 116700 22500 116800 22600
rect 116700 22600 116800 22700
rect 116700 22700 116800 22800
rect 116700 22800 116800 22900
rect 116700 22900 116800 23000
rect 116700 23900 116800 24000
rect 116700 24000 116800 24100
rect 116700 24100 116800 24200
rect 116700 24200 116800 24300
rect 116700 24300 116800 24400
rect 116700 24400 116800 24500
rect 116700 24500 116800 24600
rect 116700 24600 116800 24700
rect 116700 24700 116800 24800
rect 116700 24800 116800 24900
rect 116700 24900 116800 25000
rect 116700 25000 116800 25100
rect 116700 25100 116800 25200
rect 116700 25200 116800 25300
rect 116700 25300 116800 25400
rect 116700 25400 116800 25500
rect 116700 25500 116800 25600
rect 116700 25600 116800 25700
rect 116700 25700 116800 25800
rect 116700 25800 116800 25900
rect 116700 25900 116800 26000
rect 116700 26000 116800 26100
rect 116700 26100 116800 26200
rect 116700 26200 116800 26300
rect 116700 26300 116800 26400
rect 116700 26400 116800 26500
rect 116700 26500 116800 26600
rect 116700 26600 116800 26700
rect 116700 26700 116800 26800
rect 116700 26800 116800 26900
rect 116700 26900 116800 27000
rect 116700 27000 116800 27100
rect 116700 27100 116800 27200
rect 116700 27200 116800 27300
rect 116700 27300 116800 27400
rect 116700 27400 116800 27500
rect 116700 27500 116800 27600
rect 116700 27600 116800 27700
rect 116700 27700 116800 27800
rect 116700 27800 116800 27900
rect 116700 27900 116800 28000
rect 116800 20700 116900 20800
rect 116800 20800 116900 20900
rect 116800 20900 116900 21000
rect 116800 21000 116900 21100
rect 116800 21100 116900 21200
rect 116800 21200 116900 21300
rect 116800 21300 116900 21400
rect 116800 21400 116900 21500
rect 116800 21500 116900 21600
rect 116800 21600 116900 21700
rect 116800 21700 116900 21800
rect 116800 21800 116900 21900
rect 116800 21900 116900 22000
rect 116800 22000 116900 22100
rect 116800 22100 116900 22200
rect 116800 22200 116900 22300
rect 116800 22300 116900 22400
rect 116800 22400 116900 22500
rect 116800 22500 116900 22600
rect 116800 22600 116900 22700
rect 116800 22700 116900 22800
rect 116800 22800 116900 22900
rect 116800 23900 116900 24000
rect 116800 24000 116900 24100
rect 116800 24100 116900 24200
rect 116800 24200 116900 24300
rect 116800 24300 116900 24400
rect 116800 24400 116900 24500
rect 116800 24500 116900 24600
rect 116800 24600 116900 24700
rect 116800 24700 116900 24800
rect 116800 24800 116900 24900
rect 116800 24900 116900 25000
rect 116800 25000 116900 25100
rect 116800 25100 116900 25200
rect 116800 25200 116900 25300
rect 116800 25300 116900 25400
rect 116800 25400 116900 25500
rect 116800 25500 116900 25600
rect 116800 25600 116900 25700
rect 116800 25700 116900 25800
rect 116800 25800 116900 25900
rect 116800 25900 116900 26000
rect 116800 26000 116900 26100
rect 116800 26100 116900 26200
rect 116800 26200 116900 26300
rect 116800 26300 116900 26400
rect 116800 26400 116900 26500
rect 116800 26500 116900 26600
rect 116800 26600 116900 26700
rect 116800 26700 116900 26800
rect 116800 26800 116900 26900
rect 116800 26900 116900 27000
rect 116800 27000 116900 27100
rect 116800 27100 116900 27200
rect 116800 27200 116900 27300
rect 116800 27300 116900 27400
rect 116800 27400 116900 27500
rect 116800 27500 116900 27600
rect 116800 27600 116900 27700
rect 116900 20700 117000 20800
rect 116900 20800 117000 20900
rect 116900 20900 117000 21000
rect 116900 21000 117000 21100
rect 116900 21100 117000 21200
rect 116900 21200 117000 21300
rect 116900 21300 117000 21400
rect 116900 21400 117000 21500
rect 116900 21500 117000 21600
rect 116900 21600 117000 21700
rect 116900 21700 117000 21800
rect 116900 21800 117000 21900
rect 116900 21900 117000 22000
rect 116900 22000 117000 22100
rect 116900 22100 117000 22200
rect 116900 22200 117000 22300
rect 116900 22300 117000 22400
rect 116900 22400 117000 22500
rect 116900 22500 117000 22600
rect 116900 22600 117000 22700
rect 116900 22700 117000 22800
rect 116900 23900 117000 24000
rect 116900 24000 117000 24100
rect 116900 24100 117000 24200
rect 116900 24200 117000 24300
rect 116900 24300 117000 24400
rect 116900 24400 117000 24500
rect 116900 24500 117000 24600
rect 116900 24600 117000 24700
rect 116900 24700 117000 24800
rect 116900 24800 117000 24900
rect 116900 24900 117000 25000
rect 116900 25000 117000 25100
rect 116900 25100 117000 25200
rect 116900 25200 117000 25300
rect 116900 25300 117000 25400
rect 116900 25400 117000 25500
rect 116900 25500 117000 25600
rect 116900 25600 117000 25700
rect 116900 25700 117000 25800
rect 116900 25800 117000 25900
rect 116900 25900 117000 26000
rect 116900 26000 117000 26100
rect 116900 26100 117000 26200
rect 116900 26200 117000 26300
rect 116900 26300 117000 26400
rect 116900 26400 117000 26500
rect 116900 26500 117000 26600
rect 116900 26600 117000 26700
rect 116900 26700 117000 26800
rect 116900 26800 117000 26900
rect 116900 26900 117000 27000
rect 116900 27000 117000 27100
rect 116900 27100 117000 27200
rect 116900 27200 117000 27300
rect 116900 27300 117000 27400
rect 116900 27400 117000 27500
rect 117000 20700 117100 20800
rect 117000 20800 117100 20900
rect 117000 20900 117100 21000
rect 117000 21000 117100 21100
rect 117000 21100 117100 21200
rect 117000 21200 117100 21300
rect 117000 21300 117100 21400
rect 117000 21400 117100 21500
rect 117000 21500 117100 21600
rect 117000 21600 117100 21700
rect 117000 21700 117100 21800
rect 117000 21800 117100 21900
rect 117000 21900 117100 22000
rect 117000 22000 117100 22100
rect 117000 22100 117100 22200
rect 117000 22200 117100 22300
rect 117000 22300 117100 22400
rect 117000 22400 117100 22500
rect 117000 22500 117100 22600
rect 117000 22600 117100 22700
rect 117000 22700 117100 22800
rect 117000 23900 117100 24000
rect 117000 24000 117100 24100
rect 117000 24100 117100 24200
rect 117000 24200 117100 24300
rect 117000 24300 117100 24400
rect 117000 24400 117100 24500
rect 117000 24500 117100 24600
rect 117000 24600 117100 24700
rect 117000 24700 117100 24800
rect 117000 24800 117100 24900
rect 117000 24900 117100 25000
rect 117000 25000 117100 25100
rect 117000 25100 117100 25200
rect 117000 25200 117100 25300
rect 117000 25300 117100 25400
rect 117000 25400 117100 25500
rect 117000 25500 117100 25600
rect 117000 25600 117100 25700
rect 117000 25700 117100 25800
rect 117000 25800 117100 25900
rect 117000 25900 117100 26000
rect 117000 26000 117100 26100
rect 117000 26100 117100 26200
rect 117000 26200 117100 26300
rect 117000 26300 117100 26400
rect 117000 26400 117100 26500
rect 117000 26500 117100 26600
rect 117000 26600 117100 26700
rect 117000 26700 117100 26800
rect 117000 26800 117100 26900
rect 117000 26900 117100 27000
rect 117000 27000 117100 27100
rect 117000 27100 117100 27200
rect 117100 20700 117200 20800
rect 117100 20800 117200 20900
rect 117100 20900 117200 21000
rect 117100 21000 117200 21100
rect 117100 21100 117200 21200
rect 117100 21200 117200 21300
rect 117100 21300 117200 21400
rect 117100 21400 117200 21500
rect 117100 21500 117200 21600
rect 117100 21600 117200 21700
rect 117100 21700 117200 21800
rect 117100 21800 117200 21900
rect 117100 21900 117200 22000
rect 117100 22000 117200 22100
rect 117100 22100 117200 22200
rect 117100 22200 117200 22300
rect 117100 22300 117200 22400
rect 117100 22400 117200 22500
rect 117100 22500 117200 22600
rect 117100 22600 117200 22700
rect 117100 22700 117200 22800
rect 117100 23900 117200 24000
rect 117100 24000 117200 24100
rect 117100 24100 117200 24200
rect 117100 24200 117200 24300
rect 117100 24300 117200 24400
rect 117100 24400 117200 24500
rect 117100 24500 117200 24600
rect 117100 24600 117200 24700
rect 117100 24700 117200 24800
rect 117100 24800 117200 24900
rect 117100 24900 117200 25000
rect 117100 25000 117200 25100
rect 117100 25100 117200 25200
rect 117100 25200 117200 25300
rect 117100 25300 117200 25400
rect 117100 25400 117200 25500
rect 117100 25500 117200 25600
rect 117100 25600 117200 25700
rect 117100 25700 117200 25800
rect 117100 25800 117200 25900
rect 117100 25900 117200 26000
rect 117100 26000 117200 26100
rect 117100 26100 117200 26200
rect 117100 26200 117200 26300
rect 117100 26300 117200 26400
rect 117100 26400 117200 26500
rect 117100 26500 117200 26600
rect 117100 26600 117200 26700
rect 117100 26700 117200 26800
rect 117100 26800 117200 26900
rect 117100 26900 117200 27000
rect 117200 20800 117300 20900
rect 117200 20900 117300 21000
rect 117200 21000 117300 21100
rect 117200 21100 117300 21200
rect 117200 21200 117300 21300
rect 117200 21300 117300 21400
rect 117200 21400 117300 21500
rect 117200 21500 117300 21600
rect 117200 21600 117300 21700
rect 117200 21700 117300 21800
rect 117200 21800 117300 21900
rect 117200 21900 117300 22000
rect 117200 22000 117300 22100
rect 117200 22100 117300 22200
rect 117200 22200 117300 22300
rect 117200 22300 117300 22400
rect 117200 22400 117300 22500
rect 117200 22500 117300 22600
rect 117200 22600 117300 22700
rect 117200 23900 117300 24000
rect 117200 24000 117300 24100
rect 117200 24100 117300 24200
rect 117200 24200 117300 24300
rect 117200 24300 117300 24400
rect 117200 24400 117300 24500
rect 117200 24500 117300 24600
rect 117200 24600 117300 24700
rect 117200 24700 117300 24800
rect 117200 24800 117300 24900
rect 117200 24900 117300 25000
rect 117200 25000 117300 25100
rect 117200 25100 117300 25200
rect 117200 25200 117300 25300
rect 117200 25300 117300 25400
rect 117200 25400 117300 25500
rect 117200 25500 117300 25600
rect 117200 25600 117300 25700
rect 117200 25700 117300 25800
rect 117200 25800 117300 25900
rect 117200 25900 117300 26000
rect 117200 26000 117300 26100
rect 117200 26100 117300 26200
rect 117200 26200 117300 26300
rect 117200 26300 117300 26400
rect 117200 26400 117300 26500
rect 117200 26500 117300 26600
rect 117200 26600 117300 26700
rect 117200 26700 117300 26800
rect 117300 20800 117400 20900
rect 117300 20900 117400 21000
rect 117300 21000 117400 21100
rect 117300 21100 117400 21200
rect 117300 21200 117400 21300
rect 117300 21300 117400 21400
rect 117300 21400 117400 21500
rect 117300 21500 117400 21600
rect 117300 21600 117400 21700
rect 117300 21700 117400 21800
rect 117300 21800 117400 21900
rect 117300 21900 117400 22000
rect 117300 22000 117400 22100
rect 117300 22100 117400 22200
rect 117300 22200 117400 22300
rect 117300 22300 117400 22400
rect 117300 22400 117400 22500
rect 117300 22500 117400 22600
rect 117300 22600 117400 22700
rect 117300 23900 117400 24000
rect 117300 24000 117400 24100
rect 117300 24100 117400 24200
rect 117300 24200 117400 24300
rect 117300 24300 117400 24400
rect 117300 24400 117400 24500
rect 117300 24500 117400 24600
rect 117300 24600 117400 24700
rect 117300 24700 117400 24800
rect 117300 24800 117400 24900
rect 117300 24900 117400 25000
rect 117300 25000 117400 25100
rect 117300 25100 117400 25200
rect 117300 25200 117400 25300
rect 117300 25300 117400 25400
rect 117300 25400 117400 25500
rect 117300 25500 117400 25600
rect 117300 25600 117400 25700
rect 117300 25700 117400 25800
rect 117300 25800 117400 25900
rect 117300 25900 117400 26000
rect 117300 26000 117400 26100
rect 117300 26100 117400 26200
rect 117300 26200 117400 26300
rect 117300 26300 117400 26400
rect 117300 26400 117400 26500
rect 117300 26500 117400 26600
rect 117300 26600 117400 26700
rect 117400 20800 117500 20900
rect 117400 20900 117500 21000
rect 117400 21000 117500 21100
rect 117400 21100 117500 21200
rect 117400 21200 117500 21300
rect 117400 21300 117500 21400
rect 117400 21400 117500 21500
rect 117400 21500 117500 21600
rect 117400 21600 117500 21700
rect 117400 21700 117500 21800
rect 117400 21800 117500 21900
rect 117400 21900 117500 22000
rect 117400 22000 117500 22100
rect 117400 22100 117500 22200
rect 117400 22200 117500 22300
rect 117400 22300 117500 22400
rect 117400 22400 117500 22500
rect 117400 22500 117500 22600
rect 117400 22600 117500 22700
rect 117400 23900 117500 24000
rect 117400 24000 117500 24100
rect 117400 24100 117500 24200
rect 117400 24200 117500 24300
rect 117400 24300 117500 24400
rect 117400 24400 117500 24500
rect 117400 24500 117500 24600
rect 117400 24600 117500 24700
rect 117400 24700 117500 24800
rect 117400 24800 117500 24900
rect 117400 24900 117500 25000
rect 117400 25000 117500 25100
rect 117400 25100 117500 25200
rect 117400 25200 117500 25300
rect 117400 25300 117500 25400
rect 117400 25400 117500 25500
rect 117400 25500 117500 25600
rect 117400 25600 117500 25700
rect 117400 25700 117500 25800
rect 117400 25800 117500 25900
rect 117400 25900 117500 26000
rect 117400 26000 117500 26100
rect 117400 26100 117500 26200
rect 117400 26200 117500 26300
rect 117400 26300 117500 26400
rect 117400 26400 117500 26500
rect 117500 20800 117600 20900
rect 117500 20900 117600 21000
rect 117500 21000 117600 21100
rect 117500 21100 117600 21200
rect 117500 21200 117600 21300
rect 117500 21300 117600 21400
rect 117500 21400 117600 21500
rect 117500 21500 117600 21600
rect 117500 21600 117600 21700
rect 117500 21700 117600 21800
rect 117500 21800 117600 21900
rect 117500 21900 117600 22000
rect 117500 22000 117600 22100
rect 117500 22100 117600 22200
rect 117500 22200 117600 22300
rect 117500 22300 117600 22400
rect 117500 22400 117600 22500
rect 117500 22500 117600 22600
rect 117500 22600 117600 22700
rect 117500 22700 117600 22800
rect 117500 23800 117600 23900
rect 117500 23900 117600 24000
rect 117500 24000 117600 24100
rect 117500 24100 117600 24200
rect 117500 24200 117600 24300
rect 117500 24300 117600 24400
rect 117500 24400 117600 24500
rect 117500 24500 117600 24600
rect 117500 24600 117600 24700
rect 117500 24700 117600 24800
rect 117500 24800 117600 24900
rect 117500 24900 117600 25000
rect 117500 25000 117600 25100
rect 117500 25100 117600 25200
rect 117500 25200 117600 25300
rect 117500 25300 117600 25400
rect 117500 25400 117600 25500
rect 117500 25500 117600 25600
rect 117500 25600 117600 25700
rect 117500 25700 117600 25800
rect 117500 25800 117600 25900
rect 117500 25900 117600 26000
rect 117500 26000 117600 26100
rect 117500 26100 117600 26200
rect 117500 26200 117600 26300
rect 117500 26300 117600 26400
rect 117600 20900 117700 21000
rect 117600 21000 117700 21100
rect 117600 21100 117700 21200
rect 117600 21200 117700 21300
rect 117600 21300 117700 21400
rect 117600 21400 117700 21500
rect 117600 21500 117700 21600
rect 117600 21600 117700 21700
rect 117600 21700 117700 21800
rect 117600 21800 117700 21900
rect 117600 21900 117700 22000
rect 117600 22000 117700 22100
rect 117600 22100 117700 22200
rect 117600 22200 117700 22300
rect 117600 22300 117700 22400
rect 117600 22400 117700 22500
rect 117600 22500 117700 22600
rect 117600 22600 117700 22700
rect 117600 22700 117700 22800
rect 117600 23800 117700 23900
rect 117600 23900 117700 24000
rect 117600 24000 117700 24100
rect 117600 24100 117700 24200
rect 117600 24200 117700 24300
rect 117600 24300 117700 24400
rect 117600 24400 117700 24500
rect 117600 24500 117700 24600
rect 117600 24600 117700 24700
rect 117600 24700 117700 24800
rect 117600 24800 117700 24900
rect 117600 24900 117700 25000
rect 117600 25000 117700 25100
rect 117600 25100 117700 25200
rect 117600 25200 117700 25300
rect 117600 25300 117700 25400
rect 117600 25400 117700 25500
rect 117600 25500 117700 25600
rect 117600 25600 117700 25700
rect 117600 25700 117700 25800
rect 117600 25800 117700 25900
rect 117600 25900 117700 26000
rect 117600 26000 117700 26100
rect 117600 26100 117700 26200
rect 117600 26200 117700 26300
rect 117700 20900 117800 21000
rect 117700 21000 117800 21100
rect 117700 21100 117800 21200
rect 117700 21200 117800 21300
rect 117700 21300 117800 21400
rect 117700 21400 117800 21500
rect 117700 21500 117800 21600
rect 117700 21600 117800 21700
rect 117700 21700 117800 21800
rect 117700 21800 117800 21900
rect 117700 21900 117800 22000
rect 117700 22000 117800 22100
rect 117700 22100 117800 22200
rect 117700 22200 117800 22300
rect 117700 22300 117800 22400
rect 117700 22400 117800 22500
rect 117700 22500 117800 22600
rect 117700 22600 117800 22700
rect 117700 22700 117800 22800
rect 117700 23700 117800 23800
rect 117700 23800 117800 23900
rect 117700 23900 117800 24000
rect 117700 24000 117800 24100
rect 117700 24100 117800 24200
rect 117700 24200 117800 24300
rect 117700 24300 117800 24400
rect 117700 24400 117800 24500
rect 117700 24500 117800 24600
rect 117700 24600 117800 24700
rect 117700 24700 117800 24800
rect 117700 24800 117800 24900
rect 117700 24900 117800 25000
rect 117700 25000 117800 25100
rect 117700 25100 117800 25200
rect 117700 25200 117800 25300
rect 117700 25300 117800 25400
rect 117700 25400 117800 25500
rect 117700 25500 117800 25600
rect 117700 25600 117800 25700
rect 117700 25700 117800 25800
rect 117700 25800 117800 25900
rect 117700 25900 117800 26000
rect 117700 26000 117800 26100
rect 117700 26100 117800 26200
rect 117800 20900 117900 21000
rect 117800 21000 117900 21100
rect 117800 21100 117900 21200
rect 117800 21200 117900 21300
rect 117800 21300 117900 21400
rect 117800 21400 117900 21500
rect 117800 21500 117900 21600
rect 117800 21600 117900 21700
rect 117800 21700 117900 21800
rect 117800 21800 117900 21900
rect 117800 21900 117900 22000
rect 117800 22000 117900 22100
rect 117800 22100 117900 22200
rect 117800 22200 117900 22300
rect 117800 22300 117900 22400
rect 117800 22400 117900 22500
rect 117800 22500 117900 22600
rect 117800 22600 117900 22700
rect 117800 22700 117900 22800
rect 117800 22800 117900 22900
rect 117800 22900 117900 23000
rect 117800 23600 117900 23700
rect 117800 23700 117900 23800
rect 117800 23800 117900 23900
rect 117800 23900 117900 24000
rect 117800 24000 117900 24100
rect 117800 24100 117900 24200
rect 117800 24200 117900 24300
rect 117800 24300 117900 24400
rect 117800 24400 117900 24500
rect 117800 24500 117900 24600
rect 117800 24600 117900 24700
rect 117800 24700 117900 24800
rect 117800 24800 117900 24900
rect 117800 24900 117900 25000
rect 117800 25000 117900 25100
rect 117800 25100 117900 25200
rect 117800 25200 117900 25300
rect 117800 25300 117900 25400
rect 117800 25400 117900 25500
rect 117800 25500 117900 25600
rect 117800 25600 117900 25700
rect 117800 25700 117900 25800
rect 117800 25800 117900 25900
rect 117800 25900 117900 26000
rect 117800 26000 117900 26100
rect 117900 21000 118000 21100
rect 117900 21100 118000 21200
rect 117900 21200 118000 21300
rect 117900 21300 118000 21400
rect 117900 21400 118000 21500
rect 117900 21500 118000 21600
rect 117900 21600 118000 21700
rect 117900 21700 118000 21800
rect 117900 21800 118000 21900
rect 117900 21900 118000 22000
rect 117900 22000 118000 22100
rect 117900 22100 118000 22200
rect 117900 22200 118000 22300
rect 117900 22300 118000 22400
rect 117900 22400 118000 22500
rect 117900 22500 118000 22600
rect 117900 22600 118000 22700
rect 117900 22700 118000 22800
rect 117900 22800 118000 22900
rect 117900 22900 118000 23000
rect 117900 23000 118000 23100
rect 117900 23100 118000 23200
rect 117900 23200 118000 23300
rect 117900 23300 118000 23400
rect 117900 23400 118000 23500
rect 117900 23500 118000 23600
rect 117900 23600 118000 23700
rect 117900 23700 118000 23800
rect 117900 23800 118000 23900
rect 117900 23900 118000 24000
rect 117900 24000 118000 24100
rect 117900 24100 118000 24200
rect 117900 24200 118000 24300
rect 117900 24300 118000 24400
rect 117900 24400 118000 24500
rect 117900 24500 118000 24600
rect 117900 24600 118000 24700
rect 117900 24700 118000 24800
rect 117900 24800 118000 24900
rect 117900 24900 118000 25000
rect 117900 25000 118000 25100
rect 117900 25100 118000 25200
rect 117900 25200 118000 25300
rect 117900 25300 118000 25400
rect 117900 25400 118000 25500
rect 117900 25500 118000 25600
rect 117900 25600 118000 25700
rect 117900 25700 118000 25800
rect 117900 25800 118000 25900
rect 117900 25900 118000 26000
rect 118000 21000 118100 21100
rect 118000 21100 118100 21200
rect 118000 21200 118100 21300
rect 118000 21300 118100 21400
rect 118000 21400 118100 21500
rect 118000 21500 118100 21600
rect 118000 21600 118100 21700
rect 118000 21700 118100 21800
rect 118000 21800 118100 21900
rect 118000 21900 118100 22000
rect 118000 22000 118100 22100
rect 118000 22100 118100 22200
rect 118000 22200 118100 22300
rect 118000 22300 118100 22400
rect 118000 22400 118100 22500
rect 118000 22500 118100 22600
rect 118000 22600 118100 22700
rect 118000 22700 118100 22800
rect 118000 22800 118100 22900
rect 118000 22900 118100 23000
rect 118000 23000 118100 23100
rect 118000 23100 118100 23200
rect 118000 23200 118100 23300
rect 118000 23300 118100 23400
rect 118000 23400 118100 23500
rect 118000 23500 118100 23600
rect 118000 23600 118100 23700
rect 118000 23700 118100 23800
rect 118000 23800 118100 23900
rect 118000 23900 118100 24000
rect 118000 24000 118100 24100
rect 118000 24100 118100 24200
rect 118000 24200 118100 24300
rect 118000 24300 118100 24400
rect 118000 24400 118100 24500
rect 118000 24500 118100 24600
rect 118000 24600 118100 24700
rect 118000 24700 118100 24800
rect 118000 24800 118100 24900
rect 118000 24900 118100 25000
rect 118000 25000 118100 25100
rect 118000 25100 118100 25200
rect 118000 25200 118100 25300
rect 118000 25300 118100 25400
rect 118000 25400 118100 25500
rect 118000 25500 118100 25600
rect 118000 25600 118100 25700
rect 118000 25700 118100 25800
rect 118000 25800 118100 25900
rect 118000 25900 118100 26000
rect 118100 21100 118200 21200
rect 118100 21200 118200 21300
rect 118100 21300 118200 21400
rect 118100 21400 118200 21500
rect 118100 21500 118200 21600
rect 118100 21600 118200 21700
rect 118100 21700 118200 21800
rect 118100 21800 118200 21900
rect 118100 21900 118200 22000
rect 118100 22000 118200 22100
rect 118100 22100 118200 22200
rect 118100 22200 118200 22300
rect 118100 22300 118200 22400
rect 118100 22400 118200 22500
rect 118100 22500 118200 22600
rect 118100 22600 118200 22700
rect 118100 22700 118200 22800
rect 118100 22800 118200 22900
rect 118100 22900 118200 23000
rect 118100 23000 118200 23100
rect 118100 23100 118200 23200
rect 118100 23200 118200 23300
rect 118100 23300 118200 23400
rect 118100 23400 118200 23500
rect 118100 23500 118200 23600
rect 118100 23600 118200 23700
rect 118100 23700 118200 23800
rect 118100 23800 118200 23900
rect 118100 23900 118200 24000
rect 118100 24000 118200 24100
rect 118100 24100 118200 24200
rect 118100 24200 118200 24300
rect 118100 24300 118200 24400
rect 118100 24400 118200 24500
rect 118100 24500 118200 24600
rect 118100 24600 118200 24700
rect 118100 24700 118200 24800
rect 118100 24800 118200 24900
rect 118100 24900 118200 25000
rect 118100 25000 118200 25100
rect 118100 25100 118200 25200
rect 118100 25200 118200 25300
rect 118100 25300 118200 25400
rect 118100 25400 118200 25500
rect 118100 25500 118200 25600
rect 118100 25600 118200 25700
rect 118100 25700 118200 25800
rect 118100 25800 118200 25900
rect 118100 25900 118200 26000
rect 118200 21100 118300 21200
rect 118200 21200 118300 21300
rect 118200 21300 118300 21400
rect 118200 21400 118300 21500
rect 118200 21500 118300 21600
rect 118200 21600 118300 21700
rect 118200 21700 118300 21800
rect 118200 21800 118300 21900
rect 118200 21900 118300 22000
rect 118200 22000 118300 22100
rect 118200 22100 118300 22200
rect 118200 22200 118300 22300
rect 118200 22300 118300 22400
rect 118200 22400 118300 22500
rect 118200 22500 118300 22600
rect 118200 22600 118300 22700
rect 118200 22700 118300 22800
rect 118200 22800 118300 22900
rect 118200 22900 118300 23000
rect 118200 23000 118300 23100
rect 118200 23100 118300 23200
rect 118200 23200 118300 23300
rect 118200 23300 118300 23400
rect 118200 23400 118300 23500
rect 118200 23500 118300 23600
rect 118200 23600 118300 23700
rect 118200 23700 118300 23800
rect 118200 23800 118300 23900
rect 118200 23900 118300 24000
rect 118200 24000 118300 24100
rect 118200 24100 118300 24200
rect 118200 24200 118300 24300
rect 118200 24300 118300 24400
rect 118200 24400 118300 24500
rect 118200 24500 118300 24600
rect 118200 24600 118300 24700
rect 118200 24700 118300 24800
rect 118200 24800 118300 24900
rect 118200 24900 118300 25000
rect 118200 25000 118300 25100
rect 118200 25100 118300 25200
rect 118200 25200 118300 25300
rect 118200 25300 118300 25400
rect 118200 25400 118300 25500
rect 118200 25500 118300 25600
rect 118200 25600 118300 25700
rect 118200 25700 118300 25800
rect 118200 25800 118300 25900
rect 118200 25900 118300 26000
rect 118200 26000 118300 26100
rect 118300 21200 118400 21300
rect 118300 21300 118400 21400
rect 118300 21400 118400 21500
rect 118300 21500 118400 21600
rect 118300 21600 118400 21700
rect 118300 21700 118400 21800
rect 118300 21800 118400 21900
rect 118300 21900 118400 22000
rect 118300 22000 118400 22100
rect 118300 22100 118400 22200
rect 118300 22200 118400 22300
rect 118300 22300 118400 22400
rect 118300 22400 118400 22500
rect 118300 22500 118400 22600
rect 118300 22600 118400 22700
rect 118300 22700 118400 22800
rect 118300 22800 118400 22900
rect 118300 22900 118400 23000
rect 118300 23000 118400 23100
rect 118300 23100 118400 23200
rect 118300 23200 118400 23300
rect 118300 23300 118400 23400
rect 118300 23400 118400 23500
rect 118300 23500 118400 23600
rect 118300 23600 118400 23700
rect 118300 23700 118400 23800
rect 118300 23800 118400 23900
rect 118300 23900 118400 24000
rect 118300 24000 118400 24100
rect 118300 24100 118400 24200
rect 118300 24200 118400 24300
rect 118300 24300 118400 24400
rect 118300 24400 118400 24500
rect 118300 24500 118400 24600
rect 118300 24600 118400 24700
rect 118300 24700 118400 24800
rect 118300 24800 118400 24900
rect 118300 24900 118400 25000
rect 118300 25000 118400 25100
rect 118300 25100 118400 25200
rect 118300 25200 118400 25300
rect 118300 25300 118400 25400
rect 118300 25400 118400 25500
rect 118300 25500 118400 25600
rect 118300 25600 118400 25700
rect 118300 25700 118400 25800
rect 118300 25800 118400 25900
rect 118300 25900 118400 26000
rect 118300 26000 118400 26100
rect 118400 21300 118500 21400
rect 118400 21400 118500 21500
rect 118400 21500 118500 21600
rect 118400 21600 118500 21700
rect 118400 21700 118500 21800
rect 118400 21800 118500 21900
rect 118400 21900 118500 22000
rect 118400 22000 118500 22100
rect 118400 22100 118500 22200
rect 118400 22200 118500 22300
rect 118400 22300 118500 22400
rect 118400 22400 118500 22500
rect 118400 22500 118500 22600
rect 118400 22600 118500 22700
rect 118400 22700 118500 22800
rect 118400 22800 118500 22900
rect 118400 22900 118500 23000
rect 118400 23000 118500 23100
rect 118400 23100 118500 23200
rect 118400 23200 118500 23300
rect 118400 23300 118500 23400
rect 118400 23400 118500 23500
rect 118400 23500 118500 23600
rect 118400 23600 118500 23700
rect 118400 23700 118500 23800
rect 118400 23800 118500 23900
rect 118400 23900 118500 24000
rect 118400 24000 118500 24100
rect 118400 24100 118500 24200
rect 118400 24200 118500 24300
rect 118400 24300 118500 24400
rect 118400 24400 118500 24500
rect 118400 24500 118500 24600
rect 118400 24600 118500 24700
rect 118400 24700 118500 24800
rect 118400 24800 118500 24900
rect 118400 24900 118500 25000
rect 118400 25000 118500 25100
rect 118400 25100 118500 25200
rect 118400 25200 118500 25300
rect 118400 25300 118500 25400
rect 118400 25400 118500 25500
rect 118400 25500 118500 25600
rect 118400 25600 118500 25700
rect 118400 25700 118500 25800
rect 118400 25800 118500 25900
rect 118400 25900 118500 26000
rect 118400 26000 118500 26100
rect 118400 26100 118500 26200
rect 118500 21300 118600 21400
rect 118500 21400 118600 21500
rect 118500 21500 118600 21600
rect 118500 21600 118600 21700
rect 118500 21700 118600 21800
rect 118500 21800 118600 21900
rect 118500 21900 118600 22000
rect 118500 22000 118600 22100
rect 118500 22100 118600 22200
rect 118500 22200 118600 22300
rect 118500 22300 118600 22400
rect 118500 22400 118600 22500
rect 118500 22500 118600 22600
rect 118500 22600 118600 22700
rect 118500 22700 118600 22800
rect 118500 22800 118600 22900
rect 118500 22900 118600 23000
rect 118500 23000 118600 23100
rect 118500 23100 118600 23200
rect 118500 23200 118600 23300
rect 118500 23300 118600 23400
rect 118500 23400 118600 23500
rect 118500 23500 118600 23600
rect 118500 23600 118600 23700
rect 118500 23700 118600 23800
rect 118500 23800 118600 23900
rect 118500 23900 118600 24000
rect 118500 24000 118600 24100
rect 118500 24100 118600 24200
rect 118500 24200 118600 24300
rect 118500 24300 118600 24400
rect 118500 24400 118600 24500
rect 118500 24500 118600 24600
rect 118500 24600 118600 24700
rect 118500 24700 118600 24800
rect 118500 24800 118600 24900
rect 118500 24900 118600 25000
rect 118500 25000 118600 25100
rect 118500 25100 118600 25200
rect 118500 25200 118600 25300
rect 118500 25300 118600 25400
rect 118500 25400 118600 25500
rect 118500 25500 118600 25600
rect 118500 25600 118600 25700
rect 118500 25700 118600 25800
rect 118500 25800 118600 25900
rect 118500 25900 118600 26000
rect 118500 26000 118600 26100
rect 118500 26100 118600 26200
rect 118500 26200 118600 26300
rect 118600 21400 118700 21500
rect 118600 21500 118700 21600
rect 118600 21600 118700 21700
rect 118600 21700 118700 21800
rect 118600 21800 118700 21900
rect 118600 21900 118700 22000
rect 118600 22000 118700 22100
rect 118600 22100 118700 22200
rect 118600 22200 118700 22300
rect 118600 22300 118700 22400
rect 118600 22400 118700 22500
rect 118600 22500 118700 22600
rect 118600 22600 118700 22700
rect 118600 22700 118700 22800
rect 118600 22800 118700 22900
rect 118600 22900 118700 23000
rect 118600 23000 118700 23100
rect 118600 23100 118700 23200
rect 118600 23200 118700 23300
rect 118600 23300 118700 23400
rect 118600 23400 118700 23500
rect 118600 23500 118700 23600
rect 118600 23600 118700 23700
rect 118600 23700 118700 23800
rect 118600 23800 118700 23900
rect 118600 23900 118700 24000
rect 118600 24000 118700 24100
rect 118600 24100 118700 24200
rect 118600 24200 118700 24300
rect 118600 24300 118700 24400
rect 118600 24400 118700 24500
rect 118600 24500 118700 24600
rect 118600 24600 118700 24700
rect 118600 24700 118700 24800
rect 118600 24800 118700 24900
rect 118600 24900 118700 25000
rect 118600 25000 118700 25100
rect 118600 25100 118700 25200
rect 118600 25200 118700 25300
rect 118600 25300 118700 25400
rect 118600 25400 118700 25500
rect 118600 25500 118700 25600
rect 118600 25600 118700 25700
rect 118600 25700 118700 25800
rect 118600 25800 118700 25900
rect 118600 25900 118700 26000
rect 118600 26000 118700 26100
rect 118600 26100 118700 26200
rect 118600 26200 118700 26300
rect 118600 26300 118700 26400
rect 118700 21500 118800 21600
rect 118700 21600 118800 21700
rect 118700 21700 118800 21800
rect 118700 21800 118800 21900
rect 118700 21900 118800 22000
rect 118700 22000 118800 22100
rect 118700 22100 118800 22200
rect 118700 22200 118800 22300
rect 118700 22300 118800 22400
rect 118700 22400 118800 22500
rect 118700 22500 118800 22600
rect 118700 22600 118800 22700
rect 118700 22700 118800 22800
rect 118700 22800 118800 22900
rect 118700 22900 118800 23000
rect 118700 23000 118800 23100
rect 118700 23100 118800 23200
rect 118700 23200 118800 23300
rect 118700 23300 118800 23400
rect 118700 23400 118800 23500
rect 118700 23500 118800 23600
rect 118700 23600 118800 23700
rect 118700 23700 118800 23800
rect 118700 23800 118800 23900
rect 118700 23900 118800 24000
rect 118700 24000 118800 24100
rect 118700 24100 118800 24200
rect 118700 24200 118800 24300
rect 118700 24300 118800 24400
rect 118700 24400 118800 24500
rect 118700 24500 118800 24600
rect 118700 24600 118800 24700
rect 118700 24700 118800 24800
rect 118700 24800 118800 24900
rect 118700 24900 118800 25000
rect 118700 25000 118800 25100
rect 118700 25100 118800 25200
rect 118700 25200 118800 25300
rect 118700 25300 118800 25400
rect 118700 25400 118800 25500
rect 118700 25500 118800 25600
rect 118700 25600 118800 25700
rect 118700 25700 118800 25800
rect 118700 25800 118800 25900
rect 118700 25900 118800 26000
rect 118700 26000 118800 26100
rect 118700 26100 118800 26200
rect 118700 26200 118800 26300
rect 118700 26300 118800 26400
rect 118700 26400 118800 26500
rect 118800 21600 118900 21700
rect 118800 21700 118900 21800
rect 118800 21800 118900 21900
rect 118800 21900 118900 22000
rect 118800 22000 118900 22100
rect 118800 22100 118900 22200
rect 118800 22200 118900 22300
rect 118800 22300 118900 22400
rect 118800 22400 118900 22500
rect 118800 22500 118900 22600
rect 118800 22600 118900 22700
rect 118800 22700 118900 22800
rect 118800 22800 118900 22900
rect 118800 22900 118900 23000
rect 118800 23000 118900 23100
rect 118800 23100 118900 23200
rect 118800 23200 118900 23300
rect 118800 23300 118900 23400
rect 118800 23400 118900 23500
rect 118800 23500 118900 23600
rect 118800 23600 118900 23700
rect 118800 23700 118900 23800
rect 118800 23800 118900 23900
rect 118800 23900 118900 24000
rect 118800 24000 118900 24100
rect 118800 24100 118900 24200
rect 118800 24200 118900 24300
rect 118800 24300 118900 24400
rect 118800 24400 118900 24500
rect 118800 24500 118900 24600
rect 118800 24600 118900 24700
rect 118800 24700 118900 24800
rect 118800 24800 118900 24900
rect 118800 24900 118900 25000
rect 118800 25000 118900 25100
rect 118800 25100 118900 25200
rect 118800 25200 118900 25300
rect 118800 25300 118900 25400
rect 118800 25400 118900 25500
rect 118800 25500 118900 25600
rect 118800 25600 118900 25700
rect 118800 25700 118900 25800
rect 118800 25800 118900 25900
rect 118800 25900 118900 26000
rect 118800 26000 118900 26100
rect 118800 26100 118900 26200
rect 118800 26200 118900 26300
rect 118800 26300 118900 26400
rect 118800 26400 118900 26500
rect 118800 26500 118900 26600
rect 118900 21700 119000 21800
rect 118900 21800 119000 21900
rect 118900 21900 119000 22000
rect 118900 22000 119000 22100
rect 118900 22100 119000 22200
rect 118900 22200 119000 22300
rect 118900 22300 119000 22400
rect 118900 22400 119000 22500
rect 118900 22500 119000 22600
rect 118900 22600 119000 22700
rect 118900 22700 119000 22800
rect 118900 22800 119000 22900
rect 118900 22900 119000 23000
rect 118900 23000 119000 23100
rect 118900 23100 119000 23200
rect 118900 23200 119000 23300
rect 118900 23300 119000 23400
rect 118900 23400 119000 23500
rect 118900 23500 119000 23600
rect 118900 23600 119000 23700
rect 118900 23700 119000 23800
rect 118900 23800 119000 23900
rect 118900 23900 119000 24000
rect 118900 24000 119000 24100
rect 118900 24100 119000 24200
rect 118900 24200 119000 24300
rect 118900 24300 119000 24400
rect 118900 24400 119000 24500
rect 118900 24500 119000 24600
rect 118900 24600 119000 24700
rect 118900 24700 119000 24800
rect 118900 24800 119000 24900
rect 118900 24900 119000 25000
rect 118900 25000 119000 25100
rect 118900 25100 119000 25200
rect 118900 25200 119000 25300
rect 118900 25300 119000 25400
rect 118900 25400 119000 25500
rect 118900 25500 119000 25600
rect 118900 25600 119000 25700
rect 118900 25700 119000 25800
rect 118900 25800 119000 25900
rect 118900 25900 119000 26000
rect 118900 26000 119000 26100
rect 118900 26100 119000 26200
rect 118900 26200 119000 26300
rect 118900 26300 119000 26400
rect 118900 26400 119000 26500
rect 118900 26500 119000 26600
rect 118900 26600 119000 26700
rect 119000 21800 119100 21900
rect 119000 21900 119100 22000
rect 119000 22000 119100 22100
rect 119000 22100 119100 22200
rect 119000 22200 119100 22300
rect 119000 22300 119100 22400
rect 119000 22400 119100 22500
rect 119000 22500 119100 22600
rect 119000 22600 119100 22700
rect 119000 22700 119100 22800
rect 119000 22800 119100 22900
rect 119000 22900 119100 23000
rect 119000 23000 119100 23100
rect 119000 23100 119100 23200
rect 119000 23200 119100 23300
rect 119000 23300 119100 23400
rect 119000 23400 119100 23500
rect 119000 23500 119100 23600
rect 119000 23600 119100 23700
rect 119000 23700 119100 23800
rect 119000 23800 119100 23900
rect 119000 23900 119100 24000
rect 119000 24000 119100 24100
rect 119000 24100 119100 24200
rect 119000 24200 119100 24300
rect 119000 24300 119100 24400
rect 119000 24400 119100 24500
rect 119000 24500 119100 24600
rect 119000 24600 119100 24700
rect 119000 24700 119100 24800
rect 119000 24800 119100 24900
rect 119000 24900 119100 25000
rect 119000 25000 119100 25100
rect 119000 25100 119100 25200
rect 119000 25200 119100 25300
rect 119000 25300 119100 25400
rect 119000 25400 119100 25500
rect 119000 25500 119100 25600
rect 119000 25600 119100 25700
rect 119000 25700 119100 25800
rect 119000 25800 119100 25900
rect 119000 25900 119100 26000
rect 119000 26000 119100 26100
rect 119000 26100 119100 26200
rect 119000 26200 119100 26300
rect 119000 26300 119100 26400
rect 119000 26400 119100 26500
rect 119000 26500 119100 26600
rect 119000 26600 119100 26700
rect 119000 26700 119100 26800
rect 119100 21900 119200 22000
rect 119100 22000 119200 22100
rect 119100 22100 119200 22200
rect 119100 22200 119200 22300
rect 119100 22300 119200 22400
rect 119100 22400 119200 22500
rect 119100 22500 119200 22600
rect 119100 22600 119200 22700
rect 119100 22700 119200 22800
rect 119100 22800 119200 22900
rect 119100 22900 119200 23000
rect 119100 23000 119200 23100
rect 119100 23100 119200 23200
rect 119100 23200 119200 23300
rect 119100 23300 119200 23400
rect 119100 23400 119200 23500
rect 119100 23500 119200 23600
rect 119100 23600 119200 23700
rect 119100 23700 119200 23800
rect 119100 23800 119200 23900
rect 119100 23900 119200 24000
rect 119100 24000 119200 24100
rect 119100 24100 119200 24200
rect 119100 24200 119200 24300
rect 119100 24300 119200 24400
rect 119100 24400 119200 24500
rect 119100 24500 119200 24600
rect 119100 24600 119200 24700
rect 119100 24700 119200 24800
rect 119100 24800 119200 24900
rect 119100 24900 119200 25000
rect 119100 25000 119200 25100
rect 119100 25100 119200 25200
rect 119100 25200 119200 25300
rect 119100 25300 119200 25400
rect 119100 25400 119200 25500
rect 119100 25500 119200 25600
rect 119100 25600 119200 25700
rect 119100 25700 119200 25800
rect 119100 25800 119200 25900
rect 119100 25900 119200 26000
rect 119100 26000 119200 26100
rect 119100 26100 119200 26200
rect 119100 26200 119200 26300
rect 119100 26300 119200 26400
rect 119100 26400 119200 26500
rect 119100 26500 119200 26600
rect 119100 26600 119200 26700
rect 119100 26700 119200 26800
rect 119100 26800 119200 26900
rect 119200 22000 119300 22100
rect 119200 22100 119300 22200
rect 119200 22200 119300 22300
rect 119200 22300 119300 22400
rect 119200 22400 119300 22500
rect 119200 22500 119300 22600
rect 119200 22600 119300 22700
rect 119200 22700 119300 22800
rect 119200 22800 119300 22900
rect 119200 22900 119300 23000
rect 119200 23000 119300 23100
rect 119200 23100 119300 23200
rect 119200 23200 119300 23300
rect 119200 23300 119300 23400
rect 119200 23400 119300 23500
rect 119200 23500 119300 23600
rect 119200 23600 119300 23700
rect 119200 23700 119300 23800
rect 119200 23800 119300 23900
rect 119200 23900 119300 24000
rect 119200 24000 119300 24100
rect 119200 24100 119300 24200
rect 119200 24200 119300 24300
rect 119200 24300 119300 24400
rect 119200 24400 119300 24500
rect 119200 24500 119300 24600
rect 119200 24600 119300 24700
rect 119200 24700 119300 24800
rect 119200 24800 119300 24900
rect 119200 24900 119300 25000
rect 119200 25000 119300 25100
rect 119200 25100 119300 25200
rect 119200 25200 119300 25300
rect 119200 25300 119300 25400
rect 119200 25400 119300 25500
rect 119200 25500 119300 25600
rect 119200 25600 119300 25700
rect 119200 25700 119300 25800
rect 119200 25800 119300 25900
rect 119200 25900 119300 26000
rect 119200 26000 119300 26100
rect 119200 26100 119300 26200
rect 119200 26200 119300 26300
rect 119200 26300 119300 26400
rect 119200 26400 119300 26500
rect 119200 26500 119300 26600
rect 119200 26600 119300 26700
rect 119200 26700 119300 26800
rect 119200 26800 119300 26900
rect 119200 26900 119300 27000
rect 119300 22200 119400 22300
rect 119300 22300 119400 22400
rect 119300 22400 119400 22500
rect 119300 22500 119400 22600
rect 119300 22600 119400 22700
rect 119300 22700 119400 22800
rect 119300 22800 119400 22900
rect 119300 22900 119400 23000
rect 119300 23000 119400 23100
rect 119300 23100 119400 23200
rect 119300 23200 119400 23300
rect 119300 23300 119400 23400
rect 119300 23400 119400 23500
rect 119300 23500 119400 23600
rect 119300 23600 119400 23700
rect 119300 23700 119400 23800
rect 119300 23800 119400 23900
rect 119300 23900 119400 24000
rect 119300 24000 119400 24100
rect 119300 24100 119400 24200
rect 119300 24200 119400 24300
rect 119300 24300 119400 24400
rect 119300 24400 119400 24500
rect 119300 24500 119400 24600
rect 119300 24600 119400 24700
rect 119300 24700 119400 24800
rect 119300 24800 119400 24900
rect 119300 24900 119400 25000
rect 119300 25000 119400 25100
rect 119300 25100 119400 25200
rect 119300 25200 119400 25300
rect 119300 25300 119400 25400
rect 119300 25400 119400 25500
rect 119300 25500 119400 25600
rect 119300 25600 119400 25700
rect 119300 25700 119400 25800
rect 119300 25800 119400 25900
rect 119300 25900 119400 26000
rect 119300 26000 119400 26100
rect 119300 26100 119400 26200
rect 119300 26200 119400 26300
rect 119300 26300 119400 26400
rect 119300 26400 119400 26500
rect 119300 26500 119400 26600
rect 119300 26600 119400 26700
rect 119300 26700 119400 26800
rect 119300 26800 119400 26900
rect 119300 26900 119400 27000
rect 119300 27000 119400 27100
rect 119400 22300 119500 22400
rect 119400 22400 119500 22500
rect 119400 22500 119500 22600
rect 119400 22600 119500 22700
rect 119400 22700 119500 22800
rect 119400 22800 119500 22900
rect 119400 22900 119500 23000
rect 119400 23000 119500 23100
rect 119400 23100 119500 23200
rect 119400 23200 119500 23300
rect 119400 23300 119500 23400
rect 119400 23400 119500 23500
rect 119400 23500 119500 23600
rect 119400 23600 119500 23700
rect 119400 23700 119500 23800
rect 119400 23800 119500 23900
rect 119400 23900 119500 24000
rect 119400 24000 119500 24100
rect 119400 24100 119500 24200
rect 119400 24200 119500 24300
rect 119400 24300 119500 24400
rect 119400 24400 119500 24500
rect 119400 24500 119500 24600
rect 119400 24600 119500 24700
rect 119400 24700 119500 24800
rect 119400 24800 119500 24900
rect 119400 24900 119500 25000
rect 119400 25000 119500 25100
rect 119400 25100 119500 25200
rect 119400 25200 119500 25300
rect 119400 25300 119500 25400
rect 119400 25400 119500 25500
rect 119400 25500 119500 25600
rect 119400 25600 119500 25700
rect 119400 25700 119500 25800
rect 119400 25800 119500 25900
rect 119400 25900 119500 26000
rect 119400 26000 119500 26100
rect 119400 26100 119500 26200
rect 119400 26200 119500 26300
rect 119400 26300 119500 26400
rect 119400 26400 119500 26500
rect 119400 26500 119500 26600
rect 119400 26600 119500 26700
rect 119400 26700 119500 26800
rect 119400 26800 119500 26900
rect 119400 26900 119500 27000
rect 119400 27000 119500 27100
rect 119400 27100 119500 27200
rect 119500 22500 119600 22600
rect 119500 22600 119600 22700
rect 119500 22700 119600 22800
rect 119500 22800 119600 22900
rect 119500 22900 119600 23000
rect 119500 23000 119600 23100
rect 119500 23100 119600 23200
rect 119500 23200 119600 23300
rect 119500 23300 119600 23400
rect 119500 23400 119600 23500
rect 119500 23500 119600 23600
rect 119500 23600 119600 23700
rect 119500 23700 119600 23800
rect 119500 23800 119600 23900
rect 119500 23900 119600 24000
rect 119500 24000 119600 24100
rect 119500 24100 119600 24200
rect 119500 24200 119600 24300
rect 119500 24300 119600 24400
rect 119500 24400 119600 24500
rect 119500 24500 119600 24600
rect 119500 24600 119600 24700
rect 119500 24700 119600 24800
rect 119500 24800 119600 24900
rect 119500 24900 119600 25000
rect 119500 25000 119600 25100
rect 119500 25100 119600 25200
rect 119500 25200 119600 25300
rect 119500 25300 119600 25400
rect 119500 25400 119600 25500
rect 119500 25500 119600 25600
rect 119500 25600 119600 25700
rect 119500 25700 119600 25800
rect 119500 25800 119600 25900
rect 119500 25900 119600 26000
rect 119500 26000 119600 26100
rect 119500 26100 119600 26200
rect 119500 26200 119600 26300
rect 119500 26300 119600 26400
rect 119500 26400 119600 26500
rect 119500 26500 119600 26600
rect 119500 26600 119600 26700
rect 119500 26700 119600 26800
rect 119500 26800 119600 26900
rect 119500 26900 119600 27000
rect 119500 27000 119600 27100
rect 119500 27100 119600 27200
rect 119500 27200 119600 27300
rect 119600 22700 119700 22800
rect 119600 22800 119700 22900
rect 119600 22900 119700 23000
rect 119600 23000 119700 23100
rect 119600 23100 119700 23200
rect 119600 23200 119700 23300
rect 119600 23300 119700 23400
rect 119600 23400 119700 23500
rect 119600 23500 119700 23600
rect 119600 23600 119700 23700
rect 119600 23700 119700 23800
rect 119600 23800 119700 23900
rect 119600 23900 119700 24000
rect 119600 24000 119700 24100
rect 119600 24100 119700 24200
rect 119600 24200 119700 24300
rect 119600 24300 119700 24400
rect 119600 24400 119700 24500
rect 119600 24500 119700 24600
rect 119600 24600 119700 24700
rect 119600 24700 119700 24800
rect 119600 24800 119700 24900
rect 119600 24900 119700 25000
rect 119600 25000 119700 25100
rect 119600 25100 119700 25200
rect 119600 25200 119700 25300
rect 119600 25300 119700 25400
rect 119600 25400 119700 25500
rect 119600 25500 119700 25600
rect 119600 25600 119700 25700
rect 119600 25700 119700 25800
rect 119600 25800 119700 25900
rect 119600 25900 119700 26000
rect 119600 26000 119700 26100
rect 119600 26100 119700 26200
rect 119600 26200 119700 26300
rect 119600 26300 119700 26400
rect 119600 26400 119700 26500
rect 119600 26500 119700 26600
rect 119600 26600 119700 26700
rect 119600 26700 119700 26800
rect 119600 26800 119700 26900
rect 119600 26900 119700 27000
rect 119600 27000 119700 27100
rect 119600 27100 119700 27200
rect 119600 27200 119700 27300
rect 119600 27300 119700 27400
rect 119700 23100 119800 23200
rect 119700 23200 119800 23300
rect 119700 23300 119800 23400
rect 119700 23400 119800 23500
rect 119700 23500 119800 23600
rect 119700 23600 119800 23700
rect 119700 23700 119800 23800
rect 119700 23800 119800 23900
rect 119700 23900 119800 24000
rect 119700 24000 119800 24100
rect 119700 24100 119800 24200
rect 119700 24700 119800 24800
rect 119700 24800 119800 24900
rect 119700 24900 119800 25000
rect 119700 25000 119800 25100
rect 119700 25100 119800 25200
rect 119700 25200 119800 25300
rect 119700 25300 119800 25400
rect 119700 25400 119800 25500
rect 119700 25500 119800 25600
rect 119700 25600 119800 25700
rect 119700 25700 119800 25800
rect 119700 25800 119800 25900
rect 119700 25900 119800 26000
rect 119700 26000 119800 26100
rect 119700 26100 119800 26200
rect 119700 26200 119800 26300
rect 119700 26300 119800 26400
rect 119700 26400 119800 26500
rect 119700 26500 119800 26600
rect 119700 26600 119800 26700
rect 119700 26700 119800 26800
rect 119700 26800 119800 26900
rect 119700 26900 119800 27000
rect 119700 27000 119800 27100
rect 119700 27100 119800 27200
rect 119700 27200 119800 27300
rect 119700 27300 119800 27400
rect 119700 27400 119800 27500
rect 119700 35600 119800 35700
rect 119700 35700 119800 35800
rect 119700 35800 119800 35900
rect 119700 35900 119800 36000
rect 119700 36000 119800 36100
rect 119700 36100 119800 36200
rect 119700 36200 119800 36300
rect 119700 36300 119800 36400
rect 119700 36400 119800 36500
rect 119800 24900 119900 25000
rect 119800 25000 119900 25100
rect 119800 25100 119900 25200
rect 119800 25200 119900 25300
rect 119800 25300 119900 25400
rect 119800 25400 119900 25500
rect 119800 25500 119900 25600
rect 119800 25600 119900 25700
rect 119800 25700 119900 25800
rect 119800 25800 119900 25900
rect 119800 25900 119900 26000
rect 119800 26000 119900 26100
rect 119800 26100 119900 26200
rect 119800 26200 119900 26300
rect 119800 26300 119900 26400
rect 119800 26400 119900 26500
rect 119800 26500 119900 26600
rect 119800 26600 119900 26700
rect 119800 26700 119900 26800
rect 119800 26800 119900 26900
rect 119800 26900 119900 27000
rect 119800 27000 119900 27100
rect 119800 27100 119900 27200
rect 119800 27200 119900 27300
rect 119800 27300 119900 27400
rect 119800 27400 119900 27500
rect 119800 35200 119900 35300
rect 119800 35300 119900 35400
rect 119800 35400 119900 35500
rect 119800 35500 119900 35600
rect 119800 35600 119900 35700
rect 119800 35700 119900 35800
rect 119800 35800 119900 35900
rect 119800 35900 119900 36000
rect 119800 36000 119900 36100
rect 119800 36100 119900 36200
rect 119800 36200 119900 36300
rect 119800 36300 119900 36400
rect 119800 36400 119900 36500
rect 119800 36500 119900 36600
rect 119800 36600 119900 36700
rect 119800 36700 119900 36800
rect 119800 36800 119900 36900
rect 119900 25100 120000 25200
rect 119900 25200 120000 25300
rect 119900 25300 120000 25400
rect 119900 25400 120000 25500
rect 119900 25500 120000 25600
rect 119900 25600 120000 25700
rect 119900 25700 120000 25800
rect 119900 25800 120000 25900
rect 119900 25900 120000 26000
rect 119900 26000 120000 26100
rect 119900 26100 120000 26200
rect 119900 26200 120000 26300
rect 119900 26300 120000 26400
rect 119900 26400 120000 26500
rect 119900 26500 120000 26600
rect 119900 26600 120000 26700
rect 119900 26700 120000 26800
rect 119900 26800 120000 26900
rect 119900 26900 120000 27000
rect 119900 27000 120000 27100
rect 119900 27100 120000 27200
rect 119900 27200 120000 27300
rect 119900 27300 120000 27400
rect 119900 27400 120000 27500
rect 119900 27500 120000 27600
rect 119900 35000 120000 35100
rect 119900 35100 120000 35200
rect 119900 35200 120000 35300
rect 119900 35300 120000 35400
rect 119900 35400 120000 35500
rect 119900 35500 120000 35600
rect 119900 35600 120000 35700
rect 119900 35700 120000 35800
rect 119900 35800 120000 35900
rect 119900 35900 120000 36000
rect 119900 36000 120000 36100
rect 119900 36100 120000 36200
rect 119900 36200 120000 36300
rect 119900 36300 120000 36400
rect 119900 36400 120000 36500
rect 119900 36500 120000 36600
rect 119900 36600 120000 36700
rect 119900 36700 120000 36800
rect 119900 36800 120000 36900
rect 119900 36900 120000 37000
rect 119900 37000 120000 37100
rect 120000 25200 120100 25300
rect 120000 25300 120100 25400
rect 120000 25400 120100 25500
rect 120000 25500 120100 25600
rect 120000 25600 120100 25700
rect 120000 25700 120100 25800
rect 120000 25800 120100 25900
rect 120000 25900 120100 26000
rect 120000 26000 120100 26100
rect 120000 26100 120100 26200
rect 120000 26200 120100 26300
rect 120000 26300 120100 26400
rect 120000 26400 120100 26500
rect 120000 26500 120100 26600
rect 120000 26600 120100 26700
rect 120000 26700 120100 26800
rect 120000 26800 120100 26900
rect 120000 26900 120100 27000
rect 120000 27000 120100 27100
rect 120000 27100 120100 27200
rect 120000 27200 120100 27300
rect 120000 27300 120100 27400
rect 120000 27400 120100 27500
rect 120000 27500 120100 27600
rect 120000 27600 120100 27700
rect 120000 34800 120100 34900
rect 120000 34900 120100 35000
rect 120000 35000 120100 35100
rect 120000 35100 120100 35200
rect 120000 35200 120100 35300
rect 120000 35300 120100 35400
rect 120000 35400 120100 35500
rect 120000 35500 120100 35600
rect 120000 35600 120100 35700
rect 120000 35700 120100 35800
rect 120000 35800 120100 35900
rect 120000 35900 120100 36000
rect 120000 36000 120100 36100
rect 120000 36100 120100 36200
rect 120000 36200 120100 36300
rect 120000 36300 120100 36400
rect 120000 36400 120100 36500
rect 120000 36500 120100 36600
rect 120000 36600 120100 36700
rect 120000 36700 120100 36800
rect 120000 36800 120100 36900
rect 120000 36900 120100 37000
rect 120000 37000 120100 37100
rect 120000 37100 120100 37200
rect 120000 37200 120100 37300
rect 120100 25300 120200 25400
rect 120100 25400 120200 25500
rect 120100 25500 120200 25600
rect 120100 25600 120200 25700
rect 120100 25700 120200 25800
rect 120100 25800 120200 25900
rect 120100 25900 120200 26000
rect 120100 26000 120200 26100
rect 120100 26100 120200 26200
rect 120100 26200 120200 26300
rect 120100 26300 120200 26400
rect 120100 26400 120200 26500
rect 120100 26500 120200 26600
rect 120100 26600 120200 26700
rect 120100 26700 120200 26800
rect 120100 26800 120200 26900
rect 120100 26900 120200 27000
rect 120100 27000 120200 27100
rect 120100 27100 120200 27200
rect 120100 27200 120200 27300
rect 120100 27300 120200 27400
rect 120100 27400 120200 27500
rect 120100 27500 120200 27600
rect 120100 27600 120200 27700
rect 120100 27700 120200 27800
rect 120100 34700 120200 34800
rect 120100 34800 120200 34900
rect 120100 34900 120200 35000
rect 120100 35000 120200 35100
rect 120100 35100 120200 35200
rect 120100 35200 120200 35300
rect 120100 35300 120200 35400
rect 120100 35400 120200 35500
rect 120100 35500 120200 35600
rect 120100 35600 120200 35700
rect 120100 35700 120200 35800
rect 120100 35800 120200 35900
rect 120100 35900 120200 36000
rect 120100 36000 120200 36100
rect 120100 36100 120200 36200
rect 120100 36200 120200 36300
rect 120100 36300 120200 36400
rect 120100 36400 120200 36500
rect 120100 36500 120200 36600
rect 120100 36600 120200 36700
rect 120100 36700 120200 36800
rect 120100 36800 120200 36900
rect 120100 36900 120200 37000
rect 120100 37000 120200 37100
rect 120100 37100 120200 37200
rect 120100 37200 120200 37300
rect 120100 37300 120200 37400
rect 120200 25500 120300 25600
rect 120200 25600 120300 25700
rect 120200 25700 120300 25800
rect 120200 25800 120300 25900
rect 120200 25900 120300 26000
rect 120200 26000 120300 26100
rect 120200 26100 120300 26200
rect 120200 26200 120300 26300
rect 120200 26300 120300 26400
rect 120200 26400 120300 26500
rect 120200 26500 120300 26600
rect 120200 26600 120300 26700
rect 120200 26700 120300 26800
rect 120200 26800 120300 26900
rect 120200 26900 120300 27000
rect 120200 27000 120300 27100
rect 120200 27100 120300 27200
rect 120200 27200 120300 27300
rect 120200 27300 120300 27400
rect 120200 27400 120300 27500
rect 120200 27500 120300 27600
rect 120200 27600 120300 27700
rect 120200 27700 120300 27800
rect 120200 27800 120300 27900
rect 120200 34500 120300 34600
rect 120200 34600 120300 34700
rect 120200 34700 120300 34800
rect 120200 34800 120300 34900
rect 120200 34900 120300 35000
rect 120200 35000 120300 35100
rect 120200 35100 120300 35200
rect 120200 35200 120300 35300
rect 120200 35300 120300 35400
rect 120200 35400 120300 35500
rect 120200 35500 120300 35600
rect 120200 35600 120300 35700
rect 120200 35700 120300 35800
rect 120200 35800 120300 35900
rect 120200 35900 120300 36000
rect 120200 36000 120300 36100
rect 120200 36100 120300 36200
rect 120200 36200 120300 36300
rect 120200 36300 120300 36400
rect 120200 36400 120300 36500
rect 120200 36500 120300 36600
rect 120200 36600 120300 36700
rect 120200 36700 120300 36800
rect 120200 36800 120300 36900
rect 120200 36900 120300 37000
rect 120200 37000 120300 37100
rect 120200 37100 120300 37200
rect 120200 37200 120300 37300
rect 120200 37300 120300 37400
rect 120200 37400 120300 37500
rect 120300 25600 120400 25700
rect 120300 25700 120400 25800
rect 120300 25800 120400 25900
rect 120300 25900 120400 26000
rect 120300 26000 120400 26100
rect 120300 26100 120400 26200
rect 120300 26200 120400 26300
rect 120300 26300 120400 26400
rect 120300 26400 120400 26500
rect 120300 26500 120400 26600
rect 120300 26600 120400 26700
rect 120300 26700 120400 26800
rect 120300 26800 120400 26900
rect 120300 26900 120400 27000
rect 120300 27000 120400 27100
rect 120300 27100 120400 27200
rect 120300 27200 120400 27300
rect 120300 27300 120400 27400
rect 120300 27400 120400 27500
rect 120300 27500 120400 27600
rect 120300 27600 120400 27700
rect 120300 27700 120400 27800
rect 120300 27800 120400 27900
rect 120300 27900 120400 28000
rect 120300 34400 120400 34500
rect 120300 34500 120400 34600
rect 120300 34600 120400 34700
rect 120300 34700 120400 34800
rect 120300 34800 120400 34900
rect 120300 34900 120400 35000
rect 120300 35000 120400 35100
rect 120300 35100 120400 35200
rect 120300 35200 120400 35300
rect 120300 35300 120400 35400
rect 120300 35400 120400 35500
rect 120300 35500 120400 35600
rect 120300 35600 120400 35700
rect 120300 35700 120400 35800
rect 120300 35800 120400 35900
rect 120300 35900 120400 36000
rect 120300 36000 120400 36100
rect 120300 36100 120400 36200
rect 120300 36200 120400 36300
rect 120300 36300 120400 36400
rect 120300 36400 120400 36500
rect 120300 36500 120400 36600
rect 120300 36600 120400 36700
rect 120300 36700 120400 36800
rect 120300 36800 120400 36900
rect 120300 36900 120400 37000
rect 120300 37000 120400 37100
rect 120300 37100 120400 37200
rect 120300 37200 120400 37300
rect 120300 37300 120400 37400
rect 120300 37400 120400 37500
rect 120300 37500 120400 37600
rect 120400 25700 120500 25800
rect 120400 25800 120500 25900
rect 120400 25900 120500 26000
rect 120400 26000 120500 26100
rect 120400 26100 120500 26200
rect 120400 26200 120500 26300
rect 120400 26300 120500 26400
rect 120400 26400 120500 26500
rect 120400 26500 120500 26600
rect 120400 26600 120500 26700
rect 120400 26700 120500 26800
rect 120400 26800 120500 26900
rect 120400 26900 120500 27000
rect 120400 27000 120500 27100
rect 120400 27100 120500 27200
rect 120400 27200 120500 27300
rect 120400 27300 120500 27400
rect 120400 27400 120500 27500
rect 120400 27500 120500 27600
rect 120400 27600 120500 27700
rect 120400 27700 120500 27800
rect 120400 27800 120500 27900
rect 120400 27900 120500 28000
rect 120400 28000 120500 28100
rect 120400 34300 120500 34400
rect 120400 34400 120500 34500
rect 120400 34500 120500 34600
rect 120400 34600 120500 34700
rect 120400 34700 120500 34800
rect 120400 34800 120500 34900
rect 120400 34900 120500 35000
rect 120400 35000 120500 35100
rect 120400 35100 120500 35200
rect 120400 35200 120500 35300
rect 120400 35300 120500 35400
rect 120400 35400 120500 35500
rect 120400 35500 120500 35600
rect 120400 35600 120500 35700
rect 120400 35700 120500 35800
rect 120400 35800 120500 35900
rect 120400 35900 120500 36000
rect 120400 36000 120500 36100
rect 120400 36100 120500 36200
rect 120400 36200 120500 36300
rect 120400 36300 120500 36400
rect 120400 36400 120500 36500
rect 120400 36500 120500 36600
rect 120400 36600 120500 36700
rect 120400 36700 120500 36800
rect 120400 36800 120500 36900
rect 120400 36900 120500 37000
rect 120400 37000 120500 37100
rect 120400 37100 120500 37200
rect 120400 37200 120500 37300
rect 120400 37300 120500 37400
rect 120400 37400 120500 37500
rect 120400 37500 120500 37600
rect 120400 37600 120500 37700
rect 120500 25900 120600 26000
rect 120500 26000 120600 26100
rect 120500 26100 120600 26200
rect 120500 26200 120600 26300
rect 120500 26300 120600 26400
rect 120500 26400 120600 26500
rect 120500 26500 120600 26600
rect 120500 26600 120600 26700
rect 120500 26700 120600 26800
rect 120500 26800 120600 26900
rect 120500 26900 120600 27000
rect 120500 27000 120600 27100
rect 120500 27100 120600 27200
rect 120500 27200 120600 27300
rect 120500 27300 120600 27400
rect 120500 27400 120600 27500
rect 120500 27500 120600 27600
rect 120500 27600 120600 27700
rect 120500 27700 120600 27800
rect 120500 27800 120600 27900
rect 120500 27900 120600 28000
rect 120500 28000 120600 28100
rect 120500 28100 120600 28200
rect 120500 34200 120600 34300
rect 120500 34300 120600 34400
rect 120500 34400 120600 34500
rect 120500 34500 120600 34600
rect 120500 34600 120600 34700
rect 120500 34700 120600 34800
rect 120500 34800 120600 34900
rect 120500 34900 120600 35000
rect 120500 35000 120600 35100
rect 120500 35100 120600 35200
rect 120500 35200 120600 35300
rect 120500 35300 120600 35400
rect 120500 35400 120600 35500
rect 120500 35500 120600 35600
rect 120500 35600 120600 35700
rect 120500 35700 120600 35800
rect 120500 35800 120600 35900
rect 120500 35900 120600 36000
rect 120500 36000 120600 36100
rect 120500 36100 120600 36200
rect 120500 36200 120600 36300
rect 120500 36300 120600 36400
rect 120500 36400 120600 36500
rect 120500 36500 120600 36600
rect 120500 36600 120600 36700
rect 120500 36700 120600 36800
rect 120500 36800 120600 36900
rect 120500 36900 120600 37000
rect 120500 37000 120600 37100
rect 120500 37100 120600 37200
rect 120500 37200 120600 37300
rect 120500 37300 120600 37400
rect 120500 37400 120600 37500
rect 120500 37500 120600 37600
rect 120500 37600 120600 37700
rect 120500 37700 120600 37800
rect 120600 26000 120700 26100
rect 120600 26100 120700 26200
rect 120600 26200 120700 26300
rect 120600 26300 120700 26400
rect 120600 26400 120700 26500
rect 120600 26500 120700 26600
rect 120600 26600 120700 26700
rect 120600 26700 120700 26800
rect 120600 26800 120700 26900
rect 120600 26900 120700 27000
rect 120600 27000 120700 27100
rect 120600 27100 120700 27200
rect 120600 27200 120700 27300
rect 120600 27300 120700 27400
rect 120600 27400 120700 27500
rect 120600 27500 120700 27600
rect 120600 27600 120700 27700
rect 120600 27700 120700 27800
rect 120600 27800 120700 27900
rect 120600 27900 120700 28000
rect 120600 28000 120700 28100
rect 120600 28100 120700 28200
rect 120600 28200 120700 28300
rect 120600 34100 120700 34200
rect 120600 34200 120700 34300
rect 120600 34300 120700 34400
rect 120600 34400 120700 34500
rect 120600 34500 120700 34600
rect 120600 34600 120700 34700
rect 120600 34700 120700 34800
rect 120600 34800 120700 34900
rect 120600 34900 120700 35000
rect 120600 35000 120700 35100
rect 120600 35100 120700 35200
rect 120600 35200 120700 35300
rect 120600 35300 120700 35400
rect 120600 35400 120700 35500
rect 120600 35500 120700 35600
rect 120600 35600 120700 35700
rect 120600 35700 120700 35800
rect 120600 35800 120700 35900
rect 120600 35900 120700 36000
rect 120600 36000 120700 36100
rect 120600 36100 120700 36200
rect 120600 36200 120700 36300
rect 120600 36300 120700 36400
rect 120600 36400 120700 36500
rect 120600 36500 120700 36600
rect 120600 36600 120700 36700
rect 120600 36700 120700 36800
rect 120600 36800 120700 36900
rect 120600 36900 120700 37000
rect 120600 37000 120700 37100
rect 120600 37100 120700 37200
rect 120600 37200 120700 37300
rect 120600 37300 120700 37400
rect 120600 37400 120700 37500
rect 120600 37500 120700 37600
rect 120600 37600 120700 37700
rect 120600 37700 120700 37800
rect 120600 37800 120700 37900
rect 120700 26100 120800 26200
rect 120700 26200 120800 26300
rect 120700 26300 120800 26400
rect 120700 26400 120800 26500
rect 120700 26500 120800 26600
rect 120700 26600 120800 26700
rect 120700 26700 120800 26800
rect 120700 26800 120800 26900
rect 120700 26900 120800 27000
rect 120700 27000 120800 27100
rect 120700 27100 120800 27200
rect 120700 27200 120800 27300
rect 120700 27300 120800 27400
rect 120700 27400 120800 27500
rect 120700 27500 120800 27600
rect 120700 27600 120800 27700
rect 120700 27700 120800 27800
rect 120700 27800 120800 27900
rect 120700 27900 120800 28000
rect 120700 28000 120800 28100
rect 120700 28100 120800 28200
rect 120700 28200 120800 28300
rect 120700 28300 120800 28400
rect 120700 34000 120800 34100
rect 120700 34100 120800 34200
rect 120700 34200 120800 34300
rect 120700 34300 120800 34400
rect 120700 34400 120800 34500
rect 120700 34500 120800 34600
rect 120700 34600 120800 34700
rect 120700 34700 120800 34800
rect 120700 34800 120800 34900
rect 120700 34900 120800 35000
rect 120700 35000 120800 35100
rect 120700 35100 120800 35200
rect 120700 35200 120800 35300
rect 120700 35300 120800 35400
rect 120700 35400 120800 35500
rect 120700 35500 120800 35600
rect 120700 35600 120800 35700
rect 120700 35700 120800 35800
rect 120700 35800 120800 35900
rect 120700 35900 120800 36000
rect 120700 36000 120800 36100
rect 120700 36100 120800 36200
rect 120700 36200 120800 36300
rect 120700 36300 120800 36400
rect 120700 36400 120800 36500
rect 120700 36500 120800 36600
rect 120700 36600 120800 36700
rect 120700 36700 120800 36800
rect 120700 36800 120800 36900
rect 120700 36900 120800 37000
rect 120700 37000 120800 37100
rect 120700 37100 120800 37200
rect 120700 37200 120800 37300
rect 120700 37300 120800 37400
rect 120700 37400 120800 37500
rect 120700 37500 120800 37600
rect 120700 37600 120800 37700
rect 120700 37700 120800 37800
rect 120700 37800 120800 37900
rect 120700 37900 120800 38000
rect 120800 26200 120900 26300
rect 120800 26300 120900 26400
rect 120800 26400 120900 26500
rect 120800 26500 120900 26600
rect 120800 26600 120900 26700
rect 120800 26700 120900 26800
rect 120800 26800 120900 26900
rect 120800 26900 120900 27000
rect 120800 27000 120900 27100
rect 120800 27100 120900 27200
rect 120800 27200 120900 27300
rect 120800 27300 120900 27400
rect 120800 27400 120900 27500
rect 120800 27500 120900 27600
rect 120800 27600 120900 27700
rect 120800 27700 120900 27800
rect 120800 27800 120900 27900
rect 120800 27900 120900 28000
rect 120800 28000 120900 28100
rect 120800 28100 120900 28200
rect 120800 28200 120900 28300
rect 120800 28300 120900 28400
rect 120800 28400 120900 28500
rect 120800 34000 120900 34100
rect 120800 34100 120900 34200
rect 120800 34200 120900 34300
rect 120800 34300 120900 34400
rect 120800 34400 120900 34500
rect 120800 34500 120900 34600
rect 120800 34600 120900 34700
rect 120800 34700 120900 34800
rect 120800 34800 120900 34900
rect 120800 34900 120900 35000
rect 120800 35000 120900 35100
rect 120800 35100 120900 35200
rect 120800 35200 120900 35300
rect 120800 35300 120900 35400
rect 120800 35400 120900 35500
rect 120800 35500 120900 35600
rect 120800 35600 120900 35700
rect 120800 35700 120900 35800
rect 120800 35800 120900 35900
rect 120800 35900 120900 36000
rect 120800 36000 120900 36100
rect 120800 36100 120900 36200
rect 120800 36200 120900 36300
rect 120800 36300 120900 36400
rect 120800 36400 120900 36500
rect 120800 36500 120900 36600
rect 120800 36600 120900 36700
rect 120800 36700 120900 36800
rect 120800 36800 120900 36900
rect 120800 36900 120900 37000
rect 120800 37000 120900 37100
rect 120800 37100 120900 37200
rect 120800 37200 120900 37300
rect 120800 37300 120900 37400
rect 120800 37400 120900 37500
rect 120800 37500 120900 37600
rect 120800 37600 120900 37700
rect 120800 37700 120900 37800
rect 120800 37800 120900 37900
rect 120800 37900 120900 38000
rect 120900 26300 121000 26400
rect 120900 26400 121000 26500
rect 120900 26500 121000 26600
rect 120900 26600 121000 26700
rect 120900 26700 121000 26800
rect 120900 26800 121000 26900
rect 120900 26900 121000 27000
rect 120900 27000 121000 27100
rect 120900 27100 121000 27200
rect 120900 27200 121000 27300
rect 120900 27300 121000 27400
rect 120900 27400 121000 27500
rect 120900 27500 121000 27600
rect 120900 27600 121000 27700
rect 120900 27700 121000 27800
rect 120900 27800 121000 27900
rect 120900 27900 121000 28000
rect 120900 28000 121000 28100
rect 120900 28100 121000 28200
rect 120900 28200 121000 28300
rect 120900 28300 121000 28400
rect 120900 28400 121000 28500
rect 120900 33900 121000 34000
rect 120900 34000 121000 34100
rect 120900 34100 121000 34200
rect 120900 34200 121000 34300
rect 120900 34300 121000 34400
rect 120900 34400 121000 34500
rect 120900 34500 121000 34600
rect 120900 34600 121000 34700
rect 120900 34700 121000 34800
rect 120900 34800 121000 34900
rect 120900 34900 121000 35000
rect 120900 35000 121000 35100
rect 120900 35100 121000 35200
rect 120900 35200 121000 35300
rect 120900 35300 121000 35400
rect 120900 35400 121000 35500
rect 120900 35500 121000 35600
rect 120900 35600 121000 35700
rect 120900 35700 121000 35800
rect 120900 35800 121000 35900
rect 120900 35900 121000 36000
rect 120900 36000 121000 36100
rect 120900 36100 121000 36200
rect 120900 36200 121000 36300
rect 120900 36300 121000 36400
rect 120900 36400 121000 36500
rect 120900 36500 121000 36600
rect 120900 36600 121000 36700
rect 120900 36700 121000 36800
rect 120900 36800 121000 36900
rect 120900 36900 121000 37000
rect 120900 37000 121000 37100
rect 120900 37100 121000 37200
rect 120900 37200 121000 37300
rect 120900 37300 121000 37400
rect 120900 37400 121000 37500
rect 120900 37500 121000 37600
rect 120900 37600 121000 37700
rect 120900 37700 121000 37800
rect 120900 37800 121000 37900
rect 120900 37900 121000 38000
rect 120900 38000 121000 38100
rect 121000 26400 121100 26500
rect 121000 26500 121100 26600
rect 121000 26600 121100 26700
rect 121000 26700 121100 26800
rect 121000 26800 121100 26900
rect 121000 26900 121100 27000
rect 121000 27000 121100 27100
rect 121000 27100 121100 27200
rect 121000 27200 121100 27300
rect 121000 27300 121100 27400
rect 121000 27400 121100 27500
rect 121000 27500 121100 27600
rect 121000 27600 121100 27700
rect 121000 27700 121100 27800
rect 121000 27800 121100 27900
rect 121000 27900 121100 28000
rect 121000 28000 121100 28100
rect 121000 28100 121100 28200
rect 121000 28200 121100 28300
rect 121000 28300 121100 28400
rect 121000 28400 121100 28500
rect 121000 28500 121100 28600
rect 121000 33800 121100 33900
rect 121000 33900 121100 34000
rect 121000 34000 121100 34100
rect 121000 34100 121100 34200
rect 121000 34200 121100 34300
rect 121000 34300 121100 34400
rect 121000 34400 121100 34500
rect 121000 34500 121100 34600
rect 121000 34600 121100 34700
rect 121000 34700 121100 34800
rect 121000 34800 121100 34900
rect 121000 34900 121100 35000
rect 121000 35000 121100 35100
rect 121000 35100 121100 35200
rect 121000 35200 121100 35300
rect 121000 35300 121100 35400
rect 121000 35400 121100 35500
rect 121000 35500 121100 35600
rect 121000 35600 121100 35700
rect 121000 35700 121100 35800
rect 121000 35800 121100 35900
rect 121000 35900 121100 36000
rect 121000 36000 121100 36100
rect 121000 36100 121100 36200
rect 121000 36200 121100 36300
rect 121000 36300 121100 36400
rect 121000 36400 121100 36500
rect 121000 36500 121100 36600
rect 121000 36600 121100 36700
rect 121000 36700 121100 36800
rect 121000 36800 121100 36900
rect 121000 36900 121100 37000
rect 121000 37000 121100 37100
rect 121000 37100 121100 37200
rect 121000 37200 121100 37300
rect 121000 37300 121100 37400
rect 121000 37400 121100 37500
rect 121000 37500 121100 37600
rect 121000 37600 121100 37700
rect 121000 37700 121100 37800
rect 121000 37800 121100 37900
rect 121000 37900 121100 38000
rect 121000 38000 121100 38100
rect 121100 26500 121200 26600
rect 121100 26600 121200 26700
rect 121100 26700 121200 26800
rect 121100 26800 121200 26900
rect 121100 26900 121200 27000
rect 121100 27000 121200 27100
rect 121100 27100 121200 27200
rect 121100 27200 121200 27300
rect 121100 27300 121200 27400
rect 121100 27400 121200 27500
rect 121100 27500 121200 27600
rect 121100 27600 121200 27700
rect 121100 27700 121200 27800
rect 121100 27800 121200 27900
rect 121100 27900 121200 28000
rect 121100 28000 121200 28100
rect 121100 28100 121200 28200
rect 121100 28200 121200 28300
rect 121100 28300 121200 28400
rect 121100 28400 121200 28500
rect 121100 28500 121200 28600
rect 121100 28600 121200 28700
rect 121100 33800 121200 33900
rect 121100 33900 121200 34000
rect 121100 34000 121200 34100
rect 121100 34100 121200 34200
rect 121100 34200 121200 34300
rect 121100 34300 121200 34400
rect 121100 34400 121200 34500
rect 121100 34500 121200 34600
rect 121100 34600 121200 34700
rect 121100 34700 121200 34800
rect 121100 34800 121200 34900
rect 121100 34900 121200 35000
rect 121100 35000 121200 35100
rect 121100 35100 121200 35200
rect 121100 35200 121200 35300
rect 121100 35300 121200 35400
rect 121100 35400 121200 35500
rect 121100 35500 121200 35600
rect 121100 35600 121200 35700
rect 121100 35700 121200 35800
rect 121100 35800 121200 35900
rect 121100 35900 121200 36000
rect 121100 36000 121200 36100
rect 121100 36100 121200 36200
rect 121100 36200 121200 36300
rect 121100 36300 121200 36400
rect 121100 36400 121200 36500
rect 121100 36500 121200 36600
rect 121100 36600 121200 36700
rect 121100 36700 121200 36800
rect 121100 36800 121200 36900
rect 121100 36900 121200 37000
rect 121100 37000 121200 37100
rect 121100 37100 121200 37200
rect 121100 37200 121200 37300
rect 121100 37300 121200 37400
rect 121100 37400 121200 37500
rect 121100 37500 121200 37600
rect 121100 37600 121200 37700
rect 121100 37700 121200 37800
rect 121100 37800 121200 37900
rect 121100 37900 121200 38000
rect 121100 38000 121200 38100
rect 121100 38100 121200 38200
rect 121200 26600 121300 26700
rect 121200 26700 121300 26800
rect 121200 26800 121300 26900
rect 121200 26900 121300 27000
rect 121200 27000 121300 27100
rect 121200 27100 121300 27200
rect 121200 27200 121300 27300
rect 121200 27300 121300 27400
rect 121200 27400 121300 27500
rect 121200 27500 121300 27600
rect 121200 27600 121300 27700
rect 121200 27700 121300 27800
rect 121200 27800 121300 27900
rect 121200 27900 121300 28000
rect 121200 28000 121300 28100
rect 121200 28100 121300 28200
rect 121200 28200 121300 28300
rect 121200 28300 121300 28400
rect 121200 28400 121300 28500
rect 121200 28500 121300 28600
rect 121200 28600 121300 28700
rect 121200 28700 121300 28800
rect 121200 33700 121300 33800
rect 121200 33800 121300 33900
rect 121200 33900 121300 34000
rect 121200 34000 121300 34100
rect 121200 34100 121300 34200
rect 121200 34200 121300 34300
rect 121200 34300 121300 34400
rect 121200 34400 121300 34500
rect 121200 34500 121300 34600
rect 121200 34600 121300 34700
rect 121200 34700 121300 34800
rect 121200 34800 121300 34900
rect 121200 34900 121300 35000
rect 121200 35000 121300 35100
rect 121200 35100 121300 35200
rect 121200 35200 121300 35300
rect 121200 35300 121300 35400
rect 121200 35400 121300 35500
rect 121200 35500 121300 35600
rect 121200 35600 121300 35700
rect 121200 35700 121300 35800
rect 121200 35800 121300 35900
rect 121200 35900 121300 36000
rect 121200 36000 121300 36100
rect 121200 36100 121300 36200
rect 121200 36200 121300 36300
rect 121200 36300 121300 36400
rect 121200 36400 121300 36500
rect 121200 36500 121300 36600
rect 121200 36600 121300 36700
rect 121200 36700 121300 36800
rect 121200 36800 121300 36900
rect 121200 36900 121300 37000
rect 121200 37000 121300 37100
rect 121200 37100 121300 37200
rect 121200 37200 121300 37300
rect 121200 37300 121300 37400
rect 121200 37400 121300 37500
rect 121200 37500 121300 37600
rect 121200 37600 121300 37700
rect 121200 37700 121300 37800
rect 121200 37800 121300 37900
rect 121200 37900 121300 38000
rect 121200 38000 121300 38100
rect 121200 38100 121300 38200
rect 121300 26700 121400 26800
rect 121300 26800 121400 26900
rect 121300 26900 121400 27000
rect 121300 27000 121400 27100
rect 121300 27100 121400 27200
rect 121300 27200 121400 27300
rect 121300 27300 121400 27400
rect 121300 27400 121400 27500
rect 121300 27500 121400 27600
rect 121300 27600 121400 27700
rect 121300 27700 121400 27800
rect 121300 27800 121400 27900
rect 121300 27900 121400 28000
rect 121300 28000 121400 28100
rect 121300 28100 121400 28200
rect 121300 28200 121400 28300
rect 121300 28300 121400 28400
rect 121300 28400 121400 28500
rect 121300 28500 121400 28600
rect 121300 28600 121400 28700
rect 121300 28700 121400 28800
rect 121300 28800 121400 28900
rect 121300 33700 121400 33800
rect 121300 33800 121400 33900
rect 121300 33900 121400 34000
rect 121300 34000 121400 34100
rect 121300 34100 121400 34200
rect 121300 34200 121400 34300
rect 121300 34300 121400 34400
rect 121300 34400 121400 34500
rect 121300 34500 121400 34600
rect 121300 34600 121400 34700
rect 121300 34700 121400 34800
rect 121300 34800 121400 34900
rect 121300 34900 121400 35000
rect 121300 35000 121400 35100
rect 121300 35100 121400 35200
rect 121300 35200 121400 35300
rect 121300 35300 121400 35400
rect 121300 35400 121400 35500
rect 121300 35500 121400 35600
rect 121300 35600 121400 35700
rect 121300 35700 121400 35800
rect 121300 35800 121400 35900
rect 121300 35900 121400 36000
rect 121300 36000 121400 36100
rect 121300 36100 121400 36200
rect 121300 36200 121400 36300
rect 121300 36300 121400 36400
rect 121300 36400 121400 36500
rect 121300 36500 121400 36600
rect 121300 36600 121400 36700
rect 121300 36700 121400 36800
rect 121300 36800 121400 36900
rect 121300 36900 121400 37000
rect 121300 37000 121400 37100
rect 121300 37100 121400 37200
rect 121300 37200 121400 37300
rect 121300 37300 121400 37400
rect 121300 37400 121400 37500
rect 121300 37500 121400 37600
rect 121300 37600 121400 37700
rect 121300 37700 121400 37800
rect 121300 37800 121400 37900
rect 121300 37900 121400 38000
rect 121300 38000 121400 38100
rect 121300 38100 121400 38200
rect 121300 38200 121400 38300
rect 121400 26800 121500 26900
rect 121400 26900 121500 27000
rect 121400 27000 121500 27100
rect 121400 27100 121500 27200
rect 121400 27200 121500 27300
rect 121400 27300 121500 27400
rect 121400 27400 121500 27500
rect 121400 27500 121500 27600
rect 121400 27600 121500 27700
rect 121400 27700 121500 27800
rect 121400 27800 121500 27900
rect 121400 27900 121500 28000
rect 121400 28000 121500 28100
rect 121400 28100 121500 28200
rect 121400 28200 121500 28300
rect 121400 28300 121500 28400
rect 121400 28400 121500 28500
rect 121400 28500 121500 28600
rect 121400 28600 121500 28700
rect 121400 28700 121500 28800
rect 121400 28800 121500 28900
rect 121400 28900 121500 29000
rect 121400 33600 121500 33700
rect 121400 33700 121500 33800
rect 121400 33800 121500 33900
rect 121400 33900 121500 34000
rect 121400 34000 121500 34100
rect 121400 34100 121500 34200
rect 121400 34200 121500 34300
rect 121400 34300 121500 34400
rect 121400 34400 121500 34500
rect 121400 34500 121500 34600
rect 121400 34600 121500 34700
rect 121400 34700 121500 34800
rect 121400 34800 121500 34900
rect 121400 34900 121500 35000
rect 121400 35000 121500 35100
rect 121400 35100 121500 35200
rect 121400 35200 121500 35300
rect 121400 35300 121500 35400
rect 121400 35400 121500 35500
rect 121400 35500 121500 35600
rect 121400 35600 121500 35700
rect 121400 35700 121500 35800
rect 121400 36300 121500 36400
rect 121400 36400 121500 36500
rect 121400 36500 121500 36600
rect 121400 36600 121500 36700
rect 121400 36700 121500 36800
rect 121400 36800 121500 36900
rect 121400 36900 121500 37000
rect 121400 37000 121500 37100
rect 121400 37100 121500 37200
rect 121400 37200 121500 37300
rect 121400 37300 121500 37400
rect 121400 37400 121500 37500
rect 121400 37500 121500 37600
rect 121400 37600 121500 37700
rect 121400 37700 121500 37800
rect 121400 37800 121500 37900
rect 121400 37900 121500 38000
rect 121400 38000 121500 38100
rect 121400 38100 121500 38200
rect 121400 38200 121500 38300
rect 121500 26900 121600 27000
rect 121500 27000 121600 27100
rect 121500 27100 121600 27200
rect 121500 27200 121600 27300
rect 121500 27300 121600 27400
rect 121500 27400 121600 27500
rect 121500 27500 121600 27600
rect 121500 27600 121600 27700
rect 121500 27700 121600 27800
rect 121500 27800 121600 27900
rect 121500 27900 121600 28000
rect 121500 28000 121600 28100
rect 121500 28100 121600 28200
rect 121500 28200 121600 28300
rect 121500 28300 121600 28400
rect 121500 28400 121600 28500
rect 121500 28500 121600 28600
rect 121500 28600 121600 28700
rect 121500 28700 121600 28800
rect 121500 28800 121600 28900
rect 121500 28900 121600 29000
rect 121500 29000 121600 29100
rect 121500 33600 121600 33700
rect 121500 33700 121600 33800
rect 121500 33800 121600 33900
rect 121500 33900 121600 34000
rect 121500 34000 121600 34100
rect 121500 34100 121600 34200
rect 121500 34200 121600 34300
rect 121500 34300 121600 34400
rect 121500 34400 121600 34500
rect 121500 34500 121600 34600
rect 121500 34600 121600 34700
rect 121500 34700 121600 34800
rect 121500 34800 121600 34900
rect 121500 34900 121600 35000
rect 121500 35000 121600 35100
rect 121500 35100 121600 35200
rect 121500 35200 121600 35300
rect 121500 35300 121600 35400
rect 121500 35400 121600 35500
rect 121500 35500 121600 35600
rect 121500 35600 121600 35700
rect 121500 36500 121600 36600
rect 121500 36600 121600 36700
rect 121500 36700 121600 36800
rect 121500 36800 121600 36900
rect 121500 36900 121600 37000
rect 121500 37000 121600 37100
rect 121500 37100 121600 37200
rect 121500 37200 121600 37300
rect 121500 37300 121600 37400
rect 121500 37400 121600 37500
rect 121500 37500 121600 37600
rect 121500 37600 121600 37700
rect 121500 37700 121600 37800
rect 121500 37800 121600 37900
rect 121500 37900 121600 38000
rect 121500 38000 121600 38100
rect 121500 38100 121600 38200
rect 121500 38200 121600 38300
rect 121600 27000 121700 27100
rect 121600 27100 121700 27200
rect 121600 27200 121700 27300
rect 121600 27300 121700 27400
rect 121600 27400 121700 27500
rect 121600 27500 121700 27600
rect 121600 27600 121700 27700
rect 121600 27700 121700 27800
rect 121600 27800 121700 27900
rect 121600 27900 121700 28000
rect 121600 28000 121700 28100
rect 121600 28100 121700 28200
rect 121600 28200 121700 28300
rect 121600 28300 121700 28400
rect 121600 28400 121700 28500
rect 121600 28500 121700 28600
rect 121600 28600 121700 28700
rect 121600 28700 121700 28800
rect 121600 28800 121700 28900
rect 121600 28900 121700 29000
rect 121600 29000 121700 29100
rect 121600 33500 121700 33600
rect 121600 33600 121700 33700
rect 121600 33700 121700 33800
rect 121600 33800 121700 33900
rect 121600 33900 121700 34000
rect 121600 34000 121700 34100
rect 121600 34100 121700 34200
rect 121600 34200 121700 34300
rect 121600 34300 121700 34400
rect 121600 34400 121700 34500
rect 121600 34500 121700 34600
rect 121600 34600 121700 34700
rect 121600 34700 121700 34800
rect 121600 34800 121700 34900
rect 121600 34900 121700 35000
rect 121600 35000 121700 35100
rect 121600 35100 121700 35200
rect 121600 35200 121700 35300
rect 121600 35300 121700 35400
rect 121600 35400 121700 35500
rect 121600 35500 121700 35600
rect 121600 36600 121700 36700
rect 121600 36700 121700 36800
rect 121600 36800 121700 36900
rect 121600 36900 121700 37000
rect 121600 37000 121700 37100
rect 121600 37100 121700 37200
rect 121600 37200 121700 37300
rect 121600 37300 121700 37400
rect 121600 37400 121700 37500
rect 121600 37500 121700 37600
rect 121600 37600 121700 37700
rect 121600 37700 121700 37800
rect 121600 37800 121700 37900
rect 121600 37900 121700 38000
rect 121600 38000 121700 38100
rect 121600 38100 121700 38200
rect 121600 38200 121700 38300
rect 121700 27000 121800 27100
rect 121700 27100 121800 27200
rect 121700 27200 121800 27300
rect 121700 27300 121800 27400
rect 121700 27400 121800 27500
rect 121700 27500 121800 27600
rect 121700 27600 121800 27700
rect 121700 27700 121800 27800
rect 121700 27800 121800 27900
rect 121700 27900 121800 28000
rect 121700 28000 121800 28100
rect 121700 28100 121800 28200
rect 121700 28200 121800 28300
rect 121700 28300 121800 28400
rect 121700 28400 121800 28500
rect 121700 28500 121800 28600
rect 121700 28600 121800 28700
rect 121700 28700 121800 28800
rect 121700 28800 121800 28900
rect 121700 28900 121800 29000
rect 121700 29000 121800 29100
rect 121700 29100 121800 29200
rect 121700 33400 121800 33500
rect 121700 33500 121800 33600
rect 121700 33600 121800 33700
rect 121700 33700 121800 33800
rect 121700 33800 121800 33900
rect 121700 33900 121800 34000
rect 121700 34000 121800 34100
rect 121700 34100 121800 34200
rect 121700 34200 121800 34300
rect 121700 34300 121800 34400
rect 121700 34400 121800 34500
rect 121700 34500 121800 34600
rect 121700 34600 121800 34700
rect 121700 34700 121800 34800
rect 121700 34800 121800 34900
rect 121700 34900 121800 35000
rect 121700 35000 121800 35100
rect 121700 35100 121800 35200
rect 121700 35200 121800 35300
rect 121700 35300 121800 35400
rect 121700 35400 121800 35500
rect 121700 36700 121800 36800
rect 121700 36800 121800 36900
rect 121700 36900 121800 37000
rect 121700 37000 121800 37100
rect 121700 37100 121800 37200
rect 121700 37200 121800 37300
rect 121700 37300 121800 37400
rect 121700 37400 121800 37500
rect 121700 37500 121800 37600
rect 121700 37600 121800 37700
rect 121700 37700 121800 37800
rect 121700 37800 121800 37900
rect 121700 37900 121800 38000
rect 121700 38000 121800 38100
rect 121700 38100 121800 38200
rect 121700 38200 121800 38300
rect 121700 38300 121800 38400
rect 121800 27100 121900 27200
rect 121800 27200 121900 27300
rect 121800 27300 121900 27400
rect 121800 27400 121900 27500
rect 121800 27500 121900 27600
rect 121800 27600 121900 27700
rect 121800 27700 121900 27800
rect 121800 27800 121900 27900
rect 121800 27900 121900 28000
rect 121800 28000 121900 28100
rect 121800 28100 121900 28200
rect 121800 28200 121900 28300
rect 121800 28300 121900 28400
rect 121800 28400 121900 28500
rect 121800 28500 121900 28600
rect 121800 28600 121900 28700
rect 121800 28700 121900 28800
rect 121800 28800 121900 28900
rect 121800 28900 121900 29000
rect 121800 29000 121900 29100
rect 121800 29100 121900 29200
rect 121800 29200 121900 29300
rect 121800 33300 121900 33400
rect 121800 33400 121900 33500
rect 121800 33500 121900 33600
rect 121800 33600 121900 33700
rect 121800 33700 121900 33800
rect 121800 33800 121900 33900
rect 121800 33900 121900 34000
rect 121800 34000 121900 34100
rect 121800 34100 121900 34200
rect 121800 34200 121900 34300
rect 121800 34300 121900 34400
rect 121800 34400 121900 34500
rect 121800 34500 121900 34600
rect 121800 34600 121900 34700
rect 121800 34700 121900 34800
rect 121800 34800 121900 34900
rect 121800 34900 121900 35000
rect 121800 35000 121900 35100
rect 121800 35100 121900 35200
rect 121800 35200 121900 35300
rect 121800 35300 121900 35400
rect 121800 36700 121900 36800
rect 121800 36800 121900 36900
rect 121800 36900 121900 37000
rect 121800 37000 121900 37100
rect 121800 37100 121900 37200
rect 121800 37200 121900 37300
rect 121800 37300 121900 37400
rect 121800 37400 121900 37500
rect 121800 37500 121900 37600
rect 121800 37600 121900 37700
rect 121800 37700 121900 37800
rect 121800 37800 121900 37900
rect 121800 37900 121900 38000
rect 121800 38000 121900 38100
rect 121800 38100 121900 38200
rect 121800 38200 121900 38300
rect 121800 38300 121900 38400
rect 121900 27200 122000 27300
rect 121900 27300 122000 27400
rect 121900 27400 122000 27500
rect 121900 27500 122000 27600
rect 121900 27600 122000 27700
rect 121900 27700 122000 27800
rect 121900 27800 122000 27900
rect 121900 27900 122000 28000
rect 121900 28000 122000 28100
rect 121900 28100 122000 28200
rect 121900 28200 122000 28300
rect 121900 28300 122000 28400
rect 121900 28400 122000 28500
rect 121900 28500 122000 28600
rect 121900 28600 122000 28700
rect 121900 28700 122000 28800
rect 121900 28800 122000 28900
rect 121900 28900 122000 29000
rect 121900 29000 122000 29100
rect 121900 29100 122000 29200
rect 121900 29200 122000 29300
rect 121900 29300 122000 29400
rect 121900 33300 122000 33400
rect 121900 33400 122000 33500
rect 121900 33500 122000 33600
rect 121900 33600 122000 33700
rect 121900 33700 122000 33800
rect 121900 33800 122000 33900
rect 121900 33900 122000 34000
rect 121900 34000 122000 34100
rect 121900 34100 122000 34200
rect 121900 34200 122000 34300
rect 121900 34300 122000 34400
rect 121900 34400 122000 34500
rect 121900 34500 122000 34600
rect 121900 34600 122000 34700
rect 121900 34700 122000 34800
rect 121900 34800 122000 34900
rect 121900 34900 122000 35000
rect 121900 35000 122000 35100
rect 121900 35100 122000 35200
rect 121900 35200 122000 35300
rect 121900 35300 122000 35400
rect 121900 36800 122000 36900
rect 121900 36900 122000 37000
rect 121900 37000 122000 37100
rect 121900 37100 122000 37200
rect 121900 37200 122000 37300
rect 121900 37300 122000 37400
rect 121900 37400 122000 37500
rect 121900 37500 122000 37600
rect 121900 37600 122000 37700
rect 121900 37700 122000 37800
rect 121900 37800 122000 37900
rect 121900 37900 122000 38000
rect 121900 38000 122000 38100
rect 121900 38100 122000 38200
rect 121900 38200 122000 38300
rect 121900 38300 122000 38400
rect 122000 27300 122100 27400
rect 122000 27400 122100 27500
rect 122000 27500 122100 27600
rect 122000 27600 122100 27700
rect 122000 27700 122100 27800
rect 122000 27800 122100 27900
rect 122000 27900 122100 28000
rect 122000 28000 122100 28100
rect 122000 28100 122100 28200
rect 122000 28200 122100 28300
rect 122000 28300 122100 28400
rect 122000 28400 122100 28500
rect 122000 28500 122100 28600
rect 122000 28600 122100 28700
rect 122000 28700 122100 28800
rect 122000 28800 122100 28900
rect 122000 28900 122100 29000
rect 122000 29000 122100 29100
rect 122000 29100 122100 29200
rect 122000 29200 122100 29300
rect 122000 29300 122100 29400
rect 122000 29400 122100 29500
rect 122000 33100 122100 33200
rect 122000 33200 122100 33300
rect 122000 33300 122100 33400
rect 122000 33400 122100 33500
rect 122000 33500 122100 33600
rect 122000 33600 122100 33700
rect 122000 33700 122100 33800
rect 122000 33800 122100 33900
rect 122000 33900 122100 34000
rect 122000 34000 122100 34100
rect 122000 34100 122100 34200
rect 122000 34200 122100 34300
rect 122000 34300 122100 34400
rect 122000 34400 122100 34500
rect 122000 34500 122100 34600
rect 122000 34600 122100 34700
rect 122000 34700 122100 34800
rect 122000 34800 122100 34900
rect 122000 34900 122100 35000
rect 122000 35000 122100 35100
rect 122000 35100 122100 35200
rect 122000 35200 122100 35300
rect 122000 35300 122100 35400
rect 122000 36800 122100 36900
rect 122000 36900 122100 37000
rect 122000 37000 122100 37100
rect 122000 37100 122100 37200
rect 122000 37200 122100 37300
rect 122000 37300 122100 37400
rect 122000 37400 122100 37500
rect 122000 37500 122100 37600
rect 122000 37600 122100 37700
rect 122000 37700 122100 37800
rect 122000 37800 122100 37900
rect 122000 37900 122100 38000
rect 122000 38000 122100 38100
rect 122000 38100 122100 38200
rect 122000 38200 122100 38300
rect 122000 38300 122100 38400
rect 122100 27400 122200 27500
rect 122100 27500 122200 27600
rect 122100 27600 122200 27700
rect 122100 27700 122200 27800
rect 122100 27800 122200 27900
rect 122100 27900 122200 28000
rect 122100 28000 122200 28100
rect 122100 28100 122200 28200
rect 122100 28200 122200 28300
rect 122100 28300 122200 28400
rect 122100 28400 122200 28500
rect 122100 28500 122200 28600
rect 122100 28600 122200 28700
rect 122100 28700 122200 28800
rect 122100 28800 122200 28900
rect 122100 28900 122200 29000
rect 122100 29000 122200 29100
rect 122100 29100 122200 29200
rect 122100 29200 122200 29300
rect 122100 29300 122200 29400
rect 122100 29400 122200 29500
rect 122100 33000 122200 33100
rect 122100 33100 122200 33200
rect 122100 33200 122200 33300
rect 122100 33300 122200 33400
rect 122100 33400 122200 33500
rect 122100 33500 122200 33600
rect 122100 33600 122200 33700
rect 122100 33700 122200 33800
rect 122100 33800 122200 33900
rect 122100 33900 122200 34000
rect 122100 34000 122200 34100
rect 122100 34100 122200 34200
rect 122100 34200 122200 34300
rect 122100 34300 122200 34400
rect 122100 34400 122200 34500
rect 122100 34500 122200 34600
rect 122100 34600 122200 34700
rect 122100 34700 122200 34800
rect 122100 34800 122200 34900
rect 122100 34900 122200 35000
rect 122100 35000 122200 35100
rect 122100 35100 122200 35200
rect 122100 35200 122200 35300
rect 122100 36800 122200 36900
rect 122100 36900 122200 37000
rect 122100 37000 122200 37100
rect 122100 37100 122200 37200
rect 122100 37200 122200 37300
rect 122100 37300 122200 37400
rect 122100 37400 122200 37500
rect 122100 37500 122200 37600
rect 122100 37600 122200 37700
rect 122100 37700 122200 37800
rect 122100 37800 122200 37900
rect 122100 37900 122200 38000
rect 122100 38000 122200 38100
rect 122100 38100 122200 38200
rect 122100 38200 122200 38300
rect 122100 38300 122200 38400
rect 122200 27400 122300 27500
rect 122200 27500 122300 27600
rect 122200 27600 122300 27700
rect 122200 27700 122300 27800
rect 122200 27800 122300 27900
rect 122200 27900 122300 28000
rect 122200 28000 122300 28100
rect 122200 28100 122300 28200
rect 122200 28200 122300 28300
rect 122200 28300 122300 28400
rect 122200 28400 122300 28500
rect 122200 28500 122300 28600
rect 122200 28600 122300 28700
rect 122200 28700 122300 28800
rect 122200 28800 122300 28900
rect 122200 28900 122300 29000
rect 122200 29000 122300 29100
rect 122200 29100 122300 29200
rect 122200 29200 122300 29300
rect 122200 29300 122300 29400
rect 122200 29400 122300 29500
rect 122200 29500 122300 29600
rect 122200 32800 122300 32900
rect 122200 32900 122300 33000
rect 122200 33000 122300 33100
rect 122200 33100 122300 33200
rect 122200 33200 122300 33300
rect 122200 33300 122300 33400
rect 122200 33400 122300 33500
rect 122200 33500 122300 33600
rect 122200 33600 122300 33700
rect 122200 33700 122300 33800
rect 122200 33800 122300 33900
rect 122200 33900 122300 34000
rect 122200 34000 122300 34100
rect 122200 34100 122300 34200
rect 122200 34200 122300 34300
rect 122200 34300 122300 34400
rect 122200 34400 122300 34500
rect 122200 34500 122300 34600
rect 122200 34600 122300 34700
rect 122200 34700 122300 34800
rect 122200 34800 122300 34900
rect 122200 34900 122300 35000
rect 122200 35000 122300 35100
rect 122200 35100 122300 35200
rect 122200 35200 122300 35300
rect 122200 36900 122300 37000
rect 122200 37000 122300 37100
rect 122200 37100 122300 37200
rect 122200 37200 122300 37300
rect 122200 37300 122300 37400
rect 122200 37400 122300 37500
rect 122200 37500 122300 37600
rect 122200 37600 122300 37700
rect 122200 37700 122300 37800
rect 122200 37800 122300 37900
rect 122200 37900 122300 38000
rect 122200 38000 122300 38100
rect 122200 38100 122300 38200
rect 122200 38200 122300 38300
rect 122200 38300 122300 38400
rect 122300 27500 122400 27600
rect 122300 27600 122400 27700
rect 122300 27700 122400 27800
rect 122300 27800 122400 27900
rect 122300 27900 122400 28000
rect 122300 28000 122400 28100
rect 122300 28100 122400 28200
rect 122300 28200 122400 28300
rect 122300 28300 122400 28400
rect 122300 28400 122400 28500
rect 122300 28500 122400 28600
rect 122300 28600 122400 28700
rect 122300 28700 122400 28800
rect 122300 28800 122400 28900
rect 122300 28900 122400 29000
rect 122300 29000 122400 29100
rect 122300 29100 122400 29200
rect 122300 29200 122400 29300
rect 122300 29300 122400 29400
rect 122300 29400 122400 29500
rect 122300 29500 122400 29600
rect 122300 29600 122400 29700
rect 122300 32700 122400 32800
rect 122300 32800 122400 32900
rect 122300 32900 122400 33000
rect 122300 33000 122400 33100
rect 122300 33100 122400 33200
rect 122300 33200 122400 33300
rect 122300 33300 122400 33400
rect 122300 33400 122400 33500
rect 122300 33500 122400 33600
rect 122300 33600 122400 33700
rect 122300 33700 122400 33800
rect 122300 33800 122400 33900
rect 122300 33900 122400 34000
rect 122300 34000 122400 34100
rect 122300 34100 122400 34200
rect 122300 34200 122400 34300
rect 122300 34300 122400 34400
rect 122300 34400 122400 34500
rect 122300 34500 122400 34600
rect 122300 34600 122400 34700
rect 122300 34700 122400 34800
rect 122300 34800 122400 34900
rect 122300 34900 122400 35000
rect 122300 35000 122400 35100
rect 122300 35100 122400 35200
rect 122300 35200 122400 35300
rect 122300 36800 122400 36900
rect 122300 36900 122400 37000
rect 122300 37000 122400 37100
rect 122300 37100 122400 37200
rect 122300 37200 122400 37300
rect 122300 37300 122400 37400
rect 122300 37400 122400 37500
rect 122300 37500 122400 37600
rect 122300 37600 122400 37700
rect 122300 37700 122400 37800
rect 122300 37800 122400 37900
rect 122300 37900 122400 38000
rect 122300 38000 122400 38100
rect 122300 38100 122400 38200
rect 122300 38200 122400 38300
rect 122300 38300 122400 38400
rect 122400 27600 122500 27700
rect 122400 27700 122500 27800
rect 122400 27800 122500 27900
rect 122400 27900 122500 28000
rect 122400 28000 122500 28100
rect 122400 28100 122500 28200
rect 122400 28200 122500 28300
rect 122400 28300 122500 28400
rect 122400 28400 122500 28500
rect 122400 28500 122500 28600
rect 122400 28600 122500 28700
rect 122400 28700 122500 28800
rect 122400 28800 122500 28900
rect 122400 28900 122500 29000
rect 122400 29000 122500 29100
rect 122400 29100 122500 29200
rect 122400 29200 122500 29300
rect 122400 29300 122500 29400
rect 122400 29400 122500 29500
rect 122400 29500 122500 29600
rect 122400 29600 122500 29700
rect 122400 29700 122500 29800
rect 122400 32500 122500 32600
rect 122400 32600 122500 32700
rect 122400 32700 122500 32800
rect 122400 32800 122500 32900
rect 122400 32900 122500 33000
rect 122400 33000 122500 33100
rect 122400 33100 122500 33200
rect 122400 33200 122500 33300
rect 122400 33300 122500 33400
rect 122400 33400 122500 33500
rect 122400 33500 122500 33600
rect 122400 33600 122500 33700
rect 122400 33700 122500 33800
rect 122400 33800 122500 33900
rect 122400 33900 122500 34000
rect 122400 34000 122500 34100
rect 122400 34100 122500 34200
rect 122400 34200 122500 34300
rect 122400 34300 122500 34400
rect 122400 34400 122500 34500
rect 122400 34500 122500 34600
rect 122400 34600 122500 34700
rect 122400 34700 122500 34800
rect 122400 34800 122500 34900
rect 122400 34900 122500 35000
rect 122400 35000 122500 35100
rect 122400 35100 122500 35200
rect 122400 35200 122500 35300
rect 122400 36800 122500 36900
rect 122400 36900 122500 37000
rect 122400 37000 122500 37100
rect 122400 37100 122500 37200
rect 122400 37200 122500 37300
rect 122400 37300 122500 37400
rect 122400 37400 122500 37500
rect 122400 37500 122500 37600
rect 122400 37600 122500 37700
rect 122400 37700 122500 37800
rect 122400 37800 122500 37900
rect 122400 37900 122500 38000
rect 122400 38000 122500 38100
rect 122400 38100 122500 38200
rect 122400 38200 122500 38300
rect 122400 38300 122500 38400
rect 122500 27700 122600 27800
rect 122500 27800 122600 27900
rect 122500 27900 122600 28000
rect 122500 28000 122600 28100
rect 122500 28100 122600 28200
rect 122500 28200 122600 28300
rect 122500 28300 122600 28400
rect 122500 28400 122600 28500
rect 122500 28500 122600 28600
rect 122500 28600 122600 28700
rect 122500 28700 122600 28800
rect 122500 28800 122600 28900
rect 122500 28900 122600 29000
rect 122500 29000 122600 29100
rect 122500 29100 122600 29200
rect 122500 29200 122600 29300
rect 122500 29300 122600 29400
rect 122500 29400 122600 29500
rect 122500 29500 122600 29600
rect 122500 29600 122600 29700
rect 122500 29700 122600 29800
rect 122500 32200 122600 32300
rect 122500 32300 122600 32400
rect 122500 32400 122600 32500
rect 122500 32500 122600 32600
rect 122500 32600 122600 32700
rect 122500 32700 122600 32800
rect 122500 32800 122600 32900
rect 122500 32900 122600 33000
rect 122500 33000 122600 33100
rect 122500 33100 122600 33200
rect 122500 33200 122600 33300
rect 122500 33300 122600 33400
rect 122500 33400 122600 33500
rect 122500 33500 122600 33600
rect 122500 33600 122600 33700
rect 122500 33700 122600 33800
rect 122500 33800 122600 33900
rect 122500 33900 122600 34000
rect 122500 34000 122600 34100
rect 122500 34100 122600 34200
rect 122500 34200 122600 34300
rect 122500 34300 122600 34400
rect 122500 34400 122600 34500
rect 122500 34500 122600 34600
rect 122500 34600 122600 34700
rect 122500 34700 122600 34800
rect 122500 34800 122600 34900
rect 122500 34900 122600 35000
rect 122500 35000 122600 35100
rect 122500 35100 122600 35200
rect 122500 35200 122600 35300
rect 122500 36800 122600 36900
rect 122500 36900 122600 37000
rect 122500 37000 122600 37100
rect 122500 37100 122600 37200
rect 122500 37200 122600 37300
rect 122500 37300 122600 37400
rect 122500 37400 122600 37500
rect 122500 37500 122600 37600
rect 122500 37600 122600 37700
rect 122500 37700 122600 37800
rect 122500 37800 122600 37900
rect 122500 37900 122600 38000
rect 122500 38000 122600 38100
rect 122500 38100 122600 38200
rect 122500 38200 122600 38300
rect 122500 38300 122600 38400
rect 122600 27800 122700 27900
rect 122600 27900 122700 28000
rect 122600 28000 122700 28100
rect 122600 28100 122700 28200
rect 122600 28200 122700 28300
rect 122600 28300 122700 28400
rect 122600 28400 122700 28500
rect 122600 28500 122700 28600
rect 122600 28600 122700 28700
rect 122600 28700 122700 28800
rect 122600 28800 122700 28900
rect 122600 28900 122700 29000
rect 122600 29000 122700 29100
rect 122600 29100 122700 29200
rect 122600 29200 122700 29300
rect 122600 29300 122700 29400
rect 122600 29400 122700 29500
rect 122600 29500 122700 29600
rect 122600 29600 122700 29700
rect 122600 29700 122700 29800
rect 122600 29800 122700 29900
rect 122600 32000 122700 32100
rect 122600 32100 122700 32200
rect 122600 32200 122700 32300
rect 122600 32300 122700 32400
rect 122600 32400 122700 32500
rect 122600 32500 122700 32600
rect 122600 32600 122700 32700
rect 122600 32700 122700 32800
rect 122600 32800 122700 32900
rect 122600 32900 122700 33000
rect 122600 33000 122700 33100
rect 122600 33100 122700 33200
rect 122600 33200 122700 33300
rect 122600 33300 122700 33400
rect 122600 33400 122700 33500
rect 122600 33500 122700 33600
rect 122600 33600 122700 33700
rect 122600 33700 122700 33800
rect 122600 33800 122700 33900
rect 122600 33900 122700 34000
rect 122600 34000 122700 34100
rect 122600 34100 122700 34200
rect 122600 34200 122700 34300
rect 122600 34300 122700 34400
rect 122600 34400 122700 34500
rect 122600 34500 122700 34600
rect 122600 34600 122700 34700
rect 122600 34700 122700 34800
rect 122600 34800 122700 34900
rect 122600 34900 122700 35000
rect 122600 35000 122700 35100
rect 122600 35100 122700 35200
rect 122600 35200 122700 35300
rect 122600 36700 122700 36800
rect 122600 36800 122700 36900
rect 122600 36900 122700 37000
rect 122600 37000 122700 37100
rect 122600 37100 122700 37200
rect 122600 37200 122700 37300
rect 122600 37300 122700 37400
rect 122600 37400 122700 37500
rect 122600 37500 122700 37600
rect 122600 37600 122700 37700
rect 122600 37700 122700 37800
rect 122600 37800 122700 37900
rect 122600 37900 122700 38000
rect 122600 38000 122700 38100
rect 122600 38100 122700 38200
rect 122600 38200 122700 38300
rect 122600 38300 122700 38400
rect 122700 27800 122800 27900
rect 122700 27900 122800 28000
rect 122700 28000 122800 28100
rect 122700 28100 122800 28200
rect 122700 28200 122800 28300
rect 122700 28300 122800 28400
rect 122700 28400 122800 28500
rect 122700 28500 122800 28600
rect 122700 28600 122800 28700
rect 122700 28700 122800 28800
rect 122700 28800 122800 28900
rect 122700 28900 122800 29000
rect 122700 29000 122800 29100
rect 122700 29100 122800 29200
rect 122700 29200 122800 29300
rect 122700 29300 122800 29400
rect 122700 29400 122800 29500
rect 122700 29500 122800 29600
rect 122700 29600 122800 29700
rect 122700 29700 122800 29800
rect 122700 29800 122800 29900
rect 122700 29900 122800 30000
rect 122700 31800 122800 31900
rect 122700 31900 122800 32000
rect 122700 32000 122800 32100
rect 122700 32100 122800 32200
rect 122700 32200 122800 32300
rect 122700 32300 122800 32400
rect 122700 32400 122800 32500
rect 122700 32500 122800 32600
rect 122700 32600 122800 32700
rect 122700 32700 122800 32800
rect 122700 32800 122800 32900
rect 122700 32900 122800 33000
rect 122700 33000 122800 33100
rect 122700 33100 122800 33200
rect 122700 33200 122800 33300
rect 122700 33300 122800 33400
rect 122700 33400 122800 33500
rect 122700 33500 122800 33600
rect 122700 33600 122800 33700
rect 122700 33700 122800 33800
rect 122700 33800 122800 33900
rect 122700 33900 122800 34000
rect 122700 34000 122800 34100
rect 122700 34100 122800 34200
rect 122700 34200 122800 34300
rect 122700 34300 122800 34400
rect 122700 34400 122800 34500
rect 122700 34500 122800 34600
rect 122700 34600 122800 34700
rect 122700 34700 122800 34800
rect 122700 34800 122800 34900
rect 122700 34900 122800 35000
rect 122700 35000 122800 35100
rect 122700 35100 122800 35200
rect 122700 35200 122800 35300
rect 122700 35300 122800 35400
rect 122700 36500 122800 36600
rect 122700 36600 122800 36700
rect 122700 36700 122800 36800
rect 122700 36800 122800 36900
rect 122700 36900 122800 37000
rect 122700 37000 122800 37100
rect 122700 37100 122800 37200
rect 122700 37200 122800 37300
rect 122700 37300 122800 37400
rect 122700 37400 122800 37500
rect 122700 37500 122800 37600
rect 122700 37600 122800 37700
rect 122700 37700 122800 37800
rect 122700 37800 122800 37900
rect 122700 37900 122800 38000
rect 122700 38000 122800 38100
rect 122700 38100 122800 38200
rect 122700 38200 122800 38300
rect 122700 38300 122800 38400
rect 122800 27900 122900 28000
rect 122800 28000 122900 28100
rect 122800 28100 122900 28200
rect 122800 28200 122900 28300
rect 122800 28300 122900 28400
rect 122800 28400 122900 28500
rect 122800 28500 122900 28600
rect 122800 28600 122900 28700
rect 122800 28700 122900 28800
rect 122800 28800 122900 28900
rect 122800 28900 122900 29000
rect 122800 29000 122900 29100
rect 122800 29100 122900 29200
rect 122800 29200 122900 29300
rect 122800 29300 122900 29400
rect 122800 29400 122900 29500
rect 122800 29500 122900 29600
rect 122800 29600 122900 29700
rect 122800 29700 122900 29800
rect 122800 29800 122900 29900
rect 122800 29900 122900 30000
rect 122800 30000 122900 30100
rect 122800 31500 122900 31600
rect 122800 31600 122900 31700
rect 122800 31700 122900 31800
rect 122800 31800 122900 31900
rect 122800 31900 122900 32000
rect 122800 32000 122900 32100
rect 122800 32100 122900 32200
rect 122800 32200 122900 32300
rect 122800 32300 122900 32400
rect 122800 32400 122900 32500
rect 122800 32500 122900 32600
rect 122800 32600 122900 32700
rect 122800 32700 122900 32800
rect 122800 32800 122900 32900
rect 122800 32900 122900 33000
rect 122800 33000 122900 33100
rect 122800 33100 122900 33200
rect 122800 33200 122900 33300
rect 122800 33300 122900 33400
rect 122800 33400 122900 33500
rect 122800 33500 122900 33600
rect 122800 33600 122900 33700
rect 122800 33700 122900 33800
rect 122800 33800 122900 33900
rect 122800 33900 122900 34000
rect 122800 34000 122900 34100
rect 122800 34100 122900 34200
rect 122800 34200 122900 34300
rect 122800 34300 122900 34400
rect 122800 34400 122900 34500
rect 122800 34500 122900 34600
rect 122800 34600 122900 34700
rect 122800 34700 122900 34800
rect 122800 34800 122900 34900
rect 122800 34900 122900 35000
rect 122800 35000 122900 35100
rect 122800 35100 122900 35200
rect 122800 35200 122900 35300
rect 122800 35300 122900 35400
rect 122800 35400 122900 35500
rect 122800 36300 122900 36400
rect 122800 36400 122900 36500
rect 122800 36500 122900 36600
rect 122800 36600 122900 36700
rect 122800 36700 122900 36800
rect 122800 36800 122900 36900
rect 122800 36900 122900 37000
rect 122800 37000 122900 37100
rect 122800 37100 122900 37200
rect 122800 37200 122900 37300
rect 122800 37300 122900 37400
rect 122800 37400 122900 37500
rect 122800 37500 122900 37600
rect 122800 37600 122900 37700
rect 122800 37700 122900 37800
rect 122800 37800 122900 37900
rect 122800 37900 122900 38000
rect 122800 38000 122900 38100
rect 122800 38100 122900 38200
rect 122800 38200 122900 38300
rect 122900 28000 123000 28100
rect 122900 28100 123000 28200
rect 122900 28200 123000 28300
rect 122900 28300 123000 28400
rect 122900 28400 123000 28500
rect 122900 28500 123000 28600
rect 122900 28600 123000 28700
rect 122900 28700 123000 28800
rect 122900 28800 123000 28900
rect 122900 28900 123000 29000
rect 122900 29000 123000 29100
rect 122900 29100 123000 29200
rect 122900 29200 123000 29300
rect 122900 29300 123000 29400
rect 122900 29400 123000 29500
rect 122900 29500 123000 29600
rect 122900 29600 123000 29700
rect 122900 29700 123000 29800
rect 122900 29800 123000 29900
rect 122900 29900 123000 30000
rect 122900 30000 123000 30100
rect 122900 31200 123000 31300
rect 122900 31300 123000 31400
rect 122900 31400 123000 31500
rect 122900 31500 123000 31600
rect 122900 31600 123000 31700
rect 122900 31700 123000 31800
rect 122900 31800 123000 31900
rect 122900 31900 123000 32000
rect 122900 32000 123000 32100
rect 122900 32100 123000 32200
rect 122900 32200 123000 32300
rect 122900 32300 123000 32400
rect 122900 32400 123000 32500
rect 122900 32500 123000 32600
rect 122900 32600 123000 32700
rect 122900 32700 123000 32800
rect 122900 32800 123000 32900
rect 122900 32900 123000 33000
rect 122900 33000 123000 33100
rect 122900 33100 123000 33200
rect 122900 33200 123000 33300
rect 122900 33300 123000 33400
rect 122900 33400 123000 33500
rect 122900 33500 123000 33600
rect 122900 33600 123000 33700
rect 122900 33700 123000 33800
rect 122900 33800 123000 33900
rect 122900 33900 123000 34000
rect 122900 34000 123000 34100
rect 122900 34100 123000 34200
rect 122900 34200 123000 34300
rect 122900 34300 123000 34400
rect 122900 34400 123000 34500
rect 122900 34500 123000 34600
rect 122900 34600 123000 34700
rect 122900 34700 123000 34800
rect 122900 34800 123000 34900
rect 122900 34900 123000 35000
rect 122900 35000 123000 35100
rect 122900 35100 123000 35200
rect 122900 35200 123000 35300
rect 122900 35300 123000 35400
rect 122900 35400 123000 35500
rect 122900 35500 123000 35600
rect 122900 35600 123000 35700
rect 122900 35700 123000 35800
rect 122900 35800 123000 35900
rect 122900 35900 123000 36000
rect 122900 36000 123000 36100
rect 122900 36100 123000 36200
rect 122900 36200 123000 36300
rect 122900 36300 123000 36400
rect 122900 36400 123000 36500
rect 122900 36500 123000 36600
rect 122900 36600 123000 36700
rect 122900 36700 123000 36800
rect 122900 36800 123000 36900
rect 122900 36900 123000 37000
rect 122900 37000 123000 37100
rect 122900 37100 123000 37200
rect 122900 37200 123000 37300
rect 122900 37300 123000 37400
rect 122900 37400 123000 37500
rect 122900 37500 123000 37600
rect 122900 37600 123000 37700
rect 122900 37700 123000 37800
rect 122900 37800 123000 37900
rect 122900 37900 123000 38000
rect 122900 38000 123000 38100
rect 122900 38100 123000 38200
rect 122900 38200 123000 38300
rect 123000 28000 123100 28100
rect 123000 28100 123100 28200
rect 123000 28200 123100 28300
rect 123000 28300 123100 28400
rect 123000 28400 123100 28500
rect 123000 28500 123100 28600
rect 123000 28600 123100 28700
rect 123000 28700 123100 28800
rect 123000 28800 123100 28900
rect 123000 28900 123100 29000
rect 123000 29000 123100 29100
rect 123000 29100 123100 29200
rect 123000 29200 123100 29300
rect 123000 29300 123100 29400
rect 123000 29400 123100 29500
rect 123000 29500 123100 29600
rect 123000 29600 123100 29700
rect 123000 29700 123100 29800
rect 123000 29800 123100 29900
rect 123000 29900 123100 30000
rect 123000 30000 123100 30100
rect 123000 30100 123100 30200
rect 123000 30900 123100 31000
rect 123000 31000 123100 31100
rect 123000 31100 123100 31200
rect 123000 31200 123100 31300
rect 123000 31300 123100 31400
rect 123000 31400 123100 31500
rect 123000 31500 123100 31600
rect 123000 31600 123100 31700
rect 123000 31700 123100 31800
rect 123000 31800 123100 31900
rect 123000 31900 123100 32000
rect 123000 32000 123100 32100
rect 123000 32100 123100 32200
rect 123000 32200 123100 32300
rect 123000 32300 123100 32400
rect 123000 32400 123100 32500
rect 123000 32500 123100 32600
rect 123000 32600 123100 32700
rect 123000 32700 123100 32800
rect 123000 32800 123100 32900
rect 123000 32900 123100 33000
rect 123000 33000 123100 33100
rect 123000 33100 123100 33200
rect 123000 33200 123100 33300
rect 123000 33300 123100 33400
rect 123000 33400 123100 33500
rect 123000 33500 123100 33600
rect 123000 33600 123100 33700
rect 123000 33700 123100 33800
rect 123000 33800 123100 33900
rect 123000 33900 123100 34000
rect 123000 34000 123100 34100
rect 123000 34100 123100 34200
rect 123000 34200 123100 34300
rect 123000 34300 123100 34400
rect 123000 34400 123100 34500
rect 123000 34500 123100 34600
rect 123000 34600 123100 34700
rect 123000 34700 123100 34800
rect 123000 34800 123100 34900
rect 123000 34900 123100 35000
rect 123000 35000 123100 35100
rect 123000 35100 123100 35200
rect 123000 35200 123100 35300
rect 123000 35300 123100 35400
rect 123000 35400 123100 35500
rect 123000 35500 123100 35600
rect 123000 35600 123100 35700
rect 123000 35700 123100 35800
rect 123000 35800 123100 35900
rect 123000 35900 123100 36000
rect 123000 36000 123100 36100
rect 123000 36100 123100 36200
rect 123000 36200 123100 36300
rect 123000 36300 123100 36400
rect 123000 36400 123100 36500
rect 123000 36500 123100 36600
rect 123000 36600 123100 36700
rect 123000 36700 123100 36800
rect 123000 36800 123100 36900
rect 123000 36900 123100 37000
rect 123000 37000 123100 37100
rect 123000 37100 123100 37200
rect 123000 37200 123100 37300
rect 123000 37300 123100 37400
rect 123000 37400 123100 37500
rect 123000 37500 123100 37600
rect 123000 37600 123100 37700
rect 123000 37700 123100 37800
rect 123000 37800 123100 37900
rect 123000 37900 123100 38000
rect 123000 38000 123100 38100
rect 123000 38100 123100 38200
rect 123000 38200 123100 38300
rect 123100 28100 123200 28200
rect 123100 28200 123200 28300
rect 123100 28300 123200 28400
rect 123100 28400 123200 28500
rect 123100 28500 123200 28600
rect 123100 28600 123200 28700
rect 123100 28700 123200 28800
rect 123100 28800 123200 28900
rect 123100 28900 123200 29000
rect 123100 29000 123200 29100
rect 123100 29100 123200 29200
rect 123100 29200 123200 29300
rect 123100 29300 123200 29400
rect 123100 29400 123200 29500
rect 123100 29500 123200 29600
rect 123100 29600 123200 29700
rect 123100 29700 123200 29800
rect 123100 29800 123200 29900
rect 123100 29900 123200 30000
rect 123100 30000 123200 30100
rect 123100 30100 123200 30200
rect 123100 30200 123200 30300
rect 123100 30700 123200 30800
rect 123100 30800 123200 30900
rect 123100 30900 123200 31000
rect 123100 31000 123200 31100
rect 123100 31100 123200 31200
rect 123100 31200 123200 31300
rect 123100 31300 123200 31400
rect 123100 31400 123200 31500
rect 123100 31500 123200 31600
rect 123100 31600 123200 31700
rect 123100 31700 123200 31800
rect 123100 31800 123200 31900
rect 123100 31900 123200 32000
rect 123100 32000 123200 32100
rect 123100 32100 123200 32200
rect 123100 32200 123200 32300
rect 123100 32300 123200 32400
rect 123100 32400 123200 32500
rect 123100 32500 123200 32600
rect 123100 32600 123200 32700
rect 123100 32700 123200 32800
rect 123100 32800 123200 32900
rect 123100 32900 123200 33000
rect 123100 33000 123200 33100
rect 123100 33100 123200 33200
rect 123100 33200 123200 33300
rect 123100 33300 123200 33400
rect 123100 33400 123200 33500
rect 123100 33500 123200 33600
rect 123100 33600 123200 33700
rect 123100 33700 123200 33800
rect 123100 33800 123200 33900
rect 123100 33900 123200 34000
rect 123100 34000 123200 34100
rect 123100 34100 123200 34200
rect 123100 34200 123200 34300
rect 123100 34300 123200 34400
rect 123100 34400 123200 34500
rect 123100 34500 123200 34600
rect 123100 34600 123200 34700
rect 123100 34700 123200 34800
rect 123100 34800 123200 34900
rect 123100 34900 123200 35000
rect 123100 35000 123200 35100
rect 123100 35100 123200 35200
rect 123100 35200 123200 35300
rect 123100 35300 123200 35400
rect 123100 35400 123200 35500
rect 123100 35500 123200 35600
rect 123100 35600 123200 35700
rect 123100 35700 123200 35800
rect 123100 35800 123200 35900
rect 123100 35900 123200 36000
rect 123100 36000 123200 36100
rect 123100 36100 123200 36200
rect 123100 36200 123200 36300
rect 123100 36300 123200 36400
rect 123100 36400 123200 36500
rect 123100 36500 123200 36600
rect 123100 36600 123200 36700
rect 123100 36700 123200 36800
rect 123100 36800 123200 36900
rect 123100 36900 123200 37000
rect 123100 37000 123200 37100
rect 123100 37100 123200 37200
rect 123100 37200 123200 37300
rect 123100 37300 123200 37400
rect 123100 37400 123200 37500
rect 123100 37500 123200 37600
rect 123100 37600 123200 37700
rect 123100 37700 123200 37800
rect 123100 37800 123200 37900
rect 123100 37900 123200 38000
rect 123100 38000 123200 38100
rect 123100 38100 123200 38200
rect 123200 28200 123300 28300
rect 123200 28300 123300 28400
rect 123200 28400 123300 28500
rect 123200 28500 123300 28600
rect 123200 28600 123300 28700
rect 123200 28700 123300 28800
rect 123200 28800 123300 28900
rect 123200 28900 123300 29000
rect 123200 29000 123300 29100
rect 123200 29100 123300 29200
rect 123200 29200 123300 29300
rect 123200 29300 123300 29400
rect 123200 29400 123300 29500
rect 123200 29500 123300 29600
rect 123200 29600 123300 29700
rect 123200 29700 123300 29800
rect 123200 29800 123300 29900
rect 123200 29900 123300 30000
rect 123200 30000 123300 30100
rect 123200 30100 123300 30200
rect 123200 30200 123300 30300
rect 123200 30300 123300 30400
rect 123200 30400 123300 30500
rect 123200 30500 123300 30600
rect 123200 30600 123300 30700
rect 123200 30700 123300 30800
rect 123200 30800 123300 30900
rect 123200 30900 123300 31000
rect 123200 31000 123300 31100
rect 123200 31100 123300 31200
rect 123200 31200 123300 31300
rect 123200 31300 123300 31400
rect 123200 31400 123300 31500
rect 123200 31500 123300 31600
rect 123200 31600 123300 31700
rect 123200 31700 123300 31800
rect 123200 31800 123300 31900
rect 123200 31900 123300 32000
rect 123200 32000 123300 32100
rect 123200 32100 123300 32200
rect 123200 32200 123300 32300
rect 123200 32300 123300 32400
rect 123200 32400 123300 32500
rect 123200 32500 123300 32600
rect 123200 32600 123300 32700
rect 123200 32700 123300 32800
rect 123200 32800 123300 32900
rect 123200 32900 123300 33000
rect 123200 33000 123300 33100
rect 123200 33100 123300 33200
rect 123200 33200 123300 33300
rect 123200 33300 123300 33400
rect 123200 33400 123300 33500
rect 123200 33500 123300 33600
rect 123200 33600 123300 33700
rect 123200 33700 123300 33800
rect 123200 33800 123300 33900
rect 123200 33900 123300 34000
rect 123200 34000 123300 34100
rect 123200 34100 123300 34200
rect 123200 34200 123300 34300
rect 123200 34300 123300 34400
rect 123200 34400 123300 34500
rect 123200 34500 123300 34600
rect 123200 34600 123300 34700
rect 123200 34700 123300 34800
rect 123200 34800 123300 34900
rect 123200 34900 123300 35000
rect 123200 35000 123300 35100
rect 123200 35100 123300 35200
rect 123200 35200 123300 35300
rect 123200 35300 123300 35400
rect 123200 35400 123300 35500
rect 123200 35500 123300 35600
rect 123200 35600 123300 35700
rect 123200 35700 123300 35800
rect 123200 35800 123300 35900
rect 123200 35900 123300 36000
rect 123200 36000 123300 36100
rect 123200 36100 123300 36200
rect 123200 36200 123300 36300
rect 123200 36300 123300 36400
rect 123200 36400 123300 36500
rect 123200 36500 123300 36600
rect 123200 36600 123300 36700
rect 123200 36700 123300 36800
rect 123200 36800 123300 36900
rect 123200 36900 123300 37000
rect 123200 37000 123300 37100
rect 123200 37100 123300 37200
rect 123200 37200 123300 37300
rect 123200 37300 123300 37400
rect 123200 37400 123300 37500
rect 123200 37500 123300 37600
rect 123200 37600 123300 37700
rect 123200 37700 123300 37800
rect 123200 37800 123300 37900
rect 123200 37900 123300 38000
rect 123200 38000 123300 38100
rect 123200 38100 123300 38200
rect 123300 28200 123400 28300
rect 123300 28300 123400 28400
rect 123300 28400 123400 28500
rect 123300 28500 123400 28600
rect 123300 28600 123400 28700
rect 123300 28700 123400 28800
rect 123300 28800 123400 28900
rect 123300 28900 123400 29000
rect 123300 29000 123400 29100
rect 123300 29100 123400 29200
rect 123300 29200 123400 29300
rect 123300 29300 123400 29400
rect 123300 29400 123400 29500
rect 123300 29500 123400 29600
rect 123300 29600 123400 29700
rect 123300 29700 123400 29800
rect 123300 29800 123400 29900
rect 123300 29900 123400 30000
rect 123300 30000 123400 30100
rect 123300 30100 123400 30200
rect 123300 30200 123400 30300
rect 123300 30300 123400 30400
rect 123300 30400 123400 30500
rect 123300 30500 123400 30600
rect 123300 30600 123400 30700
rect 123300 30700 123400 30800
rect 123300 30800 123400 30900
rect 123300 30900 123400 31000
rect 123300 31000 123400 31100
rect 123300 31100 123400 31200
rect 123300 31200 123400 31300
rect 123300 31300 123400 31400
rect 123300 31400 123400 31500
rect 123300 31500 123400 31600
rect 123300 31600 123400 31700
rect 123300 31700 123400 31800
rect 123300 31800 123400 31900
rect 123300 31900 123400 32000
rect 123300 32000 123400 32100
rect 123300 32100 123400 32200
rect 123300 32200 123400 32300
rect 123300 32300 123400 32400
rect 123300 32400 123400 32500
rect 123300 32500 123400 32600
rect 123300 32600 123400 32700
rect 123300 32700 123400 32800
rect 123300 32800 123400 32900
rect 123300 32900 123400 33000
rect 123300 33000 123400 33100
rect 123300 33100 123400 33200
rect 123300 33200 123400 33300
rect 123300 33300 123400 33400
rect 123300 33400 123400 33500
rect 123300 33500 123400 33600
rect 123300 33600 123400 33700
rect 123300 33700 123400 33800
rect 123300 33800 123400 33900
rect 123300 33900 123400 34000
rect 123300 34000 123400 34100
rect 123300 34100 123400 34200
rect 123300 34200 123400 34300
rect 123300 34300 123400 34400
rect 123300 34400 123400 34500
rect 123300 34500 123400 34600
rect 123300 34600 123400 34700
rect 123300 34700 123400 34800
rect 123300 34800 123400 34900
rect 123300 34900 123400 35000
rect 123300 35000 123400 35100
rect 123300 35100 123400 35200
rect 123300 35200 123400 35300
rect 123300 35300 123400 35400
rect 123300 35400 123400 35500
rect 123300 35500 123400 35600
rect 123300 35600 123400 35700
rect 123300 35700 123400 35800
rect 123300 35800 123400 35900
rect 123300 35900 123400 36000
rect 123300 36000 123400 36100
rect 123300 36100 123400 36200
rect 123300 36200 123400 36300
rect 123300 36300 123400 36400
rect 123300 36400 123400 36500
rect 123300 36500 123400 36600
rect 123300 36600 123400 36700
rect 123300 36700 123400 36800
rect 123300 36800 123400 36900
rect 123300 36900 123400 37000
rect 123300 37000 123400 37100
rect 123300 37100 123400 37200
rect 123300 37200 123400 37300
rect 123300 37300 123400 37400
rect 123300 37400 123400 37500
rect 123300 37500 123400 37600
rect 123300 37600 123400 37700
rect 123300 37700 123400 37800
rect 123300 37800 123400 37900
rect 123300 37900 123400 38000
rect 123300 38000 123400 38100
rect 123400 28300 123500 28400
rect 123400 28400 123500 28500
rect 123400 28500 123500 28600
rect 123400 28600 123500 28700
rect 123400 28700 123500 28800
rect 123400 28800 123500 28900
rect 123400 28900 123500 29000
rect 123400 29000 123500 29100
rect 123400 29100 123500 29200
rect 123400 29200 123500 29300
rect 123400 29300 123500 29400
rect 123400 29400 123500 29500
rect 123400 29500 123500 29600
rect 123400 29600 123500 29700
rect 123400 29700 123500 29800
rect 123400 29800 123500 29900
rect 123400 29900 123500 30000
rect 123400 30000 123500 30100
rect 123400 30100 123500 30200
rect 123400 30200 123500 30300
rect 123400 30300 123500 30400
rect 123400 30400 123500 30500
rect 123400 30500 123500 30600
rect 123400 30600 123500 30700
rect 123400 30700 123500 30800
rect 123400 30800 123500 30900
rect 123400 30900 123500 31000
rect 123400 31000 123500 31100
rect 123400 31100 123500 31200
rect 123400 31200 123500 31300
rect 123400 31300 123500 31400
rect 123400 31400 123500 31500
rect 123400 31500 123500 31600
rect 123400 31600 123500 31700
rect 123400 31700 123500 31800
rect 123400 31800 123500 31900
rect 123400 31900 123500 32000
rect 123400 32000 123500 32100
rect 123400 32100 123500 32200
rect 123400 32200 123500 32300
rect 123400 32300 123500 32400
rect 123400 32400 123500 32500
rect 123400 32500 123500 32600
rect 123400 32600 123500 32700
rect 123400 32700 123500 32800
rect 123400 32800 123500 32900
rect 123400 32900 123500 33000
rect 123400 33000 123500 33100
rect 123400 33100 123500 33200
rect 123400 33200 123500 33300
rect 123400 33300 123500 33400
rect 123400 33400 123500 33500
rect 123400 33500 123500 33600
rect 123400 33600 123500 33700
rect 123400 33700 123500 33800
rect 123400 33800 123500 33900
rect 123400 33900 123500 34000
rect 123400 34000 123500 34100
rect 123400 34100 123500 34200
rect 123400 34200 123500 34300
rect 123400 34300 123500 34400
rect 123400 34400 123500 34500
rect 123400 34500 123500 34600
rect 123400 34600 123500 34700
rect 123400 34700 123500 34800
rect 123400 34800 123500 34900
rect 123400 34900 123500 35000
rect 123400 35000 123500 35100
rect 123400 35100 123500 35200
rect 123400 35200 123500 35300
rect 123400 35300 123500 35400
rect 123400 35400 123500 35500
rect 123400 35500 123500 35600
rect 123400 35600 123500 35700
rect 123400 35700 123500 35800
rect 123400 35800 123500 35900
rect 123400 35900 123500 36000
rect 123400 36000 123500 36100
rect 123400 36100 123500 36200
rect 123400 36200 123500 36300
rect 123400 36300 123500 36400
rect 123400 36400 123500 36500
rect 123400 36500 123500 36600
rect 123400 36600 123500 36700
rect 123400 36700 123500 36800
rect 123400 36800 123500 36900
rect 123400 36900 123500 37000
rect 123400 37000 123500 37100
rect 123400 37100 123500 37200
rect 123400 37200 123500 37300
rect 123400 37300 123500 37400
rect 123400 37400 123500 37500
rect 123400 37500 123500 37600
rect 123400 37600 123500 37700
rect 123400 37700 123500 37800
rect 123400 37800 123500 37900
rect 123400 37900 123500 38000
rect 123400 38000 123500 38100
rect 123500 28300 123600 28400
rect 123500 28400 123600 28500
rect 123500 28500 123600 28600
rect 123500 28600 123600 28700
rect 123500 28700 123600 28800
rect 123500 28800 123600 28900
rect 123500 28900 123600 29000
rect 123500 29000 123600 29100
rect 123500 29100 123600 29200
rect 123500 29200 123600 29300
rect 123500 29300 123600 29400
rect 123500 29400 123600 29500
rect 123500 29500 123600 29600
rect 123500 29600 123600 29700
rect 123500 29700 123600 29800
rect 123500 29800 123600 29900
rect 123500 29900 123600 30000
rect 123500 30000 123600 30100
rect 123500 30100 123600 30200
rect 123500 30200 123600 30300
rect 123500 30300 123600 30400
rect 123500 30400 123600 30500
rect 123500 30500 123600 30600
rect 123500 30600 123600 30700
rect 123500 30700 123600 30800
rect 123500 30800 123600 30900
rect 123500 30900 123600 31000
rect 123500 31000 123600 31100
rect 123500 31100 123600 31200
rect 123500 31200 123600 31300
rect 123500 31300 123600 31400
rect 123500 31400 123600 31500
rect 123500 31500 123600 31600
rect 123500 31600 123600 31700
rect 123500 31700 123600 31800
rect 123500 31800 123600 31900
rect 123500 31900 123600 32000
rect 123500 32000 123600 32100
rect 123500 32100 123600 32200
rect 123500 32200 123600 32300
rect 123500 32300 123600 32400
rect 123500 32400 123600 32500
rect 123500 32500 123600 32600
rect 123500 32600 123600 32700
rect 123500 32700 123600 32800
rect 123500 32800 123600 32900
rect 123500 32900 123600 33000
rect 123500 33000 123600 33100
rect 123500 33100 123600 33200
rect 123500 33200 123600 33300
rect 123500 33300 123600 33400
rect 123500 33400 123600 33500
rect 123500 33500 123600 33600
rect 123500 33600 123600 33700
rect 123500 33700 123600 33800
rect 123500 33800 123600 33900
rect 123500 33900 123600 34000
rect 123500 34000 123600 34100
rect 123500 34100 123600 34200
rect 123500 34200 123600 34300
rect 123500 34300 123600 34400
rect 123500 34400 123600 34500
rect 123500 34500 123600 34600
rect 123500 34600 123600 34700
rect 123500 34700 123600 34800
rect 123500 34800 123600 34900
rect 123500 34900 123600 35000
rect 123500 35000 123600 35100
rect 123500 35100 123600 35200
rect 123500 35200 123600 35300
rect 123500 35300 123600 35400
rect 123500 35400 123600 35500
rect 123500 35500 123600 35600
rect 123500 35600 123600 35700
rect 123500 35700 123600 35800
rect 123500 35800 123600 35900
rect 123500 35900 123600 36000
rect 123500 36000 123600 36100
rect 123500 36100 123600 36200
rect 123500 36200 123600 36300
rect 123500 36300 123600 36400
rect 123500 36400 123600 36500
rect 123500 36500 123600 36600
rect 123500 36600 123600 36700
rect 123500 36700 123600 36800
rect 123500 36800 123600 36900
rect 123500 36900 123600 37000
rect 123500 37000 123600 37100
rect 123500 37100 123600 37200
rect 123500 37200 123600 37300
rect 123500 37300 123600 37400
rect 123500 37400 123600 37500
rect 123500 37500 123600 37600
rect 123500 37600 123600 37700
rect 123500 37700 123600 37800
rect 123500 37800 123600 37900
rect 123500 37900 123600 38000
rect 123600 28400 123700 28500
rect 123600 28500 123700 28600
rect 123600 28600 123700 28700
rect 123600 28700 123700 28800
rect 123600 28800 123700 28900
rect 123600 28900 123700 29000
rect 123600 29000 123700 29100
rect 123600 29100 123700 29200
rect 123600 29200 123700 29300
rect 123600 29300 123700 29400
rect 123600 29400 123700 29500
rect 123600 29500 123700 29600
rect 123600 29600 123700 29700
rect 123600 29700 123700 29800
rect 123600 29800 123700 29900
rect 123600 29900 123700 30000
rect 123600 30000 123700 30100
rect 123600 30100 123700 30200
rect 123600 30200 123700 30300
rect 123600 30300 123700 30400
rect 123600 30400 123700 30500
rect 123600 30500 123700 30600
rect 123600 30600 123700 30700
rect 123600 30700 123700 30800
rect 123600 30800 123700 30900
rect 123600 30900 123700 31000
rect 123600 31000 123700 31100
rect 123600 31100 123700 31200
rect 123600 31200 123700 31300
rect 123600 31300 123700 31400
rect 123600 31400 123700 31500
rect 123600 31500 123700 31600
rect 123600 31600 123700 31700
rect 123600 31700 123700 31800
rect 123600 31800 123700 31900
rect 123600 31900 123700 32000
rect 123600 32000 123700 32100
rect 123600 32100 123700 32200
rect 123600 32200 123700 32300
rect 123600 32300 123700 32400
rect 123600 32400 123700 32500
rect 123600 32500 123700 32600
rect 123600 32600 123700 32700
rect 123600 32700 123700 32800
rect 123600 32800 123700 32900
rect 123600 32900 123700 33000
rect 123600 33000 123700 33100
rect 123600 33100 123700 33200
rect 123600 33200 123700 33300
rect 123600 33300 123700 33400
rect 123600 33400 123700 33500
rect 123600 33500 123700 33600
rect 123600 33600 123700 33700
rect 123600 33700 123700 33800
rect 123600 33800 123700 33900
rect 123600 33900 123700 34000
rect 123600 34000 123700 34100
rect 123600 34100 123700 34200
rect 123600 34200 123700 34300
rect 123600 34300 123700 34400
rect 123600 34400 123700 34500
rect 123600 34500 123700 34600
rect 123600 34600 123700 34700
rect 123600 34700 123700 34800
rect 123600 34800 123700 34900
rect 123600 34900 123700 35000
rect 123600 35000 123700 35100
rect 123600 35100 123700 35200
rect 123600 35200 123700 35300
rect 123600 35300 123700 35400
rect 123600 35400 123700 35500
rect 123600 35500 123700 35600
rect 123600 35600 123700 35700
rect 123600 35700 123700 35800
rect 123600 35800 123700 35900
rect 123600 35900 123700 36000
rect 123600 36000 123700 36100
rect 123600 36100 123700 36200
rect 123600 36200 123700 36300
rect 123600 36300 123700 36400
rect 123600 36400 123700 36500
rect 123600 36500 123700 36600
rect 123600 36600 123700 36700
rect 123600 36700 123700 36800
rect 123600 36800 123700 36900
rect 123600 36900 123700 37000
rect 123600 37000 123700 37100
rect 123600 37100 123700 37200
rect 123600 37200 123700 37300
rect 123600 37300 123700 37400
rect 123600 37400 123700 37500
rect 123600 37500 123700 37600
rect 123600 37600 123700 37700
rect 123600 37700 123700 37800
rect 123600 37800 123700 37900
rect 123600 37900 123700 38000
rect 123700 28400 123800 28500
rect 123700 28500 123800 28600
rect 123700 28600 123800 28700
rect 123700 28700 123800 28800
rect 123700 28800 123800 28900
rect 123700 28900 123800 29000
rect 123700 29000 123800 29100
rect 123700 29100 123800 29200
rect 123700 29200 123800 29300
rect 123700 29300 123800 29400
rect 123700 29400 123800 29500
rect 123700 29500 123800 29600
rect 123700 29600 123800 29700
rect 123700 29700 123800 29800
rect 123700 29800 123800 29900
rect 123700 29900 123800 30000
rect 123700 30000 123800 30100
rect 123700 30100 123800 30200
rect 123700 30200 123800 30300
rect 123700 30300 123800 30400
rect 123700 30400 123800 30500
rect 123700 30500 123800 30600
rect 123700 30600 123800 30700
rect 123700 30700 123800 30800
rect 123700 30800 123800 30900
rect 123700 30900 123800 31000
rect 123700 31000 123800 31100
rect 123700 31100 123800 31200
rect 123700 31200 123800 31300
rect 123700 31300 123800 31400
rect 123700 31400 123800 31500
rect 123700 31500 123800 31600
rect 123700 31600 123800 31700
rect 123700 31700 123800 31800
rect 123700 31800 123800 31900
rect 123700 31900 123800 32000
rect 123700 32000 123800 32100
rect 123700 32100 123800 32200
rect 123700 32200 123800 32300
rect 123700 32300 123800 32400
rect 123700 32400 123800 32500
rect 123700 32500 123800 32600
rect 123700 32600 123800 32700
rect 123700 32700 123800 32800
rect 123700 32800 123800 32900
rect 123700 32900 123800 33000
rect 123700 33000 123800 33100
rect 123700 33100 123800 33200
rect 123700 33200 123800 33300
rect 123700 33300 123800 33400
rect 123700 33400 123800 33500
rect 123700 33500 123800 33600
rect 123700 33600 123800 33700
rect 123700 33700 123800 33800
rect 123700 33800 123800 33900
rect 123700 33900 123800 34000
rect 123700 34000 123800 34100
rect 123700 34100 123800 34200
rect 123700 34200 123800 34300
rect 123700 34300 123800 34400
rect 123700 34400 123800 34500
rect 123700 34500 123800 34600
rect 123700 34600 123800 34700
rect 123700 34700 123800 34800
rect 123700 34800 123800 34900
rect 123700 34900 123800 35000
rect 123700 35000 123800 35100
rect 123700 35100 123800 35200
rect 123700 35200 123800 35300
rect 123700 35300 123800 35400
rect 123700 35400 123800 35500
rect 123700 35500 123800 35600
rect 123700 35600 123800 35700
rect 123700 35700 123800 35800
rect 123700 35800 123800 35900
rect 123700 35900 123800 36000
rect 123700 36000 123800 36100
rect 123700 36100 123800 36200
rect 123700 36200 123800 36300
rect 123700 36300 123800 36400
rect 123700 36400 123800 36500
rect 123700 36500 123800 36600
rect 123700 36600 123800 36700
rect 123700 36700 123800 36800
rect 123700 36800 123800 36900
rect 123700 36900 123800 37000
rect 123700 37000 123800 37100
rect 123700 37100 123800 37200
rect 123700 37200 123800 37300
rect 123700 37300 123800 37400
rect 123700 37400 123800 37500
rect 123700 37500 123800 37600
rect 123700 37600 123800 37700
rect 123700 37700 123800 37800
rect 123700 37800 123800 37900
rect 123800 23800 123900 23900
rect 123800 23900 123900 24000
rect 123800 24000 123900 24100
rect 123800 24100 123900 24200
rect 123800 24200 123900 24300
rect 123800 24300 123900 24400
rect 123800 24400 123900 24500
rect 123800 24500 123900 24600
rect 123800 28500 123900 28600
rect 123800 28600 123900 28700
rect 123800 28700 123900 28800
rect 123800 28800 123900 28900
rect 123800 28900 123900 29000
rect 123800 29000 123900 29100
rect 123800 29100 123900 29200
rect 123800 29200 123900 29300
rect 123800 29300 123900 29400
rect 123800 29400 123900 29500
rect 123800 29500 123900 29600
rect 123800 29600 123900 29700
rect 123800 29700 123900 29800
rect 123800 29800 123900 29900
rect 123800 29900 123900 30000
rect 123800 30000 123900 30100
rect 123800 30100 123900 30200
rect 123800 30200 123900 30300
rect 123800 30300 123900 30400
rect 123800 30400 123900 30500
rect 123800 30500 123900 30600
rect 123800 30600 123900 30700
rect 123800 30700 123900 30800
rect 123800 30800 123900 30900
rect 123800 30900 123900 31000
rect 123800 31000 123900 31100
rect 123800 31100 123900 31200
rect 123800 31200 123900 31300
rect 123800 31300 123900 31400
rect 123800 31400 123900 31500
rect 123800 31500 123900 31600
rect 123800 31600 123900 31700
rect 123800 31700 123900 31800
rect 123800 31800 123900 31900
rect 123800 31900 123900 32000
rect 123800 32000 123900 32100
rect 123800 32100 123900 32200
rect 123800 32200 123900 32300
rect 123800 32300 123900 32400
rect 123800 32400 123900 32500
rect 123800 32500 123900 32600
rect 123800 32600 123900 32700
rect 123800 32700 123900 32800
rect 123800 32800 123900 32900
rect 123800 32900 123900 33000
rect 123800 33000 123900 33100
rect 123800 33100 123900 33200
rect 123800 33200 123900 33300
rect 123800 33300 123900 33400
rect 123800 33400 123900 33500
rect 123800 33500 123900 33600
rect 123800 33600 123900 33700
rect 123800 33700 123900 33800
rect 123800 33800 123900 33900
rect 123800 33900 123900 34000
rect 123800 34000 123900 34100
rect 123800 34100 123900 34200
rect 123800 34200 123900 34300
rect 123800 34300 123900 34400
rect 123800 34400 123900 34500
rect 123800 34500 123900 34600
rect 123800 34600 123900 34700
rect 123800 34700 123900 34800
rect 123800 34800 123900 34900
rect 123800 34900 123900 35000
rect 123800 35000 123900 35100
rect 123800 35100 123900 35200
rect 123800 35200 123900 35300
rect 123800 35300 123900 35400
rect 123800 35400 123900 35500
rect 123800 35500 123900 35600
rect 123800 35600 123900 35700
rect 123800 35700 123900 35800
rect 123800 35800 123900 35900
rect 123800 35900 123900 36000
rect 123800 36000 123900 36100
rect 123800 36100 123900 36200
rect 123800 36200 123900 36300
rect 123800 36300 123900 36400
rect 123800 36400 123900 36500
rect 123800 36500 123900 36600
rect 123800 36600 123900 36700
rect 123800 36700 123900 36800
rect 123800 36800 123900 36900
rect 123800 36900 123900 37000
rect 123800 37000 123900 37100
rect 123800 37100 123900 37200
rect 123800 37200 123900 37300
rect 123800 37300 123900 37400
rect 123800 37400 123900 37500
rect 123800 37500 123900 37600
rect 123800 37600 123900 37700
rect 123800 37700 123900 37800
rect 123900 23300 124000 23400
rect 123900 23400 124000 23500
rect 123900 23500 124000 23600
rect 123900 23600 124000 23700
rect 123900 23700 124000 23800
rect 123900 23800 124000 23900
rect 123900 23900 124000 24000
rect 123900 24000 124000 24100
rect 123900 24100 124000 24200
rect 123900 24200 124000 24300
rect 123900 24300 124000 24400
rect 123900 24400 124000 24500
rect 123900 24500 124000 24600
rect 123900 24600 124000 24700
rect 123900 24700 124000 24800
rect 123900 24800 124000 24900
rect 123900 24900 124000 25000
rect 123900 28300 124000 28400
rect 123900 28400 124000 28500
rect 123900 28500 124000 28600
rect 123900 28600 124000 28700
rect 123900 28700 124000 28800
rect 123900 28800 124000 28900
rect 123900 28900 124000 29000
rect 123900 29000 124000 29100
rect 123900 29100 124000 29200
rect 123900 29200 124000 29300
rect 123900 29300 124000 29400
rect 123900 29400 124000 29500
rect 123900 29500 124000 29600
rect 123900 29600 124000 29700
rect 123900 29700 124000 29800
rect 123900 29800 124000 29900
rect 123900 29900 124000 30000
rect 123900 30000 124000 30100
rect 123900 30100 124000 30200
rect 123900 30200 124000 30300
rect 123900 30300 124000 30400
rect 123900 30400 124000 30500
rect 123900 30500 124000 30600
rect 123900 30600 124000 30700
rect 123900 30700 124000 30800
rect 123900 30800 124000 30900
rect 123900 30900 124000 31000
rect 123900 31000 124000 31100
rect 123900 31100 124000 31200
rect 123900 31200 124000 31300
rect 123900 31300 124000 31400
rect 123900 31400 124000 31500
rect 123900 31500 124000 31600
rect 123900 31600 124000 31700
rect 123900 31700 124000 31800
rect 123900 31800 124000 31900
rect 123900 31900 124000 32000
rect 123900 32000 124000 32100
rect 123900 32100 124000 32200
rect 123900 32200 124000 32300
rect 123900 32300 124000 32400
rect 123900 32400 124000 32500
rect 123900 32500 124000 32600
rect 123900 32600 124000 32700
rect 123900 32700 124000 32800
rect 123900 32800 124000 32900
rect 123900 32900 124000 33000
rect 123900 33000 124000 33100
rect 123900 33100 124000 33200
rect 123900 33200 124000 33300
rect 123900 33300 124000 33400
rect 123900 33400 124000 33500
rect 123900 33500 124000 33600
rect 123900 33600 124000 33700
rect 123900 33700 124000 33800
rect 123900 33800 124000 33900
rect 123900 33900 124000 34000
rect 123900 34000 124000 34100
rect 123900 34100 124000 34200
rect 123900 34200 124000 34300
rect 123900 34300 124000 34400
rect 123900 34400 124000 34500
rect 123900 34500 124000 34600
rect 123900 34600 124000 34700
rect 123900 34700 124000 34800
rect 123900 34800 124000 34900
rect 123900 34900 124000 35000
rect 123900 35000 124000 35100
rect 123900 35100 124000 35200
rect 123900 35200 124000 35300
rect 123900 35300 124000 35400
rect 123900 35400 124000 35500
rect 123900 35500 124000 35600
rect 123900 35600 124000 35700
rect 123900 35700 124000 35800
rect 123900 35800 124000 35900
rect 123900 35900 124000 36000
rect 123900 36000 124000 36100
rect 123900 36100 124000 36200
rect 123900 36200 124000 36300
rect 123900 36300 124000 36400
rect 123900 36400 124000 36500
rect 123900 36500 124000 36600
rect 123900 36600 124000 36700
rect 123900 36700 124000 36800
rect 123900 36800 124000 36900
rect 123900 36900 124000 37000
rect 123900 37000 124000 37100
rect 123900 37100 124000 37200
rect 123900 37200 124000 37300
rect 123900 37300 124000 37400
rect 123900 37400 124000 37500
rect 123900 37500 124000 37600
rect 123900 37600 124000 37700
rect 124000 23100 124100 23200
rect 124000 23200 124100 23300
rect 124000 23300 124100 23400
rect 124000 23400 124100 23500
rect 124000 23500 124100 23600
rect 124000 23600 124100 23700
rect 124000 23700 124100 23800
rect 124000 23800 124100 23900
rect 124000 23900 124100 24000
rect 124000 24000 124100 24100
rect 124000 24100 124100 24200
rect 124000 24200 124100 24300
rect 124000 24300 124100 24400
rect 124000 24400 124100 24500
rect 124000 24500 124100 24600
rect 124000 24600 124100 24700
rect 124000 24700 124100 24800
rect 124000 24800 124100 24900
rect 124000 24900 124100 25000
rect 124000 25000 124100 25100
rect 124000 25100 124100 25200
rect 124000 25200 124100 25300
rect 124000 28000 124100 28100
rect 124000 28100 124100 28200
rect 124000 28200 124100 28300
rect 124000 28300 124100 28400
rect 124000 28400 124100 28500
rect 124000 28500 124100 28600
rect 124000 28600 124100 28700
rect 124000 28700 124100 28800
rect 124000 28800 124100 28900
rect 124000 28900 124100 29000
rect 124000 29000 124100 29100
rect 124000 29100 124100 29200
rect 124000 29200 124100 29300
rect 124000 29300 124100 29400
rect 124000 29400 124100 29500
rect 124000 29500 124100 29600
rect 124000 29600 124100 29700
rect 124000 29700 124100 29800
rect 124000 29800 124100 29900
rect 124000 29900 124100 30000
rect 124000 30000 124100 30100
rect 124000 30100 124100 30200
rect 124000 30200 124100 30300
rect 124000 30300 124100 30400
rect 124000 30400 124100 30500
rect 124000 30500 124100 30600
rect 124000 30600 124100 30700
rect 124000 30700 124100 30800
rect 124000 30800 124100 30900
rect 124000 30900 124100 31000
rect 124000 31000 124100 31100
rect 124000 31100 124100 31200
rect 124000 31200 124100 31300
rect 124000 31300 124100 31400
rect 124000 31400 124100 31500
rect 124000 31500 124100 31600
rect 124000 31600 124100 31700
rect 124000 31700 124100 31800
rect 124000 31800 124100 31900
rect 124000 31900 124100 32000
rect 124000 32000 124100 32100
rect 124000 32100 124100 32200
rect 124000 32200 124100 32300
rect 124000 32300 124100 32400
rect 124000 32400 124100 32500
rect 124000 32500 124100 32600
rect 124000 32600 124100 32700
rect 124000 32700 124100 32800
rect 124000 32800 124100 32900
rect 124000 32900 124100 33000
rect 124000 33000 124100 33100
rect 124000 33100 124100 33200
rect 124000 33200 124100 33300
rect 124000 33300 124100 33400
rect 124000 34200 124100 34300
rect 124000 34300 124100 34400
rect 124000 34400 124100 34500
rect 124000 34500 124100 34600
rect 124000 34600 124100 34700
rect 124000 34700 124100 34800
rect 124000 34800 124100 34900
rect 124000 34900 124100 35000
rect 124000 35000 124100 35100
rect 124000 35100 124100 35200
rect 124000 35200 124100 35300
rect 124000 35300 124100 35400
rect 124000 35400 124100 35500
rect 124000 35500 124100 35600
rect 124000 35600 124100 35700
rect 124000 35700 124100 35800
rect 124000 35800 124100 35900
rect 124000 35900 124100 36000
rect 124000 36000 124100 36100
rect 124000 36100 124100 36200
rect 124000 36200 124100 36300
rect 124000 36300 124100 36400
rect 124000 36400 124100 36500
rect 124000 36500 124100 36600
rect 124000 36600 124100 36700
rect 124000 36700 124100 36800
rect 124000 36800 124100 36900
rect 124000 36900 124100 37000
rect 124000 37000 124100 37100
rect 124000 37100 124100 37200
rect 124000 37200 124100 37300
rect 124000 37300 124100 37400
rect 124000 37400 124100 37500
rect 124000 37500 124100 37600
rect 124100 22800 124200 22900
rect 124100 22900 124200 23000
rect 124100 23000 124200 23100
rect 124100 23100 124200 23200
rect 124100 23200 124200 23300
rect 124100 23300 124200 23400
rect 124100 23400 124200 23500
rect 124100 23500 124200 23600
rect 124100 23600 124200 23700
rect 124100 23700 124200 23800
rect 124100 23800 124200 23900
rect 124100 23900 124200 24000
rect 124100 24000 124200 24100
rect 124100 24100 124200 24200
rect 124100 24200 124200 24300
rect 124100 24300 124200 24400
rect 124100 24400 124200 24500
rect 124100 24500 124200 24600
rect 124100 24600 124200 24700
rect 124100 24700 124200 24800
rect 124100 24800 124200 24900
rect 124100 24900 124200 25000
rect 124100 25000 124200 25100
rect 124100 25100 124200 25200
rect 124100 25200 124200 25300
rect 124100 25300 124200 25400
rect 124100 25400 124200 25500
rect 124100 27600 124200 27700
rect 124100 27700 124200 27800
rect 124100 27800 124200 27900
rect 124100 27900 124200 28000
rect 124100 28000 124200 28100
rect 124100 28100 124200 28200
rect 124100 28200 124200 28300
rect 124100 28300 124200 28400
rect 124100 28400 124200 28500
rect 124100 28500 124200 28600
rect 124100 28600 124200 28700
rect 124100 28700 124200 28800
rect 124100 28800 124200 28900
rect 124100 28900 124200 29000
rect 124100 29000 124200 29100
rect 124100 29100 124200 29200
rect 124100 29200 124200 29300
rect 124100 29300 124200 29400
rect 124100 29400 124200 29500
rect 124100 29500 124200 29600
rect 124100 29600 124200 29700
rect 124100 29700 124200 29800
rect 124100 29800 124200 29900
rect 124100 29900 124200 30000
rect 124100 30000 124200 30100
rect 124100 30100 124200 30200
rect 124100 30200 124200 30300
rect 124100 30300 124200 30400
rect 124100 30400 124200 30500
rect 124100 30500 124200 30600
rect 124100 30600 124200 30700
rect 124100 30700 124200 30800
rect 124100 30800 124200 30900
rect 124100 30900 124200 31000
rect 124100 31000 124200 31100
rect 124100 31100 124200 31200
rect 124100 31200 124200 31300
rect 124100 31300 124200 31400
rect 124100 31400 124200 31500
rect 124100 31500 124200 31600
rect 124100 31600 124200 31700
rect 124100 31700 124200 31800
rect 124100 31800 124200 31900
rect 124100 31900 124200 32000
rect 124100 32000 124200 32100
rect 124100 32100 124200 32200
rect 124100 32200 124200 32300
rect 124100 32300 124200 32400
rect 124100 32400 124200 32500
rect 124100 32500 124200 32600
rect 124100 32600 124200 32700
rect 124100 32700 124200 32800
rect 124100 32800 124200 32900
rect 124100 34500 124200 34600
rect 124100 34600 124200 34700
rect 124100 34700 124200 34800
rect 124100 34800 124200 34900
rect 124100 34900 124200 35000
rect 124100 35000 124200 35100
rect 124100 35100 124200 35200
rect 124100 35200 124200 35300
rect 124100 35300 124200 35400
rect 124100 35400 124200 35500
rect 124100 35500 124200 35600
rect 124100 35600 124200 35700
rect 124100 35700 124200 35800
rect 124100 35800 124200 35900
rect 124100 35900 124200 36000
rect 124100 36000 124200 36100
rect 124100 36100 124200 36200
rect 124100 36200 124200 36300
rect 124100 36300 124200 36400
rect 124100 36400 124200 36500
rect 124100 36500 124200 36600
rect 124100 36600 124200 36700
rect 124100 36700 124200 36800
rect 124100 36800 124200 36900
rect 124100 36900 124200 37000
rect 124100 37000 124200 37100
rect 124100 37100 124200 37200
rect 124100 37200 124200 37300
rect 124100 37300 124200 37400
rect 124100 37400 124200 37500
rect 124200 22700 124300 22800
rect 124200 22800 124300 22900
rect 124200 22900 124300 23000
rect 124200 23000 124300 23100
rect 124200 23100 124300 23200
rect 124200 23200 124300 23300
rect 124200 23300 124300 23400
rect 124200 23400 124300 23500
rect 124200 23500 124300 23600
rect 124200 23600 124300 23700
rect 124200 23700 124300 23800
rect 124200 23800 124300 23900
rect 124200 23900 124300 24000
rect 124200 24000 124300 24100
rect 124200 24100 124300 24200
rect 124200 24200 124300 24300
rect 124200 24300 124300 24400
rect 124200 24400 124300 24500
rect 124200 24500 124300 24600
rect 124200 24600 124300 24700
rect 124200 24700 124300 24800
rect 124200 24800 124300 24900
rect 124200 24900 124300 25000
rect 124200 25000 124300 25100
rect 124200 25100 124300 25200
rect 124200 25200 124300 25300
rect 124200 25300 124300 25400
rect 124200 25400 124300 25500
rect 124200 25500 124300 25600
rect 124200 25600 124300 25700
rect 124200 27300 124300 27400
rect 124200 27400 124300 27500
rect 124200 27500 124300 27600
rect 124200 27600 124300 27700
rect 124200 27700 124300 27800
rect 124200 27800 124300 27900
rect 124200 27900 124300 28000
rect 124200 28000 124300 28100
rect 124200 28100 124300 28200
rect 124200 28200 124300 28300
rect 124200 28300 124300 28400
rect 124200 28400 124300 28500
rect 124200 28500 124300 28600
rect 124200 28600 124300 28700
rect 124200 28700 124300 28800
rect 124200 28800 124300 28900
rect 124200 28900 124300 29000
rect 124200 29000 124300 29100
rect 124200 29100 124300 29200
rect 124200 29200 124300 29300
rect 124200 29300 124300 29400
rect 124200 29400 124300 29500
rect 124200 29500 124300 29600
rect 124200 29600 124300 29700
rect 124200 29700 124300 29800
rect 124200 29800 124300 29900
rect 124200 29900 124300 30000
rect 124200 30000 124300 30100
rect 124200 30100 124300 30200
rect 124200 30200 124300 30300
rect 124200 30300 124300 30400
rect 124200 30400 124300 30500
rect 124200 30500 124300 30600
rect 124200 30600 124300 30700
rect 124200 30700 124300 30800
rect 124200 30800 124300 30900
rect 124200 30900 124300 31000
rect 124200 31000 124300 31100
rect 124200 31100 124300 31200
rect 124200 31200 124300 31300
rect 124200 31300 124300 31400
rect 124200 31400 124300 31500
rect 124200 31500 124300 31600
rect 124200 31600 124300 31700
rect 124200 31700 124300 31800
rect 124200 31800 124300 31900
rect 124200 31900 124300 32000
rect 124200 32000 124300 32100
rect 124200 32100 124300 32200
rect 124200 32200 124300 32300
rect 124200 32300 124300 32400
rect 124200 32400 124300 32500
rect 124200 32500 124300 32600
rect 124200 34700 124300 34800
rect 124200 34800 124300 34900
rect 124200 34900 124300 35000
rect 124200 35000 124300 35100
rect 124200 35100 124300 35200
rect 124200 35200 124300 35300
rect 124200 35300 124300 35400
rect 124200 35400 124300 35500
rect 124200 35500 124300 35600
rect 124200 35600 124300 35700
rect 124200 35700 124300 35800
rect 124200 35800 124300 35900
rect 124200 35900 124300 36000
rect 124200 36000 124300 36100
rect 124200 36100 124300 36200
rect 124200 36200 124300 36300
rect 124200 36300 124300 36400
rect 124200 36400 124300 36500
rect 124200 36500 124300 36600
rect 124200 36600 124300 36700
rect 124200 36700 124300 36800
rect 124200 36800 124300 36900
rect 124200 36900 124300 37000
rect 124200 37000 124300 37100
rect 124200 37100 124300 37200
rect 124200 37200 124300 37300
rect 124300 22500 124400 22600
rect 124300 22600 124400 22700
rect 124300 22700 124400 22800
rect 124300 22800 124400 22900
rect 124300 22900 124400 23000
rect 124300 23000 124400 23100
rect 124300 23100 124400 23200
rect 124300 23200 124400 23300
rect 124300 23300 124400 23400
rect 124300 23400 124400 23500
rect 124300 23500 124400 23600
rect 124300 23600 124400 23700
rect 124300 23700 124400 23800
rect 124300 23800 124400 23900
rect 124300 23900 124400 24000
rect 124300 24000 124400 24100
rect 124300 24100 124400 24200
rect 124300 24200 124400 24300
rect 124300 24300 124400 24400
rect 124300 24400 124400 24500
rect 124300 24500 124400 24600
rect 124300 24600 124400 24700
rect 124300 24700 124400 24800
rect 124300 24800 124400 24900
rect 124300 24900 124400 25000
rect 124300 25000 124400 25100
rect 124300 25100 124400 25200
rect 124300 25200 124400 25300
rect 124300 25300 124400 25400
rect 124300 25400 124400 25500
rect 124300 25500 124400 25600
rect 124300 25600 124400 25700
rect 124300 25700 124400 25800
rect 124300 25800 124400 25900
rect 124300 25900 124400 26000
rect 124300 26800 124400 26900
rect 124300 26900 124400 27000
rect 124300 27000 124400 27100
rect 124300 27100 124400 27200
rect 124300 27200 124400 27300
rect 124300 27300 124400 27400
rect 124300 27400 124400 27500
rect 124300 27500 124400 27600
rect 124300 27600 124400 27700
rect 124300 27700 124400 27800
rect 124300 27800 124400 27900
rect 124300 27900 124400 28000
rect 124300 28000 124400 28100
rect 124300 28100 124400 28200
rect 124300 28200 124400 28300
rect 124300 28300 124400 28400
rect 124300 28400 124400 28500
rect 124300 28500 124400 28600
rect 124300 28600 124400 28700
rect 124300 28700 124400 28800
rect 124300 28800 124400 28900
rect 124300 28900 124400 29000
rect 124300 29000 124400 29100
rect 124300 29100 124400 29200
rect 124300 29200 124400 29300
rect 124300 29300 124400 29400
rect 124300 29400 124400 29500
rect 124300 29500 124400 29600
rect 124300 29600 124400 29700
rect 124300 29700 124400 29800
rect 124300 29800 124400 29900
rect 124300 29900 124400 30000
rect 124300 30000 124400 30100
rect 124300 30100 124400 30200
rect 124300 30200 124400 30300
rect 124300 30300 124400 30400
rect 124300 30400 124400 30500
rect 124300 30500 124400 30600
rect 124300 30600 124400 30700
rect 124300 30700 124400 30800
rect 124300 30800 124400 30900
rect 124300 30900 124400 31000
rect 124300 31000 124400 31100
rect 124300 31100 124400 31200
rect 124300 31200 124400 31300
rect 124300 31300 124400 31400
rect 124300 31400 124400 31500
rect 124300 31500 124400 31600
rect 124300 31600 124400 31700
rect 124300 31700 124400 31800
rect 124300 31800 124400 31900
rect 124300 31900 124400 32000
rect 124300 32000 124400 32100
rect 124300 32100 124400 32200
rect 124300 34900 124400 35000
rect 124300 35000 124400 35100
rect 124300 35100 124400 35200
rect 124300 35200 124400 35300
rect 124300 35300 124400 35400
rect 124300 35400 124400 35500
rect 124300 35500 124400 35600
rect 124300 35600 124400 35700
rect 124300 35700 124400 35800
rect 124300 35800 124400 35900
rect 124300 35900 124400 36000
rect 124300 36000 124400 36100
rect 124300 36100 124400 36200
rect 124300 36200 124400 36300
rect 124300 36300 124400 36400
rect 124300 36400 124400 36500
rect 124300 36500 124400 36600
rect 124300 36600 124400 36700
rect 124300 36700 124400 36800
rect 124300 36800 124400 36900
rect 124300 36900 124400 37000
rect 124300 37000 124400 37100
rect 124300 37100 124400 37200
rect 124400 22400 124500 22500
rect 124400 22500 124500 22600
rect 124400 22600 124500 22700
rect 124400 22700 124500 22800
rect 124400 22800 124500 22900
rect 124400 22900 124500 23000
rect 124400 23000 124500 23100
rect 124400 23100 124500 23200
rect 124400 23200 124500 23300
rect 124400 23300 124500 23400
rect 124400 23400 124500 23500
rect 124400 23500 124500 23600
rect 124400 23600 124500 23700
rect 124400 23700 124500 23800
rect 124400 23800 124500 23900
rect 124400 23900 124500 24000
rect 124400 24000 124500 24100
rect 124400 24100 124500 24200
rect 124400 24200 124500 24300
rect 124400 24300 124500 24400
rect 124400 24400 124500 24500
rect 124400 24500 124500 24600
rect 124400 24600 124500 24700
rect 124400 24700 124500 24800
rect 124400 24800 124500 24900
rect 124400 24900 124500 25000
rect 124400 25000 124500 25100
rect 124400 25100 124500 25200
rect 124400 25200 124500 25300
rect 124400 25300 124500 25400
rect 124400 25400 124500 25500
rect 124400 25500 124500 25600
rect 124400 25600 124500 25700
rect 124400 25700 124500 25800
rect 124400 25800 124500 25900
rect 124400 25900 124500 26000
rect 124400 26000 124500 26100
rect 124400 26100 124500 26200
rect 124400 26200 124500 26300
rect 124400 26300 124500 26400
rect 124400 26400 124500 26500
rect 124400 26500 124500 26600
rect 124400 26600 124500 26700
rect 124400 26700 124500 26800
rect 124400 26800 124500 26900
rect 124400 26900 124500 27000
rect 124400 27000 124500 27100
rect 124400 27100 124500 27200
rect 124400 27200 124500 27300
rect 124400 27300 124500 27400
rect 124400 27400 124500 27500
rect 124400 27500 124500 27600
rect 124400 27600 124500 27700
rect 124400 27700 124500 27800
rect 124400 27800 124500 27900
rect 124400 27900 124500 28000
rect 124400 28000 124500 28100
rect 124400 28100 124500 28200
rect 124400 28200 124500 28300
rect 124400 28300 124500 28400
rect 124400 28400 124500 28500
rect 124400 28500 124500 28600
rect 124400 28600 124500 28700
rect 124400 28700 124500 28800
rect 124400 28800 124500 28900
rect 124400 28900 124500 29000
rect 124400 29000 124500 29100
rect 124400 29100 124500 29200
rect 124400 29200 124500 29300
rect 124400 29300 124500 29400
rect 124400 29400 124500 29500
rect 124400 29500 124500 29600
rect 124400 29600 124500 29700
rect 124400 29700 124500 29800
rect 124400 29800 124500 29900
rect 124400 29900 124500 30000
rect 124400 30000 124500 30100
rect 124400 30100 124500 30200
rect 124400 30200 124500 30300
rect 124400 30300 124500 30400
rect 124400 30400 124500 30500
rect 124400 30500 124500 30600
rect 124400 30600 124500 30700
rect 124400 30700 124500 30800
rect 124400 30800 124500 30900
rect 124400 30900 124500 31000
rect 124400 31000 124500 31100
rect 124400 31100 124500 31200
rect 124400 31200 124500 31300
rect 124400 31300 124500 31400
rect 124400 31400 124500 31500
rect 124400 31500 124500 31600
rect 124400 31600 124500 31700
rect 124400 31700 124500 31800
rect 124400 31800 124500 31900
rect 124400 35100 124500 35200
rect 124400 35200 124500 35300
rect 124400 35300 124500 35400
rect 124400 35400 124500 35500
rect 124400 35500 124500 35600
rect 124400 35600 124500 35700
rect 124400 35700 124500 35800
rect 124400 35800 124500 35900
rect 124400 35900 124500 36000
rect 124400 36000 124500 36100
rect 124400 36100 124500 36200
rect 124400 36200 124500 36300
rect 124400 36300 124500 36400
rect 124400 36400 124500 36500
rect 124400 36500 124500 36600
rect 124400 36600 124500 36700
rect 124400 36700 124500 36800
rect 124400 36800 124500 36900
rect 124500 22300 124600 22400
rect 124500 22400 124600 22500
rect 124500 22500 124600 22600
rect 124500 22600 124600 22700
rect 124500 22700 124600 22800
rect 124500 22800 124600 22900
rect 124500 22900 124600 23000
rect 124500 23000 124600 23100
rect 124500 23100 124600 23200
rect 124500 23200 124600 23300
rect 124500 23300 124600 23400
rect 124500 23400 124600 23500
rect 124500 23500 124600 23600
rect 124500 23600 124600 23700
rect 124500 23700 124600 23800
rect 124500 23800 124600 23900
rect 124500 23900 124600 24000
rect 124500 24000 124600 24100
rect 124500 24100 124600 24200
rect 124500 24200 124600 24300
rect 124500 24300 124600 24400
rect 124500 24400 124600 24500
rect 124500 24500 124600 24600
rect 124500 24600 124600 24700
rect 124500 24700 124600 24800
rect 124500 24800 124600 24900
rect 124500 24900 124600 25000
rect 124500 25000 124600 25100
rect 124500 25100 124600 25200
rect 124500 25200 124600 25300
rect 124500 25300 124600 25400
rect 124500 25400 124600 25500
rect 124500 25500 124600 25600
rect 124500 25600 124600 25700
rect 124500 25700 124600 25800
rect 124500 25800 124600 25900
rect 124500 25900 124600 26000
rect 124500 26000 124600 26100
rect 124500 26100 124600 26200
rect 124500 26200 124600 26300
rect 124500 26300 124600 26400
rect 124500 26400 124600 26500
rect 124500 26500 124600 26600
rect 124500 26600 124600 26700
rect 124500 26700 124600 26800
rect 124500 26800 124600 26900
rect 124500 26900 124600 27000
rect 124500 27000 124600 27100
rect 124500 27100 124600 27200
rect 124500 27200 124600 27300
rect 124500 27300 124600 27400
rect 124500 27400 124600 27500
rect 124500 27500 124600 27600
rect 124500 27600 124600 27700
rect 124500 27700 124600 27800
rect 124500 27800 124600 27900
rect 124500 27900 124600 28000
rect 124500 28000 124600 28100
rect 124500 28100 124600 28200
rect 124500 28200 124600 28300
rect 124500 28300 124600 28400
rect 124500 28400 124600 28500
rect 124500 28500 124600 28600
rect 124500 28600 124600 28700
rect 124500 28700 124600 28800
rect 124500 28800 124600 28900
rect 124500 28900 124600 29000
rect 124500 29000 124600 29100
rect 124500 29100 124600 29200
rect 124500 29200 124600 29300
rect 124500 29300 124600 29400
rect 124500 29400 124600 29500
rect 124500 29500 124600 29600
rect 124500 29600 124600 29700
rect 124500 29700 124600 29800
rect 124500 29800 124600 29900
rect 124500 29900 124600 30000
rect 124500 30000 124600 30100
rect 124500 30100 124600 30200
rect 124500 30200 124600 30300
rect 124500 30300 124600 30400
rect 124500 30400 124600 30500
rect 124500 30500 124600 30600
rect 124500 30600 124600 30700
rect 124500 30700 124600 30800
rect 124500 30800 124600 30900
rect 124500 30900 124600 31000
rect 124500 31000 124600 31100
rect 124500 31100 124600 31200
rect 124500 31200 124600 31300
rect 124500 31300 124600 31400
rect 124500 31400 124600 31500
rect 124500 31500 124600 31600
rect 124500 35400 124600 35500
rect 124500 35500 124600 35600
rect 124500 35600 124600 35700
rect 124500 35700 124600 35800
rect 124500 35800 124600 35900
rect 124500 35900 124600 36000
rect 124500 36000 124600 36100
rect 124500 36100 124600 36200
rect 124500 36200 124600 36300
rect 124500 36300 124600 36400
rect 124500 36400 124600 36500
rect 124500 36500 124600 36600
rect 124600 22200 124700 22300
rect 124600 22300 124700 22400
rect 124600 22400 124700 22500
rect 124600 22500 124700 22600
rect 124600 22600 124700 22700
rect 124600 22700 124700 22800
rect 124600 22800 124700 22900
rect 124600 22900 124700 23000
rect 124600 23000 124700 23100
rect 124600 23100 124700 23200
rect 124600 23200 124700 23300
rect 124600 23300 124700 23400
rect 124600 23400 124700 23500
rect 124600 23500 124700 23600
rect 124600 23600 124700 23700
rect 124600 23700 124700 23800
rect 124600 23800 124700 23900
rect 124600 23900 124700 24000
rect 124600 24000 124700 24100
rect 124600 24100 124700 24200
rect 124600 24200 124700 24300
rect 124600 24300 124700 24400
rect 124600 24400 124700 24500
rect 124600 24500 124700 24600
rect 124600 24600 124700 24700
rect 124600 24700 124700 24800
rect 124600 24800 124700 24900
rect 124600 24900 124700 25000
rect 124600 25000 124700 25100
rect 124600 25100 124700 25200
rect 124600 25200 124700 25300
rect 124600 25300 124700 25400
rect 124600 25400 124700 25500
rect 124600 25500 124700 25600
rect 124600 25600 124700 25700
rect 124600 25700 124700 25800
rect 124600 25800 124700 25900
rect 124600 25900 124700 26000
rect 124600 26000 124700 26100
rect 124600 26100 124700 26200
rect 124600 26200 124700 26300
rect 124600 26300 124700 26400
rect 124600 26400 124700 26500
rect 124600 26500 124700 26600
rect 124600 26600 124700 26700
rect 124600 26700 124700 26800
rect 124600 26800 124700 26900
rect 124600 26900 124700 27000
rect 124600 27000 124700 27100
rect 124600 27100 124700 27200
rect 124600 27200 124700 27300
rect 124600 27300 124700 27400
rect 124600 27400 124700 27500
rect 124600 27500 124700 27600
rect 124600 27600 124700 27700
rect 124600 27700 124700 27800
rect 124600 27800 124700 27900
rect 124600 27900 124700 28000
rect 124600 28000 124700 28100
rect 124600 28100 124700 28200
rect 124600 28200 124700 28300
rect 124600 28300 124700 28400
rect 124600 28400 124700 28500
rect 124600 28500 124700 28600
rect 124600 28600 124700 28700
rect 124600 28700 124700 28800
rect 124600 28800 124700 28900
rect 124600 28900 124700 29000
rect 124600 29000 124700 29100
rect 124600 29100 124700 29200
rect 124600 29200 124700 29300
rect 124600 29300 124700 29400
rect 124600 29400 124700 29500
rect 124600 29500 124700 29600
rect 124600 29600 124700 29700
rect 124600 29700 124700 29800
rect 124600 29800 124700 29900
rect 124600 29900 124700 30000
rect 124600 30000 124700 30100
rect 124600 30100 124700 30200
rect 124600 30200 124700 30300
rect 124600 30300 124700 30400
rect 124600 30400 124700 30500
rect 124600 30500 124700 30600
rect 124600 30600 124700 30700
rect 124600 30700 124700 30800
rect 124600 30800 124700 30900
rect 124600 30900 124700 31000
rect 124600 31000 124700 31100
rect 124600 31100 124700 31200
rect 124600 31200 124700 31300
rect 124700 22100 124800 22200
rect 124700 22200 124800 22300
rect 124700 22300 124800 22400
rect 124700 22400 124800 22500
rect 124700 22500 124800 22600
rect 124700 22600 124800 22700
rect 124700 22700 124800 22800
rect 124700 22800 124800 22900
rect 124700 22900 124800 23000
rect 124700 23000 124800 23100
rect 124700 23100 124800 23200
rect 124700 23200 124800 23300
rect 124700 23300 124800 23400
rect 124700 23400 124800 23500
rect 124700 23500 124800 23600
rect 124700 23600 124800 23700
rect 124700 23700 124800 23800
rect 124700 23800 124800 23900
rect 124700 23900 124800 24000
rect 124700 24000 124800 24100
rect 124700 24100 124800 24200
rect 124700 24200 124800 24300
rect 124700 24300 124800 24400
rect 124700 24400 124800 24500
rect 124700 24500 124800 24600
rect 124700 24600 124800 24700
rect 124700 24700 124800 24800
rect 124700 24800 124800 24900
rect 124700 24900 124800 25000
rect 124700 25000 124800 25100
rect 124700 25100 124800 25200
rect 124700 25200 124800 25300
rect 124700 25300 124800 25400
rect 124700 25400 124800 25500
rect 124700 25500 124800 25600
rect 124700 25600 124800 25700
rect 124700 25700 124800 25800
rect 124700 25800 124800 25900
rect 124700 25900 124800 26000
rect 124700 26000 124800 26100
rect 124700 26100 124800 26200
rect 124700 26200 124800 26300
rect 124700 26300 124800 26400
rect 124700 26400 124800 26500
rect 124700 26500 124800 26600
rect 124700 26600 124800 26700
rect 124700 26700 124800 26800
rect 124700 26800 124800 26900
rect 124700 26900 124800 27000
rect 124700 27000 124800 27100
rect 124700 27100 124800 27200
rect 124700 27200 124800 27300
rect 124700 27300 124800 27400
rect 124700 27400 124800 27500
rect 124700 27500 124800 27600
rect 124700 27600 124800 27700
rect 124700 27700 124800 27800
rect 124700 27800 124800 27900
rect 124700 27900 124800 28000
rect 124700 28000 124800 28100
rect 124700 28100 124800 28200
rect 124700 28200 124800 28300
rect 124700 28300 124800 28400
rect 124700 28400 124800 28500
rect 124700 28500 124800 28600
rect 124700 28600 124800 28700
rect 124700 28700 124800 28800
rect 124700 28800 124800 28900
rect 124700 28900 124800 29000
rect 124700 29000 124800 29100
rect 124700 29100 124800 29200
rect 124700 29200 124800 29300
rect 124700 29300 124800 29400
rect 124700 29400 124800 29500
rect 124700 29500 124800 29600
rect 124700 29600 124800 29700
rect 124700 29700 124800 29800
rect 124700 29800 124800 29900
rect 124700 29900 124800 30000
rect 124700 30000 124800 30100
rect 124700 30100 124800 30200
rect 124700 30200 124800 30300
rect 124700 30300 124800 30400
rect 124700 30400 124800 30500
rect 124700 30500 124800 30600
rect 124700 30600 124800 30700
rect 124700 30700 124800 30800
rect 124700 30800 124800 30900
rect 124700 30900 124800 31000
rect 124800 22000 124900 22100
rect 124800 22100 124900 22200
rect 124800 22200 124900 22300
rect 124800 22300 124900 22400
rect 124800 22400 124900 22500
rect 124800 22500 124900 22600
rect 124800 22600 124900 22700
rect 124800 22700 124900 22800
rect 124800 22800 124900 22900
rect 124800 22900 124900 23000
rect 124800 23000 124900 23100
rect 124800 23100 124900 23200
rect 124800 23200 124900 23300
rect 124800 23300 124900 23400
rect 124800 23400 124900 23500
rect 124800 23500 124900 23600
rect 124800 23600 124900 23700
rect 124800 23700 124900 23800
rect 124800 23800 124900 23900
rect 124800 23900 124900 24000
rect 124800 24000 124900 24100
rect 124800 24100 124900 24200
rect 124800 24200 124900 24300
rect 124800 24300 124900 24400
rect 124800 24400 124900 24500
rect 124800 24500 124900 24600
rect 124800 24600 124900 24700
rect 124800 24700 124900 24800
rect 124800 24800 124900 24900
rect 124800 24900 124900 25000
rect 124800 25000 124900 25100
rect 124800 25100 124900 25200
rect 124800 25200 124900 25300
rect 124800 25300 124900 25400
rect 124800 25400 124900 25500
rect 124800 25500 124900 25600
rect 124800 25600 124900 25700
rect 124800 25700 124900 25800
rect 124800 25800 124900 25900
rect 124800 25900 124900 26000
rect 124800 26000 124900 26100
rect 124800 26100 124900 26200
rect 124800 26200 124900 26300
rect 124800 26300 124900 26400
rect 124800 26400 124900 26500
rect 124800 26500 124900 26600
rect 124800 26600 124900 26700
rect 124800 26700 124900 26800
rect 124800 26800 124900 26900
rect 124800 26900 124900 27000
rect 124800 27000 124900 27100
rect 124800 27100 124900 27200
rect 124800 27200 124900 27300
rect 124800 27300 124900 27400
rect 124800 27400 124900 27500
rect 124800 27500 124900 27600
rect 124800 27600 124900 27700
rect 124800 27700 124900 27800
rect 124800 27800 124900 27900
rect 124800 27900 124900 28000
rect 124800 28000 124900 28100
rect 124800 28100 124900 28200
rect 124800 28200 124900 28300
rect 124800 28300 124900 28400
rect 124800 28400 124900 28500
rect 124800 28500 124900 28600
rect 124800 28600 124900 28700
rect 124800 28700 124900 28800
rect 124800 28800 124900 28900
rect 124800 28900 124900 29000
rect 124800 29000 124900 29100
rect 124800 29100 124900 29200
rect 124800 29200 124900 29300
rect 124800 29300 124900 29400
rect 124800 29400 124900 29500
rect 124800 29500 124900 29600
rect 124800 29600 124900 29700
rect 124800 29700 124900 29800
rect 124800 29800 124900 29900
rect 124800 29900 124900 30000
rect 124800 30000 124900 30100
rect 124800 30100 124900 30200
rect 124800 30200 124900 30300
rect 124800 30300 124900 30400
rect 124800 30400 124900 30500
rect 124800 30500 124900 30600
rect 124800 30600 124900 30700
rect 124900 22000 125000 22100
rect 124900 22100 125000 22200
rect 124900 22200 125000 22300
rect 124900 22300 125000 22400
rect 124900 22400 125000 22500
rect 124900 22500 125000 22600
rect 124900 22600 125000 22700
rect 124900 22700 125000 22800
rect 124900 22800 125000 22900
rect 124900 22900 125000 23000
rect 124900 23000 125000 23100
rect 124900 23100 125000 23200
rect 124900 23200 125000 23300
rect 124900 23300 125000 23400
rect 124900 23400 125000 23500
rect 124900 23500 125000 23600
rect 124900 23600 125000 23700
rect 124900 23700 125000 23800
rect 124900 23800 125000 23900
rect 124900 23900 125000 24000
rect 124900 24000 125000 24100
rect 124900 24100 125000 24200
rect 124900 24200 125000 24300
rect 124900 24300 125000 24400
rect 124900 24400 125000 24500
rect 124900 24500 125000 24600
rect 124900 24600 125000 24700
rect 124900 24700 125000 24800
rect 124900 24800 125000 24900
rect 124900 24900 125000 25000
rect 124900 25000 125000 25100
rect 124900 25100 125000 25200
rect 124900 25200 125000 25300
rect 124900 25300 125000 25400
rect 124900 25400 125000 25500
rect 124900 25500 125000 25600
rect 124900 25600 125000 25700
rect 124900 25700 125000 25800
rect 124900 25800 125000 25900
rect 124900 25900 125000 26000
rect 124900 26000 125000 26100
rect 124900 26100 125000 26200
rect 124900 26200 125000 26300
rect 124900 26300 125000 26400
rect 124900 26400 125000 26500
rect 124900 26500 125000 26600
rect 124900 26600 125000 26700
rect 124900 26700 125000 26800
rect 124900 26800 125000 26900
rect 124900 26900 125000 27000
rect 124900 27000 125000 27100
rect 124900 27100 125000 27200
rect 124900 27200 125000 27300
rect 124900 27300 125000 27400
rect 124900 27400 125000 27500
rect 124900 27500 125000 27600
rect 124900 27600 125000 27700
rect 124900 27700 125000 27800
rect 124900 27800 125000 27900
rect 124900 27900 125000 28000
rect 124900 28000 125000 28100
rect 124900 28100 125000 28200
rect 124900 28200 125000 28300
rect 124900 28300 125000 28400
rect 124900 28400 125000 28500
rect 124900 28500 125000 28600
rect 124900 28600 125000 28700
rect 124900 28700 125000 28800
rect 124900 28800 125000 28900
rect 124900 28900 125000 29000
rect 124900 29000 125000 29100
rect 124900 29100 125000 29200
rect 124900 29200 125000 29300
rect 124900 29300 125000 29400
rect 124900 29400 125000 29500
rect 124900 29500 125000 29600
rect 124900 29600 125000 29700
rect 124900 29700 125000 29800
rect 124900 29800 125000 29900
rect 124900 29900 125000 30000
rect 124900 30000 125000 30100
rect 124900 30100 125000 30200
rect 124900 30200 125000 30300
rect 124900 30300 125000 30400
rect 125000 21900 125100 22000
rect 125000 22000 125100 22100
rect 125000 22100 125100 22200
rect 125000 22200 125100 22300
rect 125000 22300 125100 22400
rect 125000 22400 125100 22500
rect 125000 22500 125100 22600
rect 125000 22600 125100 22700
rect 125000 22700 125100 22800
rect 125000 22800 125100 22900
rect 125000 22900 125100 23000
rect 125000 23000 125100 23100
rect 125000 23100 125100 23200
rect 125000 23200 125100 23300
rect 125000 23300 125100 23400
rect 125000 23400 125100 23500
rect 125000 23500 125100 23600
rect 125000 23600 125100 23700
rect 125000 23700 125100 23800
rect 125000 23800 125100 23900
rect 125000 23900 125100 24000
rect 125000 24000 125100 24100
rect 125000 24100 125100 24200
rect 125000 24200 125100 24300
rect 125000 24300 125100 24400
rect 125000 24400 125100 24500
rect 125000 24500 125100 24600
rect 125000 24600 125100 24700
rect 125000 24700 125100 24800
rect 125000 24800 125100 24900
rect 125000 24900 125100 25000
rect 125000 25000 125100 25100
rect 125000 25100 125100 25200
rect 125000 25200 125100 25300
rect 125000 25300 125100 25400
rect 125000 25400 125100 25500
rect 125000 25500 125100 25600
rect 125000 25600 125100 25700
rect 125000 25700 125100 25800
rect 125000 25800 125100 25900
rect 125000 25900 125100 26000
rect 125000 26000 125100 26100
rect 125000 26100 125100 26200
rect 125000 26200 125100 26300
rect 125000 26300 125100 26400
rect 125000 26400 125100 26500
rect 125000 26500 125100 26600
rect 125000 26600 125100 26700
rect 125000 26700 125100 26800
rect 125000 26800 125100 26900
rect 125000 26900 125100 27000
rect 125000 27000 125100 27100
rect 125000 27100 125100 27200
rect 125000 27200 125100 27300
rect 125000 27300 125100 27400
rect 125000 27400 125100 27500
rect 125000 27500 125100 27600
rect 125000 27600 125100 27700
rect 125000 27700 125100 27800
rect 125000 27800 125100 27900
rect 125000 27900 125100 28000
rect 125000 28000 125100 28100
rect 125000 28100 125100 28200
rect 125000 28200 125100 28300
rect 125000 28300 125100 28400
rect 125000 28400 125100 28500
rect 125000 28500 125100 28600
rect 125000 28600 125100 28700
rect 125000 28700 125100 28800
rect 125000 28800 125100 28900
rect 125000 28900 125100 29000
rect 125000 29000 125100 29100
rect 125000 29100 125100 29200
rect 125000 29200 125100 29300
rect 125000 29300 125100 29400
rect 125000 29400 125100 29500
rect 125000 29500 125100 29600
rect 125000 29600 125100 29700
rect 125000 29700 125100 29800
rect 125000 29800 125100 29900
rect 125000 29900 125100 30000
rect 125000 30000 125100 30100
rect 125100 21900 125200 22000
rect 125100 22000 125200 22100
rect 125100 22100 125200 22200
rect 125100 22200 125200 22300
rect 125100 22300 125200 22400
rect 125100 22400 125200 22500
rect 125100 22500 125200 22600
rect 125100 22600 125200 22700
rect 125100 22700 125200 22800
rect 125100 22800 125200 22900
rect 125100 22900 125200 23000
rect 125100 23000 125200 23100
rect 125100 23100 125200 23200
rect 125100 23200 125200 23300
rect 125100 23300 125200 23400
rect 125100 23400 125200 23500
rect 125100 23500 125200 23600
rect 125100 23600 125200 23700
rect 125100 23700 125200 23800
rect 125100 23800 125200 23900
rect 125100 23900 125200 24000
rect 125100 24000 125200 24100
rect 125100 24100 125200 24200
rect 125100 24200 125200 24300
rect 125100 24300 125200 24400
rect 125100 24400 125200 24500
rect 125100 24500 125200 24600
rect 125100 24600 125200 24700
rect 125100 24700 125200 24800
rect 125100 24800 125200 24900
rect 125100 24900 125200 25000
rect 125100 25000 125200 25100
rect 125100 25100 125200 25200
rect 125100 25200 125200 25300
rect 125100 25300 125200 25400
rect 125100 25400 125200 25500
rect 125100 25500 125200 25600
rect 125100 25600 125200 25700
rect 125100 25700 125200 25800
rect 125100 25800 125200 25900
rect 125100 25900 125200 26000
rect 125100 26000 125200 26100
rect 125100 26100 125200 26200
rect 125100 26200 125200 26300
rect 125100 26300 125200 26400
rect 125100 26400 125200 26500
rect 125100 26500 125200 26600
rect 125100 26600 125200 26700
rect 125100 26700 125200 26800
rect 125100 26800 125200 26900
rect 125100 26900 125200 27000
rect 125100 27000 125200 27100
rect 125100 27100 125200 27200
rect 125100 27200 125200 27300
rect 125100 27300 125200 27400
rect 125100 27400 125200 27500
rect 125100 27500 125200 27600
rect 125100 27600 125200 27700
rect 125100 27700 125200 27800
rect 125100 27800 125200 27900
rect 125100 27900 125200 28000
rect 125100 28000 125200 28100
rect 125100 28100 125200 28200
rect 125100 28200 125200 28300
rect 125100 28300 125200 28400
rect 125100 28400 125200 28500
rect 125100 28500 125200 28600
rect 125100 28600 125200 28700
rect 125100 28700 125200 28800
rect 125100 28800 125200 28900
rect 125100 28900 125200 29000
rect 125100 29000 125200 29100
rect 125100 29100 125200 29200
rect 125100 29200 125200 29300
rect 125100 29300 125200 29400
rect 125100 29400 125200 29500
rect 125100 29500 125200 29600
rect 125100 29600 125200 29700
rect 125100 29700 125200 29800
rect 125200 21900 125300 22000
rect 125200 22000 125300 22100
rect 125200 22100 125300 22200
rect 125200 22200 125300 22300
rect 125200 22300 125300 22400
rect 125200 22400 125300 22500
rect 125200 22500 125300 22600
rect 125200 22600 125300 22700
rect 125200 22700 125300 22800
rect 125200 22800 125300 22900
rect 125200 22900 125300 23000
rect 125200 23000 125300 23100
rect 125200 23100 125300 23200
rect 125200 23200 125300 23300
rect 125200 23300 125300 23400
rect 125200 23400 125300 23500
rect 125200 23500 125300 23600
rect 125200 23600 125300 23700
rect 125200 23700 125300 23800
rect 125200 23800 125300 23900
rect 125200 23900 125300 24000
rect 125200 24000 125300 24100
rect 125200 24100 125300 24200
rect 125200 24200 125300 24300
rect 125200 24300 125300 24400
rect 125200 24400 125300 24500
rect 125200 24500 125300 24600
rect 125200 24600 125300 24700
rect 125200 24700 125300 24800
rect 125200 24800 125300 24900
rect 125200 24900 125300 25000
rect 125200 25000 125300 25100
rect 125200 25100 125300 25200
rect 125200 25200 125300 25300
rect 125200 25300 125300 25400
rect 125200 25400 125300 25500
rect 125200 25500 125300 25600
rect 125200 25600 125300 25700
rect 125200 25700 125300 25800
rect 125200 25800 125300 25900
rect 125200 25900 125300 26000
rect 125200 26000 125300 26100
rect 125200 26100 125300 26200
rect 125200 26200 125300 26300
rect 125200 26300 125300 26400
rect 125200 26400 125300 26500
rect 125200 26500 125300 26600
rect 125200 26600 125300 26700
rect 125200 26700 125300 26800
rect 125200 26800 125300 26900
rect 125200 26900 125300 27000
rect 125200 27000 125300 27100
rect 125200 27100 125300 27200
rect 125200 27200 125300 27300
rect 125200 27300 125300 27400
rect 125200 27400 125300 27500
rect 125200 27500 125300 27600
rect 125200 27600 125300 27700
rect 125200 27700 125300 27800
rect 125200 27800 125300 27900
rect 125200 27900 125300 28000
rect 125200 28000 125300 28100
rect 125200 28100 125300 28200
rect 125200 28200 125300 28300
rect 125200 28300 125300 28400
rect 125200 28400 125300 28500
rect 125200 28500 125300 28600
rect 125200 28600 125300 28700
rect 125200 28700 125300 28800
rect 125200 28800 125300 28900
rect 125200 28900 125300 29000
rect 125200 29000 125300 29100
rect 125200 29100 125300 29200
rect 125200 29200 125300 29300
rect 125200 29300 125300 29400
rect 125200 29400 125300 29500
rect 125200 29500 125300 29600
rect 125300 21800 125400 21900
rect 125300 21900 125400 22000
rect 125300 22000 125400 22100
rect 125300 22100 125400 22200
rect 125300 22200 125400 22300
rect 125300 22300 125400 22400
rect 125300 22400 125400 22500
rect 125300 22500 125400 22600
rect 125300 22600 125400 22700
rect 125300 22700 125400 22800
rect 125300 22800 125400 22900
rect 125300 22900 125400 23000
rect 125300 23000 125400 23100
rect 125300 23100 125400 23200
rect 125300 23200 125400 23300
rect 125300 23300 125400 23400
rect 125300 23400 125400 23500
rect 125300 23500 125400 23600
rect 125300 23600 125400 23700
rect 125300 23700 125400 23800
rect 125300 23800 125400 23900
rect 125300 23900 125400 24000
rect 125300 24000 125400 24100
rect 125300 24100 125400 24200
rect 125300 24200 125400 24300
rect 125300 24300 125400 24400
rect 125300 24400 125400 24500
rect 125300 24500 125400 24600
rect 125300 24600 125400 24700
rect 125300 24700 125400 24800
rect 125300 24800 125400 24900
rect 125300 24900 125400 25000
rect 125300 25000 125400 25100
rect 125300 25100 125400 25200
rect 125300 25200 125400 25300
rect 125300 25300 125400 25400
rect 125300 25400 125400 25500
rect 125300 25500 125400 25600
rect 125300 25600 125400 25700
rect 125300 25700 125400 25800
rect 125300 25800 125400 25900
rect 125300 25900 125400 26000
rect 125300 26000 125400 26100
rect 125300 26100 125400 26200
rect 125300 26200 125400 26300
rect 125300 26300 125400 26400
rect 125300 26400 125400 26500
rect 125300 26500 125400 26600
rect 125300 26600 125400 26700
rect 125300 26700 125400 26800
rect 125300 26800 125400 26900
rect 125300 26900 125400 27000
rect 125300 27000 125400 27100
rect 125300 27100 125400 27200
rect 125300 27200 125400 27300
rect 125300 27300 125400 27400
rect 125300 27400 125400 27500
rect 125300 27500 125400 27600
rect 125300 27600 125400 27700
rect 125300 27700 125400 27800
rect 125300 27800 125400 27900
rect 125300 27900 125400 28000
rect 125300 28000 125400 28100
rect 125300 28100 125400 28200
rect 125300 28200 125400 28300
rect 125300 28300 125400 28400
rect 125300 28400 125400 28500
rect 125300 28500 125400 28600
rect 125300 28600 125400 28700
rect 125300 28700 125400 28800
rect 125300 28800 125400 28900
rect 125300 28900 125400 29000
rect 125300 29000 125400 29100
rect 125300 29100 125400 29200
rect 125300 29200 125400 29300
rect 125400 21800 125500 21900
rect 125400 21900 125500 22000
rect 125400 22000 125500 22100
rect 125400 22100 125500 22200
rect 125400 22200 125500 22300
rect 125400 22300 125500 22400
rect 125400 22400 125500 22500
rect 125400 22500 125500 22600
rect 125400 22600 125500 22700
rect 125400 22700 125500 22800
rect 125400 22800 125500 22900
rect 125400 22900 125500 23000
rect 125400 23000 125500 23100
rect 125400 23100 125500 23200
rect 125400 23200 125500 23300
rect 125400 23300 125500 23400
rect 125400 23400 125500 23500
rect 125400 23500 125500 23600
rect 125400 23600 125500 23700
rect 125400 23700 125500 23800
rect 125400 23800 125500 23900
rect 125400 23900 125500 24000
rect 125400 24300 125500 24400
rect 125400 24400 125500 24500
rect 125400 24500 125500 24600
rect 125400 24600 125500 24700
rect 125400 24700 125500 24800
rect 125400 24800 125500 24900
rect 125400 24900 125500 25000
rect 125400 25000 125500 25100
rect 125400 25100 125500 25200
rect 125400 25200 125500 25300
rect 125400 25300 125500 25400
rect 125400 25400 125500 25500
rect 125400 25500 125500 25600
rect 125400 25600 125500 25700
rect 125400 25700 125500 25800
rect 125400 25800 125500 25900
rect 125400 25900 125500 26000
rect 125400 26000 125500 26100
rect 125400 26100 125500 26200
rect 125400 26200 125500 26300
rect 125400 26300 125500 26400
rect 125400 26400 125500 26500
rect 125400 26500 125500 26600
rect 125400 26600 125500 26700
rect 125400 26700 125500 26800
rect 125400 26800 125500 26900
rect 125400 26900 125500 27000
rect 125400 27000 125500 27100
rect 125400 27100 125500 27200
rect 125400 27200 125500 27300
rect 125400 27300 125500 27400
rect 125400 27400 125500 27500
rect 125400 27500 125500 27600
rect 125400 27600 125500 27700
rect 125400 27700 125500 27800
rect 125400 27800 125500 27900
rect 125400 27900 125500 28000
rect 125400 28000 125500 28100
rect 125400 28100 125500 28200
rect 125400 28200 125500 28300
rect 125400 28300 125500 28400
rect 125400 28400 125500 28500
rect 125400 28500 125500 28600
rect 125400 28600 125500 28700
rect 125400 28700 125500 28800
rect 125400 28800 125500 28900
rect 125400 28900 125500 29000
rect 125500 21800 125600 21900
rect 125500 21900 125600 22000
rect 125500 22000 125600 22100
rect 125500 22100 125600 22200
rect 125500 22200 125600 22300
rect 125500 22300 125600 22400
rect 125500 22400 125600 22500
rect 125500 22500 125600 22600
rect 125500 22600 125600 22700
rect 125500 22700 125600 22800
rect 125500 22800 125600 22900
rect 125500 22900 125600 23000
rect 125500 23000 125600 23100
rect 125500 23100 125600 23200
rect 125500 23200 125600 23300
rect 125500 23300 125600 23400
rect 125500 23400 125600 23500
rect 125500 23500 125600 23600
rect 125500 23600 125600 23700
rect 125500 24600 125600 24700
rect 125500 24700 125600 24800
rect 125500 24800 125600 24900
rect 125500 24900 125600 25000
rect 125500 25000 125600 25100
rect 125500 25100 125600 25200
rect 125500 25200 125600 25300
rect 125500 25300 125600 25400
rect 125500 25400 125600 25500
rect 125500 25500 125600 25600
rect 125500 25600 125600 25700
rect 125500 25700 125600 25800
rect 125500 25800 125600 25900
rect 125500 25900 125600 26000
rect 125500 26000 125600 26100
rect 125500 26100 125600 26200
rect 125500 26200 125600 26300
rect 125500 26300 125600 26400
rect 125500 26400 125600 26500
rect 125500 26500 125600 26600
rect 125500 26600 125600 26700
rect 125500 26700 125600 26800
rect 125500 26800 125600 26900
rect 125500 26900 125600 27000
rect 125500 27000 125600 27100
rect 125500 27100 125600 27200
rect 125500 27200 125600 27300
rect 125500 27300 125600 27400
rect 125500 27400 125600 27500
rect 125500 27500 125600 27600
rect 125500 27600 125600 27700
rect 125500 27700 125600 27800
rect 125500 27800 125600 27900
rect 125500 27900 125600 28000
rect 125500 28000 125600 28100
rect 125500 28100 125600 28200
rect 125500 28200 125600 28300
rect 125500 28300 125600 28400
rect 125500 28400 125600 28500
rect 125500 28500 125600 28600
rect 125500 28600 125600 28700
rect 125600 21800 125700 21900
rect 125600 21900 125700 22000
rect 125600 22000 125700 22100
rect 125600 22100 125700 22200
rect 125600 22200 125700 22300
rect 125600 22300 125700 22400
rect 125600 22400 125700 22500
rect 125600 22500 125700 22600
rect 125600 22600 125700 22700
rect 125600 22700 125700 22800
rect 125600 22800 125700 22900
rect 125600 22900 125700 23000
rect 125600 23000 125700 23100
rect 125600 23100 125700 23200
rect 125600 23200 125700 23300
rect 125600 23300 125700 23400
rect 125600 23400 125700 23500
rect 125600 23500 125700 23600
rect 125600 24800 125700 24900
rect 125600 24900 125700 25000
rect 125600 25000 125700 25100
rect 125600 25100 125700 25200
rect 125600 25200 125700 25300
rect 125600 25300 125700 25400
rect 125600 25400 125700 25500
rect 125600 25500 125700 25600
rect 125600 25600 125700 25700
rect 125600 25700 125700 25800
rect 125600 25800 125700 25900
rect 125600 25900 125700 26000
rect 125600 26000 125700 26100
rect 125600 26100 125700 26200
rect 125600 26200 125700 26300
rect 125600 26300 125700 26400
rect 125600 26400 125700 26500
rect 125600 26500 125700 26600
rect 125600 26600 125700 26700
rect 125600 26700 125700 26800
rect 125600 26800 125700 26900
rect 125600 26900 125700 27000
rect 125600 27000 125700 27100
rect 125600 27100 125700 27200
rect 125600 27200 125700 27300
rect 125600 27300 125700 27400
rect 125600 27400 125700 27500
rect 125600 27500 125700 27600
rect 125600 27600 125700 27700
rect 125600 27700 125700 27800
rect 125600 27800 125700 27900
rect 125600 27900 125700 28000
rect 125600 28000 125700 28100
rect 125600 28100 125700 28200
rect 125600 28200 125700 28300
rect 125600 28300 125700 28400
rect 125600 28400 125700 28500
rect 125700 21700 125800 21800
rect 125700 21800 125800 21900
rect 125700 21900 125800 22000
rect 125700 22000 125800 22100
rect 125700 22100 125800 22200
rect 125700 22200 125800 22300
rect 125700 22300 125800 22400
rect 125700 22400 125800 22500
rect 125700 22500 125800 22600
rect 125700 22600 125800 22700
rect 125700 22700 125800 22800
rect 125700 22800 125800 22900
rect 125700 22900 125800 23000
rect 125700 23000 125800 23100
rect 125700 23100 125800 23200
rect 125700 23200 125800 23300
rect 125700 23300 125800 23400
rect 125700 23400 125800 23500
rect 125700 24900 125800 25000
rect 125700 25000 125800 25100
rect 125700 25100 125800 25200
rect 125700 25200 125800 25300
rect 125700 25300 125800 25400
rect 125700 25400 125800 25500
rect 125700 25500 125800 25600
rect 125700 25600 125800 25700
rect 125700 25700 125800 25800
rect 125700 25800 125800 25900
rect 125700 25900 125800 26000
rect 125700 26000 125800 26100
rect 125700 26100 125800 26200
rect 125700 26200 125800 26300
rect 125700 26300 125800 26400
rect 125700 26400 125800 26500
rect 125700 26500 125800 26600
rect 125700 26600 125800 26700
rect 125700 26700 125800 26800
rect 125700 26800 125800 26900
rect 125700 26900 125800 27000
rect 125700 27000 125800 27100
rect 125700 27100 125800 27200
rect 125700 27200 125800 27300
rect 125700 27300 125800 27400
rect 125700 27400 125800 27500
rect 125700 27500 125800 27600
rect 125700 27600 125800 27700
rect 125700 27700 125800 27800
rect 125700 27800 125800 27900
rect 125700 27900 125800 28000
rect 125700 28000 125800 28100
rect 125700 28100 125800 28200
rect 125800 21700 125900 21800
rect 125800 21800 125900 21900
rect 125800 21900 125900 22000
rect 125800 22000 125900 22100
rect 125800 22100 125900 22200
rect 125800 22200 125900 22300
rect 125800 22300 125900 22400
rect 125800 22400 125900 22500
rect 125800 22500 125900 22600
rect 125800 22600 125900 22700
rect 125800 22700 125900 22800
rect 125800 22800 125900 22900
rect 125800 22900 125900 23000
rect 125800 23000 125900 23100
rect 125800 23100 125900 23200
rect 125800 23200 125900 23300
rect 125800 23300 125900 23400
rect 125800 24900 125900 25000
rect 125800 25000 125900 25100
rect 125800 25100 125900 25200
rect 125800 25200 125900 25300
rect 125800 25300 125900 25400
rect 125800 25400 125900 25500
rect 125800 25500 125900 25600
rect 125800 25600 125900 25700
rect 125800 25700 125900 25800
rect 125800 25800 125900 25900
rect 125800 25900 125900 26000
rect 125800 26000 125900 26100
rect 125800 26100 125900 26200
rect 125800 26200 125900 26300
rect 125800 26300 125900 26400
rect 125800 26400 125900 26500
rect 125800 26500 125900 26600
rect 125800 26600 125900 26700
rect 125800 26700 125900 26800
rect 125800 26800 125900 26900
rect 125800 26900 125900 27000
rect 125800 27000 125900 27100
rect 125800 27100 125900 27200
rect 125800 27200 125900 27300
rect 125800 27300 125900 27400
rect 125800 27400 125900 27500
rect 125800 27500 125900 27600
rect 125800 27600 125900 27700
rect 125800 27700 125900 27800
rect 125800 27800 125900 27900
rect 125800 27900 125900 28000
rect 125900 21700 126000 21800
rect 125900 21800 126000 21900
rect 125900 21900 126000 22000
rect 125900 22000 126000 22100
rect 125900 22100 126000 22200
rect 125900 22200 126000 22300
rect 125900 22300 126000 22400
rect 125900 22400 126000 22500
rect 125900 22500 126000 22600
rect 125900 22600 126000 22700
rect 125900 22700 126000 22800
rect 125900 22800 126000 22900
rect 125900 22900 126000 23000
rect 125900 23000 126000 23100
rect 125900 23100 126000 23200
rect 125900 23200 126000 23300
rect 125900 23300 126000 23400
rect 125900 24900 126000 25000
rect 125900 25000 126000 25100
rect 125900 25100 126000 25200
rect 125900 25200 126000 25300
rect 125900 25300 126000 25400
rect 125900 25400 126000 25500
rect 125900 25500 126000 25600
rect 125900 25600 126000 25700
rect 125900 25700 126000 25800
rect 125900 25800 126000 25900
rect 125900 25900 126000 26000
rect 125900 26000 126000 26100
rect 125900 26100 126000 26200
rect 125900 26200 126000 26300
rect 125900 26300 126000 26400
rect 125900 26400 126000 26500
rect 125900 26500 126000 26600
rect 125900 26600 126000 26700
rect 125900 26700 126000 26800
rect 125900 26800 126000 26900
rect 125900 26900 126000 27000
rect 125900 27000 126000 27100
rect 125900 27100 126000 27200
rect 125900 27200 126000 27300
rect 125900 27300 126000 27400
rect 125900 27400 126000 27500
rect 125900 27500 126000 27600
rect 125900 27600 126000 27700
rect 126000 21700 126100 21800
rect 126000 21800 126100 21900
rect 126000 21900 126100 22000
rect 126000 22000 126100 22100
rect 126000 22100 126100 22200
rect 126000 22200 126100 22300
rect 126000 22300 126100 22400
rect 126000 22400 126100 22500
rect 126000 22500 126100 22600
rect 126000 22600 126100 22700
rect 126000 22700 126100 22800
rect 126000 22800 126100 22900
rect 126000 22900 126100 23000
rect 126000 23000 126100 23100
rect 126000 23100 126100 23200
rect 126000 23200 126100 23300
rect 126000 23300 126100 23400
rect 126000 24900 126100 25000
rect 126000 25000 126100 25100
rect 126000 25100 126100 25200
rect 126000 25200 126100 25300
rect 126000 25300 126100 25400
rect 126000 25400 126100 25500
rect 126000 25500 126100 25600
rect 126000 25600 126100 25700
rect 126000 25700 126100 25800
rect 126000 25800 126100 25900
rect 126000 25900 126100 26000
rect 126000 26000 126100 26100
rect 126000 26100 126100 26200
rect 126000 26200 126100 26300
rect 126000 26300 126100 26400
rect 126000 26400 126100 26500
rect 126000 26500 126100 26600
rect 126000 26600 126100 26700
rect 126000 26700 126100 26800
rect 126000 26800 126100 26900
rect 126000 26900 126100 27000
rect 126000 27000 126100 27100
rect 126000 27100 126100 27200
rect 126000 27200 126100 27300
rect 126000 27300 126100 27400
rect 126000 27400 126100 27500
rect 126100 21700 126200 21800
rect 126100 21800 126200 21900
rect 126100 21900 126200 22000
rect 126100 22000 126200 22100
rect 126100 22100 126200 22200
rect 126100 22200 126200 22300
rect 126100 22300 126200 22400
rect 126100 22400 126200 22500
rect 126100 22500 126200 22600
rect 126100 22600 126200 22700
rect 126100 22700 126200 22800
rect 126100 22800 126200 22900
rect 126100 22900 126200 23000
rect 126100 23000 126200 23100
rect 126100 23100 126200 23200
rect 126100 23200 126200 23300
rect 126100 24900 126200 25000
rect 126100 25000 126200 25100
rect 126100 25100 126200 25200
rect 126100 25200 126200 25300
rect 126100 25300 126200 25400
rect 126100 25400 126200 25500
rect 126100 25500 126200 25600
rect 126100 25600 126200 25700
rect 126100 25700 126200 25800
rect 126100 25800 126200 25900
rect 126100 25900 126200 26000
rect 126100 26000 126200 26100
rect 126100 26100 126200 26200
rect 126100 26200 126200 26300
rect 126100 26300 126200 26400
rect 126100 26400 126200 26500
rect 126100 26500 126200 26600
rect 126100 26600 126200 26700
rect 126100 26700 126200 26800
rect 126100 26800 126200 26900
rect 126100 26900 126200 27000
rect 126100 27000 126200 27100
rect 126100 27100 126200 27200
rect 126100 27200 126200 27300
rect 126200 21700 126300 21800
rect 126200 21800 126300 21900
rect 126200 21900 126300 22000
rect 126200 22000 126300 22100
rect 126200 22100 126300 22200
rect 126200 22200 126300 22300
rect 126200 22300 126300 22400
rect 126200 22400 126300 22500
rect 126200 22500 126300 22600
rect 126200 22600 126300 22700
rect 126200 22700 126300 22800
rect 126200 22800 126300 22900
rect 126200 22900 126300 23000
rect 126200 23000 126300 23100
rect 126200 23100 126300 23200
rect 126200 23200 126300 23300
rect 126200 23300 126300 23400
rect 126200 24900 126300 25000
rect 126200 25000 126300 25100
rect 126200 25100 126300 25200
rect 126200 25200 126300 25300
rect 126200 25300 126300 25400
rect 126200 25400 126300 25500
rect 126200 25500 126300 25600
rect 126200 25600 126300 25700
rect 126200 25700 126300 25800
rect 126200 25800 126300 25900
rect 126200 25900 126300 26000
rect 126200 26000 126300 26100
rect 126200 26100 126300 26200
rect 126200 26200 126300 26300
rect 126200 26300 126300 26400
rect 126200 26400 126300 26500
rect 126200 26500 126300 26600
rect 126200 26600 126300 26700
rect 126200 26700 126300 26800
rect 126200 26800 126300 26900
rect 126200 26900 126300 27000
rect 126200 27000 126300 27100
rect 126200 27100 126300 27200
rect 126300 21800 126400 21900
rect 126300 21900 126400 22000
rect 126300 22000 126400 22100
rect 126300 22100 126400 22200
rect 126300 22200 126400 22300
rect 126300 22300 126400 22400
rect 126300 22400 126400 22500
rect 126300 22500 126400 22600
rect 126300 22600 126400 22700
rect 126300 22700 126400 22800
rect 126300 22800 126400 22900
rect 126300 22900 126400 23000
rect 126300 23000 126400 23100
rect 126300 23100 126400 23200
rect 126300 23200 126400 23300
rect 126300 23300 126400 23400
rect 126300 24800 126400 24900
rect 126300 24900 126400 25000
rect 126300 25000 126400 25100
rect 126300 25100 126400 25200
rect 126300 25200 126400 25300
rect 126300 25300 126400 25400
rect 126300 25400 126400 25500
rect 126300 25500 126400 25600
rect 126300 25600 126400 25700
rect 126300 25700 126400 25800
rect 126300 25800 126400 25900
rect 126300 25900 126400 26000
rect 126300 26000 126400 26100
rect 126300 26100 126400 26200
rect 126300 26200 126400 26300
rect 126300 26300 126400 26400
rect 126300 26400 126400 26500
rect 126300 26500 126400 26600
rect 126300 26600 126400 26700
rect 126300 26700 126400 26800
rect 126300 26800 126400 26900
rect 126300 26900 126400 27000
rect 126400 21800 126500 21900
rect 126400 21900 126500 22000
rect 126400 22000 126500 22100
rect 126400 22100 126500 22200
rect 126400 22200 126500 22300
rect 126400 22300 126500 22400
rect 126400 22400 126500 22500
rect 126400 22500 126500 22600
rect 126400 22600 126500 22700
rect 126400 22700 126500 22800
rect 126400 22800 126500 22900
rect 126400 22900 126500 23000
rect 126400 23000 126500 23100
rect 126400 23100 126500 23200
rect 126400 23200 126500 23300
rect 126400 23300 126500 23400
rect 126400 24800 126500 24900
rect 126400 24900 126500 25000
rect 126400 25000 126500 25100
rect 126400 25100 126500 25200
rect 126400 25200 126500 25300
rect 126400 25300 126500 25400
rect 126400 25400 126500 25500
rect 126400 25500 126500 25600
rect 126400 25600 126500 25700
rect 126400 25700 126500 25800
rect 126400 25800 126500 25900
rect 126400 25900 126500 26000
rect 126400 26000 126500 26100
rect 126400 26100 126500 26200
rect 126400 26200 126500 26300
rect 126400 26300 126500 26400
rect 126400 26400 126500 26500
rect 126400 26500 126500 26600
rect 126400 26600 126500 26700
rect 126400 26700 126500 26800
rect 126400 26800 126500 26900
rect 126400 26900 126500 27000
rect 126400 27000 126500 27100
rect 126500 21800 126600 21900
rect 126500 21900 126600 22000
rect 126500 22000 126600 22100
rect 126500 22100 126600 22200
rect 126500 22200 126600 22300
rect 126500 22300 126600 22400
rect 126500 22400 126600 22500
rect 126500 22500 126600 22600
rect 126500 22600 126600 22700
rect 126500 22700 126600 22800
rect 126500 22800 126600 22900
rect 126500 22900 126600 23000
rect 126500 23000 126600 23100
rect 126500 23100 126600 23200
rect 126500 23200 126600 23300
rect 126500 23300 126600 23400
rect 126500 24700 126600 24800
rect 126500 24800 126600 24900
rect 126500 24900 126600 25000
rect 126500 25000 126600 25100
rect 126500 25100 126600 25200
rect 126500 25200 126600 25300
rect 126500 25300 126600 25400
rect 126500 25400 126600 25500
rect 126500 25500 126600 25600
rect 126500 25600 126600 25700
rect 126500 25700 126600 25800
rect 126500 25800 126600 25900
rect 126500 25900 126600 26000
rect 126500 26000 126600 26100
rect 126500 26100 126600 26200
rect 126500 26200 126600 26300
rect 126500 26300 126600 26400
rect 126500 26400 126600 26500
rect 126500 26500 126600 26600
rect 126500 26600 126600 26700
rect 126500 26700 126600 26800
rect 126500 26800 126600 26900
rect 126500 26900 126600 27000
rect 126500 27000 126600 27100
rect 126500 27100 126600 27200
rect 126500 27200 126600 27300
rect 126600 21800 126700 21900
rect 126600 21900 126700 22000
rect 126600 22000 126700 22100
rect 126600 22100 126700 22200
rect 126600 22200 126700 22300
rect 126600 22300 126700 22400
rect 126600 22400 126700 22500
rect 126600 22500 126700 22600
rect 126600 22600 126700 22700
rect 126600 22700 126700 22800
rect 126600 22800 126700 22900
rect 126600 22900 126700 23000
rect 126600 23000 126700 23100
rect 126600 23100 126700 23200
rect 126600 23200 126700 23300
rect 126600 23300 126700 23400
rect 126600 23400 126700 23500
rect 126600 24700 126700 24800
rect 126600 24800 126700 24900
rect 126600 24900 126700 25000
rect 126600 25000 126700 25100
rect 126600 25100 126700 25200
rect 126600 25200 126700 25300
rect 126600 25300 126700 25400
rect 126600 25400 126700 25500
rect 126600 25500 126700 25600
rect 126600 25600 126700 25700
rect 126600 25700 126700 25800
rect 126600 25800 126700 25900
rect 126600 25900 126700 26000
rect 126600 26000 126700 26100
rect 126600 26100 126700 26200
rect 126600 26200 126700 26300
rect 126600 26300 126700 26400
rect 126600 26400 126700 26500
rect 126600 26500 126700 26600
rect 126600 26600 126700 26700
rect 126600 26700 126700 26800
rect 126600 26800 126700 26900
rect 126600 26900 126700 27000
rect 126600 27000 126700 27100
rect 126600 27100 126700 27200
rect 126600 27200 126700 27300
rect 126600 27300 126700 27400
rect 126600 27400 126700 27500
rect 126600 27500 126700 27600
rect 126700 21800 126800 21900
rect 126700 21900 126800 22000
rect 126700 22000 126800 22100
rect 126700 22100 126800 22200
rect 126700 22200 126800 22300
rect 126700 22300 126800 22400
rect 126700 22400 126800 22500
rect 126700 22500 126800 22600
rect 126700 22600 126800 22700
rect 126700 22700 126800 22800
rect 126700 22800 126800 22900
rect 126700 22900 126800 23000
rect 126700 23000 126800 23100
rect 126700 23100 126800 23200
rect 126700 23200 126800 23300
rect 126700 23300 126800 23400
rect 126700 23400 126800 23500
rect 126700 23500 126800 23600
rect 126700 24600 126800 24700
rect 126700 24700 126800 24800
rect 126700 24800 126800 24900
rect 126700 24900 126800 25000
rect 126700 25000 126800 25100
rect 126700 25100 126800 25200
rect 126700 25200 126800 25300
rect 126700 25300 126800 25400
rect 126700 25400 126800 25500
rect 126700 25500 126800 25600
rect 126700 25600 126800 25700
rect 126700 25700 126800 25800
rect 126700 25800 126800 25900
rect 126700 25900 126800 26000
rect 126700 26000 126800 26100
rect 126700 26100 126800 26200
rect 126700 26200 126800 26300
rect 126700 26300 126800 26400
rect 126700 26400 126800 26500
rect 126700 26500 126800 26600
rect 126700 26600 126800 26700
rect 126700 26700 126800 26800
rect 126700 26800 126800 26900
rect 126700 26900 126800 27000
rect 126700 27000 126800 27100
rect 126700 27100 126800 27200
rect 126700 27200 126800 27300
rect 126700 27300 126800 27400
rect 126700 27400 126800 27500
rect 126700 27500 126800 27600
rect 126700 27600 126800 27700
rect 126700 27700 126800 27800
rect 126700 27800 126800 27900
rect 126800 21900 126900 22000
rect 126800 22000 126900 22100
rect 126800 22100 126900 22200
rect 126800 22200 126900 22300
rect 126800 22300 126900 22400
rect 126800 22400 126900 22500
rect 126800 22500 126900 22600
rect 126800 22600 126900 22700
rect 126800 22700 126900 22800
rect 126800 22800 126900 22900
rect 126800 22900 126900 23000
rect 126800 23000 126900 23100
rect 126800 23100 126900 23200
rect 126800 23200 126900 23300
rect 126800 23300 126900 23400
rect 126800 23400 126900 23500
rect 126800 23500 126900 23600
rect 126800 23600 126900 23700
rect 126800 24500 126900 24600
rect 126800 24600 126900 24700
rect 126800 24700 126900 24800
rect 126800 24800 126900 24900
rect 126800 24900 126900 25000
rect 126800 25000 126900 25100
rect 126800 25100 126900 25200
rect 126800 25200 126900 25300
rect 126800 25300 126900 25400
rect 126800 25400 126900 25500
rect 126800 25500 126900 25600
rect 126800 25600 126900 25700
rect 126800 25700 126900 25800
rect 126800 25800 126900 25900
rect 126800 25900 126900 26000
rect 126800 26000 126900 26100
rect 126800 26100 126900 26200
rect 126800 26200 126900 26300
rect 126800 26300 126900 26400
rect 126800 26400 126900 26500
rect 126800 26500 126900 26600
rect 126800 26600 126900 26700
rect 126800 26700 126900 26800
rect 126800 26800 126900 26900
rect 126800 26900 126900 27000
rect 126800 27000 126900 27100
rect 126800 27100 126900 27200
rect 126800 27200 126900 27300
rect 126800 27300 126900 27400
rect 126800 27400 126900 27500
rect 126800 27500 126900 27600
rect 126800 27600 126900 27700
rect 126800 27700 126900 27800
rect 126800 27800 126900 27900
rect 126800 27900 126900 28000
rect 126800 28000 126900 28100
rect 126800 28100 126900 28200
rect 126900 21900 127000 22000
rect 126900 22000 127000 22100
rect 126900 22100 127000 22200
rect 126900 22200 127000 22300
rect 126900 22300 127000 22400
rect 126900 22400 127000 22500
rect 126900 22500 127000 22600
rect 126900 22600 127000 22700
rect 126900 22700 127000 22800
rect 126900 22800 127000 22900
rect 126900 22900 127000 23000
rect 126900 23000 127000 23100
rect 126900 23100 127000 23200
rect 126900 23200 127000 23300
rect 126900 23300 127000 23400
rect 126900 23400 127000 23500
rect 126900 23500 127000 23600
rect 126900 23600 127000 23700
rect 126900 23700 127000 23800
rect 126900 24400 127000 24500
rect 126900 24500 127000 24600
rect 126900 24600 127000 24700
rect 126900 24700 127000 24800
rect 126900 24800 127000 24900
rect 126900 24900 127000 25000
rect 126900 25000 127000 25100
rect 126900 25100 127000 25200
rect 126900 25200 127000 25300
rect 126900 25300 127000 25400
rect 126900 25400 127000 25500
rect 126900 25500 127000 25600
rect 126900 25600 127000 25700
rect 126900 25700 127000 25800
rect 126900 25800 127000 25900
rect 126900 25900 127000 26000
rect 126900 26000 127000 26100
rect 126900 26100 127000 26200
rect 126900 26200 127000 26300
rect 126900 26300 127000 26400
rect 126900 26400 127000 26500
rect 126900 26500 127000 26600
rect 126900 26600 127000 26700
rect 126900 26700 127000 26800
rect 126900 26800 127000 26900
rect 126900 26900 127000 27000
rect 126900 27000 127000 27100
rect 126900 27100 127000 27200
rect 126900 27200 127000 27300
rect 126900 27300 127000 27400
rect 126900 27400 127000 27500
rect 126900 27500 127000 27600
rect 126900 27600 127000 27700
rect 126900 27700 127000 27800
rect 126900 27800 127000 27900
rect 126900 27900 127000 28000
rect 126900 28000 127000 28100
rect 126900 28100 127000 28200
rect 126900 28200 127000 28300
rect 126900 28300 127000 28400
rect 127000 21900 127100 22000
rect 127000 22000 127100 22100
rect 127000 22100 127100 22200
rect 127000 22200 127100 22300
rect 127000 22300 127100 22400
rect 127000 22400 127100 22500
rect 127000 22500 127100 22600
rect 127000 22600 127100 22700
rect 127000 22700 127100 22800
rect 127000 22800 127100 22900
rect 127000 22900 127100 23000
rect 127000 23000 127100 23100
rect 127000 23100 127100 23200
rect 127000 23200 127100 23300
rect 127000 23300 127100 23400
rect 127000 23400 127100 23500
rect 127000 23500 127100 23600
rect 127000 23600 127100 23700
rect 127000 23700 127100 23800
rect 127000 23800 127100 23900
rect 127000 23900 127100 24000
rect 127000 24000 127100 24100
rect 127000 24100 127100 24200
rect 127000 24200 127100 24300
rect 127000 24300 127100 24400
rect 127000 24400 127100 24500
rect 127000 24500 127100 24600
rect 127000 24600 127100 24700
rect 127000 24700 127100 24800
rect 127000 24800 127100 24900
rect 127000 24900 127100 25000
rect 127000 25000 127100 25100
rect 127000 25100 127100 25200
rect 127000 25200 127100 25300
rect 127000 25300 127100 25400
rect 127000 25400 127100 25500
rect 127000 25500 127100 25600
rect 127000 25600 127100 25700
rect 127000 25700 127100 25800
rect 127000 25800 127100 25900
rect 127000 25900 127100 26000
rect 127000 26000 127100 26100
rect 127000 26100 127100 26200
rect 127000 26200 127100 26300
rect 127000 26300 127100 26400
rect 127000 26400 127100 26500
rect 127000 26500 127100 26600
rect 127000 26600 127100 26700
rect 127000 26700 127100 26800
rect 127000 26800 127100 26900
rect 127000 26900 127100 27000
rect 127000 27000 127100 27100
rect 127000 27100 127100 27200
rect 127000 27200 127100 27300
rect 127000 27300 127100 27400
rect 127000 27400 127100 27500
rect 127000 27500 127100 27600
rect 127000 27600 127100 27700
rect 127000 27700 127100 27800
rect 127000 27800 127100 27900
rect 127000 27900 127100 28000
rect 127000 28000 127100 28100
rect 127000 28100 127100 28200
rect 127000 28200 127100 28300
rect 127000 28300 127100 28400
rect 127000 28400 127100 28500
rect 127000 28500 127100 28600
rect 127000 28600 127100 28700
rect 127100 22000 127200 22100
rect 127100 22100 127200 22200
rect 127100 22200 127200 22300
rect 127100 22300 127200 22400
rect 127100 22400 127200 22500
rect 127100 22500 127200 22600
rect 127100 22600 127200 22700
rect 127100 22700 127200 22800
rect 127100 22800 127200 22900
rect 127100 22900 127200 23000
rect 127100 23000 127200 23100
rect 127100 23100 127200 23200
rect 127100 23200 127200 23300
rect 127100 23300 127200 23400
rect 127100 23400 127200 23500
rect 127100 23500 127200 23600
rect 127100 23600 127200 23700
rect 127100 23700 127200 23800
rect 127100 23800 127200 23900
rect 127100 23900 127200 24000
rect 127100 24000 127200 24100
rect 127100 24100 127200 24200
rect 127100 24200 127200 24300
rect 127100 24300 127200 24400
rect 127100 24400 127200 24500
rect 127100 24500 127200 24600
rect 127100 24600 127200 24700
rect 127100 24700 127200 24800
rect 127100 24800 127200 24900
rect 127100 24900 127200 25000
rect 127100 25000 127200 25100
rect 127100 25100 127200 25200
rect 127100 25200 127200 25300
rect 127100 25300 127200 25400
rect 127100 25400 127200 25500
rect 127100 25500 127200 25600
rect 127100 25600 127200 25700
rect 127100 25700 127200 25800
rect 127100 25800 127200 25900
rect 127100 25900 127200 26000
rect 127100 26000 127200 26100
rect 127100 26100 127200 26200
rect 127100 26200 127200 26300
rect 127100 26300 127200 26400
rect 127100 26400 127200 26500
rect 127100 26500 127200 26600
rect 127100 26600 127200 26700
rect 127100 26700 127200 26800
rect 127100 26800 127200 26900
rect 127100 26900 127200 27000
rect 127100 27000 127200 27100
rect 127100 27100 127200 27200
rect 127100 27200 127200 27300
rect 127100 27300 127200 27400
rect 127100 27400 127200 27500
rect 127100 27500 127200 27600
rect 127100 27600 127200 27700
rect 127100 27700 127200 27800
rect 127100 27800 127200 27900
rect 127100 27900 127200 28000
rect 127100 28000 127200 28100
rect 127100 28100 127200 28200
rect 127100 28200 127200 28300
rect 127100 28300 127200 28400
rect 127100 28400 127200 28500
rect 127100 28500 127200 28600
rect 127100 28600 127200 28700
rect 127100 28700 127200 28800
rect 127100 28800 127200 28900
rect 127100 28900 127200 29000
rect 127200 22000 127300 22100
rect 127200 22100 127300 22200
rect 127200 22200 127300 22300
rect 127200 22300 127300 22400
rect 127200 22400 127300 22500
rect 127200 22500 127300 22600
rect 127200 22600 127300 22700
rect 127200 22700 127300 22800
rect 127200 22800 127300 22900
rect 127200 22900 127300 23000
rect 127200 23000 127300 23100
rect 127200 23100 127300 23200
rect 127200 23200 127300 23300
rect 127200 23300 127300 23400
rect 127200 23400 127300 23500
rect 127200 23500 127300 23600
rect 127200 23600 127300 23700
rect 127200 23700 127300 23800
rect 127200 23800 127300 23900
rect 127200 23900 127300 24000
rect 127200 24000 127300 24100
rect 127200 24100 127300 24200
rect 127200 24200 127300 24300
rect 127200 24300 127300 24400
rect 127200 24400 127300 24500
rect 127200 24500 127300 24600
rect 127200 24600 127300 24700
rect 127200 24700 127300 24800
rect 127200 24800 127300 24900
rect 127200 24900 127300 25000
rect 127200 25000 127300 25100
rect 127200 25100 127300 25200
rect 127200 25200 127300 25300
rect 127200 25300 127300 25400
rect 127200 25400 127300 25500
rect 127200 25500 127300 25600
rect 127200 25600 127300 25700
rect 127200 25700 127300 25800
rect 127200 25800 127300 25900
rect 127200 25900 127300 26000
rect 127200 26000 127300 26100
rect 127200 26100 127300 26200
rect 127200 26200 127300 26300
rect 127200 26300 127300 26400
rect 127200 26400 127300 26500
rect 127200 26500 127300 26600
rect 127200 26600 127300 26700
rect 127200 26700 127300 26800
rect 127200 26800 127300 26900
rect 127200 26900 127300 27000
rect 127200 27000 127300 27100
rect 127200 27100 127300 27200
rect 127200 27200 127300 27300
rect 127200 27300 127300 27400
rect 127200 27400 127300 27500
rect 127200 27500 127300 27600
rect 127200 27600 127300 27700
rect 127200 27700 127300 27800
rect 127200 27800 127300 27900
rect 127200 27900 127300 28000
rect 127200 28000 127300 28100
rect 127200 28100 127300 28200
rect 127200 28200 127300 28300
rect 127200 28300 127300 28400
rect 127200 28400 127300 28500
rect 127200 28500 127300 28600
rect 127200 28600 127300 28700
rect 127200 28700 127300 28800
rect 127200 28800 127300 28900
rect 127200 28900 127300 29000
rect 127200 29000 127300 29100
rect 127200 29100 127300 29200
rect 127200 29200 127300 29300
rect 127300 22100 127400 22200
rect 127300 22200 127400 22300
rect 127300 22300 127400 22400
rect 127300 22400 127400 22500
rect 127300 22500 127400 22600
rect 127300 22600 127400 22700
rect 127300 22700 127400 22800
rect 127300 22800 127400 22900
rect 127300 22900 127400 23000
rect 127300 23000 127400 23100
rect 127300 23100 127400 23200
rect 127300 23200 127400 23300
rect 127300 23300 127400 23400
rect 127300 23400 127400 23500
rect 127300 23500 127400 23600
rect 127300 23600 127400 23700
rect 127300 23700 127400 23800
rect 127300 23800 127400 23900
rect 127300 23900 127400 24000
rect 127300 24000 127400 24100
rect 127300 24100 127400 24200
rect 127300 24200 127400 24300
rect 127300 24300 127400 24400
rect 127300 24400 127400 24500
rect 127300 24500 127400 24600
rect 127300 24600 127400 24700
rect 127300 24700 127400 24800
rect 127300 24800 127400 24900
rect 127300 24900 127400 25000
rect 127300 25000 127400 25100
rect 127300 25100 127400 25200
rect 127300 25200 127400 25300
rect 127300 25300 127400 25400
rect 127300 25400 127400 25500
rect 127300 25500 127400 25600
rect 127300 25600 127400 25700
rect 127300 25700 127400 25800
rect 127300 25800 127400 25900
rect 127300 25900 127400 26000
rect 127300 26000 127400 26100
rect 127300 26100 127400 26200
rect 127300 26200 127400 26300
rect 127300 26300 127400 26400
rect 127300 26400 127400 26500
rect 127300 26500 127400 26600
rect 127300 26600 127400 26700
rect 127300 26700 127400 26800
rect 127300 26800 127400 26900
rect 127300 26900 127400 27000
rect 127300 27000 127400 27100
rect 127300 27100 127400 27200
rect 127300 27200 127400 27300
rect 127300 27300 127400 27400
rect 127300 27400 127400 27500
rect 127300 27500 127400 27600
rect 127300 27600 127400 27700
rect 127300 27700 127400 27800
rect 127300 27800 127400 27900
rect 127300 27900 127400 28000
rect 127300 28000 127400 28100
rect 127300 28100 127400 28200
rect 127300 28200 127400 28300
rect 127300 28300 127400 28400
rect 127300 28400 127400 28500
rect 127300 28500 127400 28600
rect 127300 28600 127400 28700
rect 127300 28700 127400 28800
rect 127300 28800 127400 28900
rect 127300 28900 127400 29000
rect 127300 29000 127400 29100
rect 127300 29100 127400 29200
rect 127300 29200 127400 29300
rect 127300 29300 127400 29400
rect 127300 29400 127400 29500
rect 127400 22100 127500 22200
rect 127400 22200 127500 22300
rect 127400 22300 127500 22400
rect 127400 22400 127500 22500
rect 127400 22500 127500 22600
rect 127400 22600 127500 22700
rect 127400 22700 127500 22800
rect 127400 22800 127500 22900
rect 127400 22900 127500 23000
rect 127400 23000 127500 23100
rect 127400 23100 127500 23200
rect 127400 23200 127500 23300
rect 127400 23300 127500 23400
rect 127400 23400 127500 23500
rect 127400 23500 127500 23600
rect 127400 23600 127500 23700
rect 127400 23700 127500 23800
rect 127400 23800 127500 23900
rect 127400 23900 127500 24000
rect 127400 24000 127500 24100
rect 127400 24100 127500 24200
rect 127400 24200 127500 24300
rect 127400 24300 127500 24400
rect 127400 24400 127500 24500
rect 127400 24500 127500 24600
rect 127400 24600 127500 24700
rect 127400 24700 127500 24800
rect 127400 24800 127500 24900
rect 127400 24900 127500 25000
rect 127400 25000 127500 25100
rect 127400 25100 127500 25200
rect 127400 25200 127500 25300
rect 127400 25300 127500 25400
rect 127400 25400 127500 25500
rect 127400 25500 127500 25600
rect 127400 25600 127500 25700
rect 127400 25700 127500 25800
rect 127400 25800 127500 25900
rect 127400 25900 127500 26000
rect 127400 26000 127500 26100
rect 127400 26100 127500 26200
rect 127400 26200 127500 26300
rect 127400 26300 127500 26400
rect 127400 26400 127500 26500
rect 127400 26500 127500 26600
rect 127400 26600 127500 26700
rect 127400 26700 127500 26800
rect 127400 26800 127500 26900
rect 127400 26900 127500 27000
rect 127400 27000 127500 27100
rect 127400 27100 127500 27200
rect 127400 27200 127500 27300
rect 127400 27300 127500 27400
rect 127400 27400 127500 27500
rect 127400 27500 127500 27600
rect 127400 27600 127500 27700
rect 127400 27700 127500 27800
rect 127400 27800 127500 27900
rect 127400 27900 127500 28000
rect 127400 28000 127500 28100
rect 127400 28100 127500 28200
rect 127400 28200 127500 28300
rect 127400 28300 127500 28400
rect 127400 28400 127500 28500
rect 127400 28500 127500 28600
rect 127400 28600 127500 28700
rect 127400 28700 127500 28800
rect 127400 28800 127500 28900
rect 127400 28900 127500 29000
rect 127400 29000 127500 29100
rect 127400 29100 127500 29200
rect 127400 29200 127500 29300
rect 127400 29300 127500 29400
rect 127400 29400 127500 29500
rect 127400 29500 127500 29600
rect 127400 29600 127500 29700
rect 127400 29700 127500 29800
rect 127500 22200 127600 22300
rect 127500 22300 127600 22400
rect 127500 22400 127600 22500
rect 127500 22500 127600 22600
rect 127500 22600 127600 22700
rect 127500 22700 127600 22800
rect 127500 22800 127600 22900
rect 127500 22900 127600 23000
rect 127500 23000 127600 23100
rect 127500 23100 127600 23200
rect 127500 23200 127600 23300
rect 127500 23300 127600 23400
rect 127500 23400 127600 23500
rect 127500 23500 127600 23600
rect 127500 23600 127600 23700
rect 127500 23700 127600 23800
rect 127500 23800 127600 23900
rect 127500 23900 127600 24000
rect 127500 24000 127600 24100
rect 127500 24100 127600 24200
rect 127500 24200 127600 24300
rect 127500 24300 127600 24400
rect 127500 24400 127600 24500
rect 127500 24500 127600 24600
rect 127500 24600 127600 24700
rect 127500 24700 127600 24800
rect 127500 24800 127600 24900
rect 127500 24900 127600 25000
rect 127500 25000 127600 25100
rect 127500 25100 127600 25200
rect 127500 25200 127600 25300
rect 127500 25300 127600 25400
rect 127500 25400 127600 25500
rect 127500 25500 127600 25600
rect 127500 25600 127600 25700
rect 127500 25700 127600 25800
rect 127500 25800 127600 25900
rect 127500 25900 127600 26000
rect 127500 26000 127600 26100
rect 127500 26100 127600 26200
rect 127500 26200 127600 26300
rect 127500 26300 127600 26400
rect 127500 26400 127600 26500
rect 127500 26500 127600 26600
rect 127500 26600 127600 26700
rect 127500 26700 127600 26800
rect 127500 26800 127600 26900
rect 127500 26900 127600 27000
rect 127500 27000 127600 27100
rect 127500 27100 127600 27200
rect 127500 27200 127600 27300
rect 127500 27300 127600 27400
rect 127500 27400 127600 27500
rect 127500 27500 127600 27600
rect 127500 27600 127600 27700
rect 127500 27700 127600 27800
rect 127500 27800 127600 27900
rect 127500 27900 127600 28000
rect 127500 28000 127600 28100
rect 127500 28100 127600 28200
rect 127500 28200 127600 28300
rect 127500 28300 127600 28400
rect 127500 28400 127600 28500
rect 127500 28500 127600 28600
rect 127500 28600 127600 28700
rect 127500 28700 127600 28800
rect 127500 28800 127600 28900
rect 127500 28900 127600 29000
rect 127500 29000 127600 29100
rect 127500 29100 127600 29200
rect 127500 29200 127600 29300
rect 127500 29300 127600 29400
rect 127500 29400 127600 29500
rect 127500 29500 127600 29600
rect 127500 29600 127600 29700
rect 127500 29700 127600 29800
rect 127500 29800 127600 29900
rect 127500 29900 127600 30000
rect 127500 30000 127600 30100
rect 127600 22200 127700 22300
rect 127600 22300 127700 22400
rect 127600 22400 127700 22500
rect 127600 22500 127700 22600
rect 127600 22600 127700 22700
rect 127600 22700 127700 22800
rect 127600 22800 127700 22900
rect 127600 22900 127700 23000
rect 127600 23000 127700 23100
rect 127600 23100 127700 23200
rect 127600 23200 127700 23300
rect 127600 23300 127700 23400
rect 127600 23400 127700 23500
rect 127600 23500 127700 23600
rect 127600 23600 127700 23700
rect 127600 23700 127700 23800
rect 127600 23800 127700 23900
rect 127600 23900 127700 24000
rect 127600 24000 127700 24100
rect 127600 24100 127700 24200
rect 127600 24200 127700 24300
rect 127600 24300 127700 24400
rect 127600 24400 127700 24500
rect 127600 24500 127700 24600
rect 127600 24600 127700 24700
rect 127600 24700 127700 24800
rect 127600 24800 127700 24900
rect 127600 24900 127700 25000
rect 127600 25000 127700 25100
rect 127600 25100 127700 25200
rect 127600 25200 127700 25300
rect 127600 25300 127700 25400
rect 127600 25400 127700 25500
rect 127600 25500 127700 25600
rect 127600 25600 127700 25700
rect 127600 25700 127700 25800
rect 127600 25800 127700 25900
rect 127600 25900 127700 26000
rect 127600 26000 127700 26100
rect 127600 26100 127700 26200
rect 127600 26200 127700 26300
rect 127600 26300 127700 26400
rect 127600 26400 127700 26500
rect 127600 26500 127700 26600
rect 127600 26600 127700 26700
rect 127600 26700 127700 26800
rect 127600 26800 127700 26900
rect 127600 26900 127700 27000
rect 127600 27000 127700 27100
rect 127600 27100 127700 27200
rect 127600 27200 127700 27300
rect 127600 27300 127700 27400
rect 127600 27400 127700 27500
rect 127600 27500 127700 27600
rect 127600 27600 127700 27700
rect 127600 27700 127700 27800
rect 127600 27800 127700 27900
rect 127600 27900 127700 28000
rect 127600 28000 127700 28100
rect 127600 28100 127700 28200
rect 127600 28200 127700 28300
rect 127600 28300 127700 28400
rect 127600 28400 127700 28500
rect 127600 28500 127700 28600
rect 127600 28600 127700 28700
rect 127600 28700 127700 28800
rect 127600 28800 127700 28900
rect 127600 28900 127700 29000
rect 127600 29000 127700 29100
rect 127600 29100 127700 29200
rect 127600 29200 127700 29300
rect 127600 29300 127700 29400
rect 127600 29400 127700 29500
rect 127600 29500 127700 29600
rect 127600 29600 127700 29700
rect 127600 29700 127700 29800
rect 127600 29800 127700 29900
rect 127600 29900 127700 30000
rect 127600 30000 127700 30100
rect 127600 30100 127700 30200
rect 127600 30200 127700 30300
rect 127600 30300 127700 30400
rect 127700 22300 127800 22400
rect 127700 22400 127800 22500
rect 127700 22500 127800 22600
rect 127700 22600 127800 22700
rect 127700 22700 127800 22800
rect 127700 22800 127800 22900
rect 127700 22900 127800 23000
rect 127700 23000 127800 23100
rect 127700 23100 127800 23200
rect 127700 23200 127800 23300
rect 127700 23300 127800 23400
rect 127700 23400 127800 23500
rect 127700 23500 127800 23600
rect 127700 23600 127800 23700
rect 127700 23700 127800 23800
rect 127700 23800 127800 23900
rect 127700 23900 127800 24000
rect 127700 24000 127800 24100
rect 127700 24100 127800 24200
rect 127700 24200 127800 24300
rect 127700 24300 127800 24400
rect 127700 24400 127800 24500
rect 127700 24500 127800 24600
rect 127700 24600 127800 24700
rect 127700 24700 127800 24800
rect 127700 24800 127800 24900
rect 127700 24900 127800 25000
rect 127700 25000 127800 25100
rect 127700 25100 127800 25200
rect 127700 25200 127800 25300
rect 127700 25300 127800 25400
rect 127700 25400 127800 25500
rect 127700 25500 127800 25600
rect 127700 25600 127800 25700
rect 127700 25700 127800 25800
rect 127700 25800 127800 25900
rect 127700 25900 127800 26000
rect 127700 26000 127800 26100
rect 127700 26100 127800 26200
rect 127700 26200 127800 26300
rect 127700 26300 127800 26400
rect 127700 26400 127800 26500
rect 127700 26500 127800 26600
rect 127700 26600 127800 26700
rect 127700 26700 127800 26800
rect 127700 26800 127800 26900
rect 127700 26900 127800 27000
rect 127700 27000 127800 27100
rect 127700 27100 127800 27200
rect 127700 27200 127800 27300
rect 127700 27300 127800 27400
rect 127700 27400 127800 27500
rect 127700 27500 127800 27600
rect 127700 27600 127800 27700
rect 127700 27700 127800 27800
rect 127700 27800 127800 27900
rect 127700 27900 127800 28000
rect 127700 28000 127800 28100
rect 127700 28100 127800 28200
rect 127700 28200 127800 28300
rect 127700 28300 127800 28400
rect 127700 28400 127800 28500
rect 127700 28500 127800 28600
rect 127700 28600 127800 28700
rect 127700 28700 127800 28800
rect 127700 28800 127800 28900
rect 127700 28900 127800 29000
rect 127700 29000 127800 29100
rect 127700 29100 127800 29200
rect 127700 29200 127800 29300
rect 127700 29300 127800 29400
rect 127700 29400 127800 29500
rect 127700 29500 127800 29600
rect 127700 29600 127800 29700
rect 127700 29700 127800 29800
rect 127700 29800 127800 29900
rect 127700 29900 127800 30000
rect 127700 30000 127800 30100
rect 127700 30100 127800 30200
rect 127700 30200 127800 30300
rect 127700 30300 127800 30400
rect 127700 30400 127800 30500
rect 127700 30500 127800 30600
rect 127700 30600 127800 30700
rect 127800 22400 127900 22500
rect 127800 22500 127900 22600
rect 127800 22600 127900 22700
rect 127800 22700 127900 22800
rect 127800 22800 127900 22900
rect 127800 22900 127900 23000
rect 127800 23000 127900 23100
rect 127800 23100 127900 23200
rect 127800 23200 127900 23300
rect 127800 23300 127900 23400
rect 127800 23400 127900 23500
rect 127800 23500 127900 23600
rect 127800 23600 127900 23700
rect 127800 23700 127900 23800
rect 127800 23800 127900 23900
rect 127800 23900 127900 24000
rect 127800 24000 127900 24100
rect 127800 24100 127900 24200
rect 127800 24200 127900 24300
rect 127800 24300 127900 24400
rect 127800 24400 127900 24500
rect 127800 24500 127900 24600
rect 127800 24600 127900 24700
rect 127800 24700 127900 24800
rect 127800 24800 127900 24900
rect 127800 24900 127900 25000
rect 127800 25000 127900 25100
rect 127800 25100 127900 25200
rect 127800 25200 127900 25300
rect 127800 25300 127900 25400
rect 127800 25400 127900 25500
rect 127800 25500 127900 25600
rect 127800 25600 127900 25700
rect 127800 25700 127900 25800
rect 127800 25800 127900 25900
rect 127800 25900 127900 26000
rect 127800 26000 127900 26100
rect 127800 26100 127900 26200
rect 127800 26200 127900 26300
rect 127800 26300 127900 26400
rect 127800 26400 127900 26500
rect 127800 26500 127900 26600
rect 127800 26600 127900 26700
rect 127800 26700 127900 26800
rect 127800 26800 127900 26900
rect 127800 26900 127900 27000
rect 127800 27000 127900 27100
rect 127800 27100 127900 27200
rect 127800 27200 127900 27300
rect 127800 27300 127900 27400
rect 127800 27400 127900 27500
rect 127800 27500 127900 27600
rect 127800 27600 127900 27700
rect 127800 27700 127900 27800
rect 127800 27800 127900 27900
rect 127800 27900 127900 28000
rect 127800 28000 127900 28100
rect 127800 28100 127900 28200
rect 127800 28200 127900 28300
rect 127800 28300 127900 28400
rect 127800 28400 127900 28500
rect 127800 28500 127900 28600
rect 127800 28600 127900 28700
rect 127800 28700 127900 28800
rect 127800 28800 127900 28900
rect 127800 28900 127900 29000
rect 127800 29000 127900 29100
rect 127800 29100 127900 29200
rect 127800 29200 127900 29300
rect 127800 29300 127900 29400
rect 127800 29400 127900 29500
rect 127800 29500 127900 29600
rect 127800 29600 127900 29700
rect 127800 29700 127900 29800
rect 127800 29800 127900 29900
rect 127800 29900 127900 30000
rect 127800 30000 127900 30100
rect 127800 30100 127900 30200
rect 127800 30200 127900 30300
rect 127800 30300 127900 30400
rect 127800 30400 127900 30500
rect 127800 30500 127900 30600
rect 127800 30600 127900 30700
rect 127800 30700 127900 30800
rect 127800 30800 127900 30900
rect 127800 30900 127900 31000
rect 127900 22500 128000 22600
rect 127900 22600 128000 22700
rect 127900 22700 128000 22800
rect 127900 22800 128000 22900
rect 127900 22900 128000 23000
rect 127900 23000 128000 23100
rect 127900 23100 128000 23200
rect 127900 23200 128000 23300
rect 127900 23300 128000 23400
rect 127900 23400 128000 23500
rect 127900 23500 128000 23600
rect 127900 23600 128000 23700
rect 127900 23700 128000 23800
rect 127900 23800 128000 23900
rect 127900 23900 128000 24000
rect 127900 24000 128000 24100
rect 127900 24100 128000 24200
rect 127900 24200 128000 24300
rect 127900 24300 128000 24400
rect 127900 24400 128000 24500
rect 127900 24500 128000 24600
rect 127900 24600 128000 24700
rect 127900 24700 128000 24800
rect 127900 24800 128000 24900
rect 127900 24900 128000 25000
rect 127900 25000 128000 25100
rect 127900 25100 128000 25200
rect 127900 25200 128000 25300
rect 127900 25300 128000 25400
rect 127900 25400 128000 25500
rect 127900 25500 128000 25600
rect 127900 25600 128000 25700
rect 127900 25700 128000 25800
rect 127900 25800 128000 25900
rect 127900 26200 128000 26300
rect 127900 26300 128000 26400
rect 127900 26400 128000 26500
rect 127900 26500 128000 26600
rect 127900 26600 128000 26700
rect 127900 26700 128000 26800
rect 127900 26800 128000 26900
rect 127900 26900 128000 27000
rect 127900 27000 128000 27100
rect 127900 27100 128000 27200
rect 127900 27200 128000 27300
rect 127900 27300 128000 27400
rect 127900 27400 128000 27500
rect 127900 27500 128000 27600
rect 127900 27600 128000 27700
rect 127900 27700 128000 27800
rect 127900 27800 128000 27900
rect 127900 27900 128000 28000
rect 127900 28000 128000 28100
rect 127900 28100 128000 28200
rect 127900 28200 128000 28300
rect 127900 28300 128000 28400
rect 127900 28400 128000 28500
rect 127900 28500 128000 28600
rect 127900 28600 128000 28700
rect 127900 28700 128000 28800
rect 127900 28800 128000 28900
rect 127900 28900 128000 29000
rect 127900 29000 128000 29100
rect 127900 29100 128000 29200
rect 127900 29200 128000 29300
rect 127900 29300 128000 29400
rect 127900 29400 128000 29500
rect 127900 29500 128000 29600
rect 127900 29600 128000 29700
rect 127900 29700 128000 29800
rect 127900 29800 128000 29900
rect 127900 29900 128000 30000
rect 127900 30000 128000 30100
rect 127900 30100 128000 30200
rect 127900 30200 128000 30300
rect 127900 30300 128000 30400
rect 127900 30400 128000 30500
rect 127900 30500 128000 30600
rect 127900 30600 128000 30700
rect 127900 30700 128000 30800
rect 127900 30800 128000 30900
rect 127900 30900 128000 31000
rect 127900 31000 128000 31100
rect 127900 31100 128000 31200
rect 127900 31200 128000 31300
rect 128000 22600 128100 22700
rect 128000 22700 128100 22800
rect 128000 22800 128100 22900
rect 128000 22900 128100 23000
rect 128000 23000 128100 23100
rect 128000 23100 128100 23200
rect 128000 23200 128100 23300
rect 128000 23300 128100 23400
rect 128000 23400 128100 23500
rect 128000 23500 128100 23600
rect 128000 23600 128100 23700
rect 128000 23700 128100 23800
rect 128000 23800 128100 23900
rect 128000 23900 128100 24000
rect 128000 24000 128100 24100
rect 128000 24100 128100 24200
rect 128000 24200 128100 24300
rect 128000 24300 128100 24400
rect 128000 24400 128100 24500
rect 128000 24500 128100 24600
rect 128000 24600 128100 24700
rect 128000 24700 128100 24800
rect 128000 24800 128100 24900
rect 128000 24900 128100 25000
rect 128000 25000 128100 25100
rect 128000 25100 128100 25200
rect 128000 25200 128100 25300
rect 128000 25300 128100 25400
rect 128000 25400 128100 25500
rect 128000 25500 128100 25600
rect 128000 25600 128100 25700
rect 128000 25700 128100 25800
rect 128000 26500 128100 26600
rect 128000 26600 128100 26700
rect 128000 26700 128100 26800
rect 128000 26800 128100 26900
rect 128000 26900 128100 27000
rect 128000 27000 128100 27100
rect 128000 27100 128100 27200
rect 128000 27200 128100 27300
rect 128000 27300 128100 27400
rect 128000 27400 128100 27500
rect 128000 27500 128100 27600
rect 128000 27600 128100 27700
rect 128000 27700 128100 27800
rect 128000 27800 128100 27900
rect 128000 27900 128100 28000
rect 128000 28000 128100 28100
rect 128000 28100 128100 28200
rect 128000 28200 128100 28300
rect 128000 28300 128100 28400
rect 128000 28400 128100 28500
rect 128000 28500 128100 28600
rect 128000 28600 128100 28700
rect 128000 28700 128100 28800
rect 128000 28800 128100 28900
rect 128000 28900 128100 29000
rect 128000 29000 128100 29100
rect 128000 29100 128100 29200
rect 128000 29200 128100 29300
rect 128000 29300 128100 29400
rect 128000 29400 128100 29500
rect 128000 29500 128100 29600
rect 128000 29600 128100 29700
rect 128000 29700 128100 29800
rect 128000 29800 128100 29900
rect 128000 29900 128100 30000
rect 128000 30000 128100 30100
rect 128000 30100 128100 30200
rect 128000 30200 128100 30300
rect 128000 30300 128100 30400
rect 128000 30400 128100 30500
rect 128000 30500 128100 30600
rect 128000 30600 128100 30700
rect 128000 30700 128100 30800
rect 128000 30800 128100 30900
rect 128000 30900 128100 31000
rect 128000 31000 128100 31100
rect 128000 31100 128100 31200
rect 128000 31200 128100 31300
rect 128000 31300 128100 31400
rect 128000 31400 128100 31500
rect 128100 22700 128200 22800
rect 128100 22800 128200 22900
rect 128100 22900 128200 23000
rect 128100 23000 128200 23100
rect 128100 23100 128200 23200
rect 128100 23200 128200 23300
rect 128100 23300 128200 23400
rect 128100 23400 128200 23500
rect 128100 23500 128200 23600
rect 128100 23600 128200 23700
rect 128100 23700 128200 23800
rect 128100 23800 128200 23900
rect 128100 23900 128200 24000
rect 128100 24000 128200 24100
rect 128100 24100 128200 24200
rect 128100 24200 128200 24300
rect 128100 24300 128200 24400
rect 128100 24400 128200 24500
rect 128100 24500 128200 24600
rect 128100 24600 128200 24700
rect 128100 24700 128200 24800
rect 128100 24800 128200 24900
rect 128100 24900 128200 25000
rect 128100 25000 128200 25100
rect 128100 25100 128200 25200
rect 128100 25200 128200 25300
rect 128100 25300 128200 25400
rect 128100 25400 128200 25500
rect 128100 25500 128200 25600
rect 128100 25600 128200 25700
rect 128100 26800 128200 26900
rect 128100 26900 128200 27000
rect 128100 27000 128200 27100
rect 128100 27100 128200 27200
rect 128100 27200 128200 27300
rect 128100 27300 128200 27400
rect 128100 27400 128200 27500
rect 128100 27500 128200 27600
rect 128100 27600 128200 27700
rect 128100 27700 128200 27800
rect 128100 27800 128200 27900
rect 128100 27900 128200 28000
rect 128100 28000 128200 28100
rect 128100 28100 128200 28200
rect 128100 28200 128200 28300
rect 128100 28300 128200 28400
rect 128100 28400 128200 28500
rect 128100 28500 128200 28600
rect 128100 28600 128200 28700
rect 128100 28700 128200 28800
rect 128100 28800 128200 28900
rect 128100 28900 128200 29000
rect 128100 29000 128200 29100
rect 128100 29100 128200 29200
rect 128100 29200 128200 29300
rect 128100 29300 128200 29400
rect 128100 29400 128200 29500
rect 128100 29500 128200 29600
rect 128100 29600 128200 29700
rect 128100 29700 128200 29800
rect 128100 29800 128200 29900
rect 128100 29900 128200 30000
rect 128100 30000 128200 30100
rect 128100 30100 128200 30200
rect 128100 30200 128200 30300
rect 128100 30300 128200 30400
rect 128100 30400 128200 30500
rect 128100 30500 128200 30600
rect 128100 30600 128200 30700
rect 128100 30700 128200 30800
rect 128100 30800 128200 30900
rect 128100 30900 128200 31000
rect 128100 31000 128200 31100
rect 128100 31100 128200 31200
rect 128100 31200 128200 31300
rect 128100 31300 128200 31400
rect 128100 31400 128200 31500
rect 128100 31500 128200 31600
rect 128100 31600 128200 31700
rect 128100 31700 128200 31800
rect 128200 22800 128300 22900
rect 128200 22900 128300 23000
rect 128200 23000 128300 23100
rect 128200 23100 128300 23200
rect 128200 23200 128300 23300
rect 128200 23300 128300 23400
rect 128200 23400 128300 23500
rect 128200 23500 128300 23600
rect 128200 23600 128300 23700
rect 128200 23700 128300 23800
rect 128200 23800 128300 23900
rect 128200 23900 128300 24000
rect 128200 24000 128300 24100
rect 128200 24100 128300 24200
rect 128200 24200 128300 24300
rect 128200 24300 128300 24400
rect 128200 24400 128300 24500
rect 128200 24500 128300 24600
rect 128200 24600 128300 24700
rect 128200 24700 128300 24800
rect 128200 24800 128300 24900
rect 128200 24900 128300 25000
rect 128200 25000 128300 25100
rect 128200 25100 128300 25200
rect 128200 25200 128300 25300
rect 128200 25300 128300 25400
rect 128200 25400 128300 25500
rect 128200 27100 128300 27200
rect 128200 27200 128300 27300
rect 128200 27300 128300 27400
rect 128200 27400 128300 27500
rect 128200 27500 128300 27600
rect 128200 27600 128300 27700
rect 128200 27700 128300 27800
rect 128200 27800 128300 27900
rect 128200 27900 128300 28000
rect 128200 28000 128300 28100
rect 128200 28100 128300 28200
rect 128200 28200 128300 28300
rect 128200 28300 128300 28400
rect 128200 28400 128300 28500
rect 128200 28500 128300 28600
rect 128200 28600 128300 28700
rect 128200 28700 128300 28800
rect 128200 28800 128300 28900
rect 128200 28900 128300 29000
rect 128200 29000 128300 29100
rect 128200 29100 128300 29200
rect 128200 29200 128300 29300
rect 128200 29300 128300 29400
rect 128200 29400 128300 29500
rect 128200 29500 128300 29600
rect 128200 29600 128300 29700
rect 128200 29700 128300 29800
rect 128200 29800 128300 29900
rect 128200 29900 128300 30000
rect 128200 30000 128300 30100
rect 128200 30100 128300 30200
rect 128200 30200 128300 30300
rect 128200 30300 128300 30400
rect 128200 30400 128300 30500
rect 128200 30500 128300 30600
rect 128200 30600 128300 30700
rect 128200 30700 128300 30800
rect 128200 30800 128300 30900
rect 128200 30900 128300 31000
rect 128200 31000 128300 31100
rect 128200 31100 128300 31200
rect 128200 31200 128300 31300
rect 128200 31300 128300 31400
rect 128200 31400 128300 31500
rect 128200 31500 128300 31600
rect 128200 31600 128300 31700
rect 128200 31700 128300 31800
rect 128200 31800 128300 31900
rect 128200 31900 128300 32000
rect 128200 32000 128300 32100
rect 128300 23000 128400 23100
rect 128300 23100 128400 23200
rect 128300 23200 128400 23300
rect 128300 23300 128400 23400
rect 128300 23400 128400 23500
rect 128300 23500 128400 23600
rect 128300 23600 128400 23700
rect 128300 23700 128400 23800
rect 128300 23800 128400 23900
rect 128300 23900 128400 24000
rect 128300 24000 128400 24100
rect 128300 24100 128400 24200
rect 128300 24200 128400 24300
rect 128300 24300 128400 24400
rect 128300 24400 128400 24500
rect 128300 24500 128400 24600
rect 128300 24600 128400 24700
rect 128300 24700 128400 24800
rect 128300 24800 128400 24900
rect 128300 24900 128400 25000
rect 128300 25000 128400 25100
rect 128300 25100 128400 25200
rect 128300 25200 128400 25300
rect 128300 25300 128400 25400
rect 128300 27400 128400 27500
rect 128300 27500 128400 27600
rect 128300 27600 128400 27700
rect 128300 27700 128400 27800
rect 128300 27800 128400 27900
rect 128300 27900 128400 28000
rect 128300 28000 128400 28100
rect 128300 28100 128400 28200
rect 128300 28200 128400 28300
rect 128300 28300 128400 28400
rect 128300 28400 128400 28500
rect 128300 28500 128400 28600
rect 128300 28600 128400 28700
rect 128300 28700 128400 28800
rect 128300 28800 128400 28900
rect 128300 28900 128400 29000
rect 128300 29000 128400 29100
rect 128300 29100 128400 29200
rect 128300 29200 128400 29300
rect 128300 29300 128400 29400
rect 128300 29400 128400 29500
rect 128300 29500 128400 29600
rect 128300 29600 128400 29700
rect 128300 29700 128400 29800
rect 128300 29800 128400 29900
rect 128300 29900 128400 30000
rect 128300 30000 128400 30100
rect 128300 30100 128400 30200
rect 128300 30200 128400 30300
rect 128300 30300 128400 30400
rect 128300 30400 128400 30500
rect 128300 30500 128400 30600
rect 128300 30600 128400 30700
rect 128300 30700 128400 30800
rect 128300 30800 128400 30900
rect 128300 30900 128400 31000
rect 128300 31000 128400 31100
rect 128300 31100 128400 31200
rect 128300 31200 128400 31300
rect 128300 31300 128400 31400
rect 128300 31400 128400 31500
rect 128300 31500 128400 31600
rect 128300 31600 128400 31700
rect 128300 31700 128400 31800
rect 128300 31800 128400 31900
rect 128300 31900 128400 32000
rect 128300 32000 128400 32100
rect 128300 32100 128400 32200
rect 128300 32200 128400 32300
rect 128300 32300 128400 32400
rect 128400 23200 128500 23300
rect 128400 23300 128500 23400
rect 128400 23400 128500 23500
rect 128400 23500 128500 23600
rect 128400 23600 128500 23700
rect 128400 23700 128500 23800
rect 128400 23800 128500 23900
rect 128400 23900 128500 24000
rect 128400 24000 128500 24100
rect 128400 24100 128500 24200
rect 128400 24200 128500 24300
rect 128400 24300 128500 24400
rect 128400 24400 128500 24500
rect 128400 24500 128500 24600
rect 128400 24600 128500 24700
rect 128400 24700 128500 24800
rect 128400 24800 128500 24900
rect 128400 24900 128500 25000
rect 128400 25000 128500 25100
rect 128400 25100 128500 25200
rect 128400 27600 128500 27700
rect 128400 27700 128500 27800
rect 128400 27800 128500 27900
rect 128400 27900 128500 28000
rect 128400 28000 128500 28100
rect 128400 28100 128500 28200
rect 128400 28200 128500 28300
rect 128400 28300 128500 28400
rect 128400 28400 128500 28500
rect 128400 28500 128500 28600
rect 128400 28600 128500 28700
rect 128400 28700 128500 28800
rect 128400 28800 128500 28900
rect 128400 28900 128500 29000
rect 128400 29000 128500 29100
rect 128400 29100 128500 29200
rect 128400 29200 128500 29300
rect 128400 29300 128500 29400
rect 128400 29400 128500 29500
rect 128400 29500 128500 29600
rect 128400 29600 128500 29700
rect 128400 29700 128500 29800
rect 128400 29800 128500 29900
rect 128400 29900 128500 30000
rect 128400 30000 128500 30100
rect 128400 30100 128500 30200
rect 128400 30200 128500 30300
rect 128400 30300 128500 30400
rect 128400 30400 128500 30500
rect 128400 30500 128500 30600
rect 128400 30600 128500 30700
rect 128400 30700 128500 30800
rect 128400 30800 128500 30900
rect 128400 30900 128500 31000
rect 128400 31000 128500 31100
rect 128400 31100 128500 31200
rect 128400 31200 128500 31300
rect 128400 31300 128500 31400
rect 128400 31400 128500 31500
rect 128400 31500 128500 31600
rect 128400 31600 128500 31700
rect 128400 31700 128500 31800
rect 128400 31800 128500 31900
rect 128400 31900 128500 32000
rect 128400 32000 128500 32100
rect 128400 32100 128500 32200
rect 128400 32200 128500 32300
rect 128400 32300 128500 32400
rect 128400 32400 128500 32500
rect 128400 32500 128500 32600
rect 128400 32600 128500 32700
rect 128500 23500 128600 23600
rect 128500 23600 128600 23700
rect 128500 23700 128600 23800
rect 128500 23800 128600 23900
rect 128500 23900 128600 24000
rect 128500 24000 128600 24100
rect 128500 24100 128600 24200
rect 128500 24200 128600 24300
rect 128500 24300 128600 24400
rect 128500 24400 128600 24500
rect 128500 24500 128600 24600
rect 128500 24600 128600 24700
rect 128500 24700 128600 24800
rect 128500 24800 128600 24900
rect 128500 27900 128600 28000
rect 128500 28000 128600 28100
rect 128500 28100 128600 28200
rect 128500 28200 128600 28300
rect 128500 28300 128600 28400
rect 128500 28400 128600 28500
rect 128500 28500 128600 28600
rect 128500 28600 128600 28700
rect 128500 28700 128600 28800
rect 128500 28800 128600 28900
rect 128500 28900 128600 29000
rect 128500 29000 128600 29100
rect 128500 29100 128600 29200
rect 128500 29200 128600 29300
rect 128500 29300 128600 29400
rect 128500 29400 128600 29500
rect 128500 29500 128600 29600
rect 128500 29600 128600 29700
rect 128500 29700 128600 29800
rect 128500 29800 128600 29900
rect 128500 29900 128600 30000
rect 128500 30000 128600 30100
rect 128500 30100 128600 30200
rect 128500 30200 128600 30300
rect 128500 30300 128600 30400
rect 128500 30400 128600 30500
rect 128500 30500 128600 30600
rect 128500 30600 128600 30700
rect 128500 30700 128600 30800
rect 128500 30800 128600 30900
rect 128500 30900 128600 31000
rect 128500 31000 128600 31100
rect 128500 31100 128600 31200
rect 128500 31200 128600 31300
rect 128500 31300 128600 31400
rect 128500 31400 128600 31500
rect 128500 31500 128600 31600
rect 128500 31600 128600 31700
rect 128500 31700 128600 31800
rect 128500 31800 128600 31900
rect 128500 31900 128600 32000
rect 128500 32000 128600 32100
rect 128500 32100 128600 32200
rect 128500 32200 128600 32300
rect 128500 32300 128600 32400
rect 128500 32400 128600 32500
rect 128500 32500 128600 32600
rect 128500 32600 128600 32700
rect 128500 32700 128600 32800
rect 128500 32800 128600 32900
rect 128500 32900 128600 33000
rect 128500 36500 128600 36600
rect 128500 36600 128600 36700
rect 128500 36700 128600 36800
rect 128500 36800 128600 36900
rect 128500 36900 128600 37000
rect 128500 37000 128600 37100
rect 128500 37100 128600 37200
rect 128500 37200 128600 37300
rect 128500 37300 128600 37400
rect 128500 37400 128600 37500
rect 128500 37500 128600 37600
rect 128500 37600 128600 37700
rect 128600 24000 128700 24100
rect 128600 24100 128700 24200
rect 128600 24200 128700 24300
rect 128600 24300 128700 24400
rect 128600 24400 128700 24500
rect 128600 24500 128700 24600
rect 128600 28200 128700 28300
rect 128600 28300 128700 28400
rect 128600 28400 128700 28500
rect 128600 28500 128700 28600
rect 128600 28600 128700 28700
rect 128600 28700 128700 28800
rect 128600 28800 128700 28900
rect 128600 28900 128700 29000
rect 128600 29000 128700 29100
rect 128600 29100 128700 29200
rect 128600 29200 128700 29300
rect 128600 29300 128700 29400
rect 128600 29400 128700 29500
rect 128600 29500 128700 29600
rect 128600 29600 128700 29700
rect 128600 29700 128700 29800
rect 128600 29800 128700 29900
rect 128600 29900 128700 30000
rect 128600 30000 128700 30100
rect 128600 30100 128700 30200
rect 128600 30200 128700 30300
rect 128600 30300 128700 30400
rect 128600 30400 128700 30500
rect 128600 30500 128700 30600
rect 128600 30600 128700 30700
rect 128600 30700 128700 30800
rect 128600 30800 128700 30900
rect 128600 30900 128700 31000
rect 128600 31000 128700 31100
rect 128600 31100 128700 31200
rect 128600 31200 128700 31300
rect 128600 31300 128700 31400
rect 128600 31400 128700 31500
rect 128600 31500 128700 31600
rect 128600 31600 128700 31700
rect 128600 31700 128700 31800
rect 128600 31800 128700 31900
rect 128600 31900 128700 32000
rect 128600 32000 128700 32100
rect 128600 32100 128700 32200
rect 128600 32200 128700 32300
rect 128600 32300 128700 32400
rect 128600 32400 128700 32500
rect 128600 32500 128700 32600
rect 128600 32600 128700 32700
rect 128600 32700 128700 32800
rect 128600 32800 128700 32900
rect 128600 32900 128700 33000
rect 128600 33000 128700 33100
rect 128600 33100 128700 33200
rect 128600 33200 128700 33300
rect 128600 33300 128700 33400
rect 128600 36200 128700 36300
rect 128600 36300 128700 36400
rect 128600 36400 128700 36500
rect 128600 36500 128700 36600
rect 128600 36600 128700 36700
rect 128600 36700 128700 36800
rect 128600 36800 128700 36900
rect 128600 36900 128700 37000
rect 128600 37000 128700 37100
rect 128600 37100 128700 37200
rect 128600 37200 128700 37300
rect 128600 37300 128700 37400
rect 128600 37400 128700 37500
rect 128600 37500 128700 37600
rect 128600 37600 128700 37700
rect 128600 37700 128700 37800
rect 128600 37800 128700 37900
rect 128600 37900 128700 38000
rect 128700 28500 128800 28600
rect 128700 28600 128800 28700
rect 128700 28700 128800 28800
rect 128700 28800 128800 28900
rect 128700 28900 128800 29000
rect 128700 29000 128800 29100
rect 128700 29100 128800 29200
rect 128700 29200 128800 29300
rect 128700 29300 128800 29400
rect 128700 29400 128800 29500
rect 128700 29500 128800 29600
rect 128700 29600 128800 29700
rect 128700 29700 128800 29800
rect 128700 29800 128800 29900
rect 128700 29900 128800 30000
rect 128700 30000 128800 30100
rect 128700 30100 128800 30200
rect 128700 30200 128800 30300
rect 128700 30300 128800 30400
rect 128700 30400 128800 30500
rect 128700 30500 128800 30600
rect 128700 30600 128800 30700
rect 128700 30700 128800 30800
rect 128700 30800 128800 30900
rect 128700 30900 128800 31000
rect 128700 31000 128800 31100
rect 128700 31100 128800 31200
rect 128700 31200 128800 31300
rect 128700 31300 128800 31400
rect 128700 31400 128800 31500
rect 128700 31500 128800 31600
rect 128700 31600 128800 31700
rect 128700 31700 128800 31800
rect 128700 31800 128800 31900
rect 128700 31900 128800 32000
rect 128700 32000 128800 32100
rect 128700 32100 128800 32200
rect 128700 32200 128800 32300
rect 128700 32300 128800 32400
rect 128700 32400 128800 32500
rect 128700 32500 128800 32600
rect 128700 32600 128800 32700
rect 128700 32700 128800 32800
rect 128700 32800 128800 32900
rect 128700 32900 128800 33000
rect 128700 33000 128800 33100
rect 128700 33100 128800 33200
rect 128700 33200 128800 33300
rect 128700 33300 128800 33400
rect 128700 33400 128800 33500
rect 128700 33500 128800 33600
rect 128700 33600 128800 33700
rect 128700 35900 128800 36000
rect 128700 36000 128800 36100
rect 128700 36100 128800 36200
rect 128700 36200 128800 36300
rect 128700 36300 128800 36400
rect 128700 36400 128800 36500
rect 128700 36500 128800 36600
rect 128700 36600 128800 36700
rect 128700 36700 128800 36800
rect 128700 36800 128800 36900
rect 128700 36900 128800 37000
rect 128700 37000 128800 37100
rect 128700 37100 128800 37200
rect 128700 37200 128800 37300
rect 128700 37300 128800 37400
rect 128700 37400 128800 37500
rect 128700 37500 128800 37600
rect 128700 37600 128800 37700
rect 128700 37700 128800 37800
rect 128700 37800 128800 37900
rect 128700 37900 128800 38000
rect 128700 38000 128800 38100
rect 128700 38100 128800 38200
rect 128800 28700 128900 28800
rect 128800 28800 128900 28900
rect 128800 28900 128900 29000
rect 128800 29000 128900 29100
rect 128800 29100 128900 29200
rect 128800 29200 128900 29300
rect 128800 29300 128900 29400
rect 128800 29400 128900 29500
rect 128800 29500 128900 29600
rect 128800 29600 128900 29700
rect 128800 29700 128900 29800
rect 128800 29800 128900 29900
rect 128800 29900 128900 30000
rect 128800 30000 128900 30100
rect 128800 30100 128900 30200
rect 128800 30200 128900 30300
rect 128800 30300 128900 30400
rect 128800 30400 128900 30500
rect 128800 30500 128900 30600
rect 128800 30600 128900 30700
rect 128800 30700 128900 30800
rect 128800 30800 128900 30900
rect 128800 30900 128900 31000
rect 128800 31000 128900 31100
rect 128800 31100 128900 31200
rect 128800 31200 128900 31300
rect 128800 31300 128900 31400
rect 128800 31400 128900 31500
rect 128800 31500 128900 31600
rect 128800 31600 128900 31700
rect 128800 31700 128900 31800
rect 128800 31800 128900 31900
rect 128800 31900 128900 32000
rect 128800 32000 128900 32100
rect 128800 32100 128900 32200
rect 128800 32200 128900 32300
rect 128800 32300 128900 32400
rect 128800 32400 128900 32500
rect 128800 32500 128900 32600
rect 128800 32600 128900 32700
rect 128800 32700 128900 32800
rect 128800 32800 128900 32900
rect 128800 32900 128900 33000
rect 128800 33000 128900 33100
rect 128800 33100 128900 33200
rect 128800 33200 128900 33300
rect 128800 33300 128900 33400
rect 128800 33400 128900 33500
rect 128800 33500 128900 33600
rect 128800 33600 128900 33700
rect 128800 33700 128900 33800
rect 128800 33800 128900 33900
rect 128800 33900 128900 34000
rect 128800 34000 128900 34100
rect 128800 35700 128900 35800
rect 128800 35800 128900 35900
rect 128800 35900 128900 36000
rect 128800 36000 128900 36100
rect 128800 36100 128900 36200
rect 128800 36200 128900 36300
rect 128800 36300 128900 36400
rect 128800 36400 128900 36500
rect 128800 36500 128900 36600
rect 128800 36600 128900 36700
rect 128800 36700 128900 36800
rect 128800 36800 128900 36900
rect 128800 36900 128900 37000
rect 128800 37000 128900 37100
rect 128800 37100 128900 37200
rect 128800 37200 128900 37300
rect 128800 37300 128900 37400
rect 128800 37400 128900 37500
rect 128800 37500 128900 37600
rect 128800 37600 128900 37700
rect 128800 37700 128900 37800
rect 128800 37800 128900 37900
rect 128800 37900 128900 38000
rect 128800 38000 128900 38100
rect 128800 38100 128900 38200
rect 128800 38200 128900 38300
rect 128800 38300 128900 38400
rect 128900 29000 129000 29100
rect 128900 29100 129000 29200
rect 128900 29200 129000 29300
rect 128900 29300 129000 29400
rect 128900 29400 129000 29500
rect 128900 29500 129000 29600
rect 128900 29600 129000 29700
rect 128900 29700 129000 29800
rect 128900 29800 129000 29900
rect 128900 29900 129000 30000
rect 128900 30000 129000 30100
rect 128900 30100 129000 30200
rect 128900 30200 129000 30300
rect 128900 30300 129000 30400
rect 128900 30400 129000 30500
rect 128900 30500 129000 30600
rect 128900 30600 129000 30700
rect 128900 30700 129000 30800
rect 128900 30800 129000 30900
rect 128900 30900 129000 31000
rect 128900 31000 129000 31100
rect 128900 31100 129000 31200
rect 128900 31200 129000 31300
rect 128900 31300 129000 31400
rect 128900 31400 129000 31500
rect 128900 31500 129000 31600
rect 128900 31600 129000 31700
rect 128900 31700 129000 31800
rect 128900 31800 129000 31900
rect 128900 31900 129000 32000
rect 128900 32000 129000 32100
rect 128900 32100 129000 32200
rect 128900 32200 129000 32300
rect 128900 32300 129000 32400
rect 128900 32400 129000 32500
rect 128900 32500 129000 32600
rect 128900 32600 129000 32700
rect 128900 32700 129000 32800
rect 128900 32800 129000 32900
rect 128900 32900 129000 33000
rect 128900 33000 129000 33100
rect 128900 33100 129000 33200
rect 128900 33200 129000 33300
rect 128900 33300 129000 33400
rect 128900 33400 129000 33500
rect 128900 33500 129000 33600
rect 128900 33600 129000 33700
rect 128900 33700 129000 33800
rect 128900 33800 129000 33900
rect 128900 33900 129000 34000
rect 128900 34000 129000 34100
rect 128900 34100 129000 34200
rect 128900 34200 129000 34300
rect 128900 34300 129000 34400
rect 128900 34400 129000 34500
rect 128900 35400 129000 35500
rect 128900 35500 129000 35600
rect 128900 35600 129000 35700
rect 128900 35700 129000 35800
rect 128900 35800 129000 35900
rect 128900 35900 129000 36000
rect 128900 36000 129000 36100
rect 128900 36100 129000 36200
rect 128900 36200 129000 36300
rect 128900 36300 129000 36400
rect 128900 36400 129000 36500
rect 128900 36500 129000 36600
rect 128900 36600 129000 36700
rect 128900 36700 129000 36800
rect 128900 36800 129000 36900
rect 128900 36900 129000 37000
rect 128900 37000 129000 37100
rect 128900 37100 129000 37200
rect 128900 37200 129000 37300
rect 128900 37300 129000 37400
rect 128900 37400 129000 37500
rect 128900 37500 129000 37600
rect 128900 37600 129000 37700
rect 128900 37700 129000 37800
rect 128900 37800 129000 37900
rect 128900 37900 129000 38000
rect 128900 38000 129000 38100
rect 128900 38100 129000 38200
rect 128900 38200 129000 38300
rect 128900 38300 129000 38400
rect 128900 38400 129000 38500
rect 129000 29300 129100 29400
rect 129000 29400 129100 29500
rect 129000 29500 129100 29600
rect 129000 29600 129100 29700
rect 129000 29700 129100 29800
rect 129000 29800 129100 29900
rect 129000 29900 129100 30000
rect 129000 30000 129100 30100
rect 129000 30100 129100 30200
rect 129000 30200 129100 30300
rect 129000 30300 129100 30400
rect 129000 30400 129100 30500
rect 129000 30500 129100 30600
rect 129000 30600 129100 30700
rect 129000 30700 129100 30800
rect 129000 30800 129100 30900
rect 129000 30900 129100 31000
rect 129000 31000 129100 31100
rect 129000 31100 129100 31200
rect 129000 31200 129100 31300
rect 129000 31300 129100 31400
rect 129000 31400 129100 31500
rect 129000 31500 129100 31600
rect 129000 31600 129100 31700
rect 129000 31700 129100 31800
rect 129000 31800 129100 31900
rect 129000 31900 129100 32000
rect 129000 32000 129100 32100
rect 129000 32100 129100 32200
rect 129000 32200 129100 32300
rect 129000 32300 129100 32400
rect 129000 32400 129100 32500
rect 129000 32500 129100 32600
rect 129000 32600 129100 32700
rect 129000 32700 129100 32800
rect 129000 32800 129100 32900
rect 129000 32900 129100 33000
rect 129000 33000 129100 33100
rect 129000 33100 129100 33200
rect 129000 33200 129100 33300
rect 129000 33300 129100 33400
rect 129000 33400 129100 33500
rect 129000 33500 129100 33600
rect 129000 33600 129100 33700
rect 129000 33700 129100 33800
rect 129000 33800 129100 33900
rect 129000 33900 129100 34000
rect 129000 34000 129100 34100
rect 129000 34100 129100 34200
rect 129000 34200 129100 34300
rect 129000 34300 129100 34400
rect 129000 34400 129100 34500
rect 129000 34500 129100 34600
rect 129000 34600 129100 34700
rect 129000 34700 129100 34800
rect 129000 34800 129100 34900
rect 129000 34900 129100 35000
rect 129000 35000 129100 35100
rect 129000 35100 129100 35200
rect 129000 35200 129100 35300
rect 129000 35300 129100 35400
rect 129000 35400 129100 35500
rect 129000 35500 129100 35600
rect 129000 35600 129100 35700
rect 129000 35700 129100 35800
rect 129000 35800 129100 35900
rect 129000 35900 129100 36000
rect 129000 36000 129100 36100
rect 129000 36100 129100 36200
rect 129000 36200 129100 36300
rect 129000 36300 129100 36400
rect 129000 36400 129100 36500
rect 129000 36500 129100 36600
rect 129000 36600 129100 36700
rect 129000 36700 129100 36800
rect 129000 36800 129100 36900
rect 129000 36900 129100 37000
rect 129000 37000 129100 37100
rect 129000 37100 129100 37200
rect 129000 37200 129100 37300
rect 129000 37300 129100 37400
rect 129000 37400 129100 37500
rect 129000 37500 129100 37600
rect 129000 37600 129100 37700
rect 129000 37700 129100 37800
rect 129000 37800 129100 37900
rect 129000 37900 129100 38000
rect 129000 38000 129100 38100
rect 129000 38100 129100 38200
rect 129000 38200 129100 38300
rect 129000 38300 129100 38400
rect 129000 38400 129100 38500
rect 129000 38500 129100 38600
rect 129000 38600 129100 38700
rect 129100 29600 129200 29700
rect 129100 29700 129200 29800
rect 129100 29800 129200 29900
rect 129100 29900 129200 30000
rect 129100 30000 129200 30100
rect 129100 30100 129200 30200
rect 129100 30200 129200 30300
rect 129100 30300 129200 30400
rect 129100 30400 129200 30500
rect 129100 30500 129200 30600
rect 129100 30600 129200 30700
rect 129100 30700 129200 30800
rect 129100 30800 129200 30900
rect 129100 30900 129200 31000
rect 129100 31000 129200 31100
rect 129100 31100 129200 31200
rect 129100 31200 129200 31300
rect 129100 31300 129200 31400
rect 129100 31400 129200 31500
rect 129100 31500 129200 31600
rect 129100 31600 129200 31700
rect 129100 31700 129200 31800
rect 129100 31800 129200 31900
rect 129100 31900 129200 32000
rect 129100 32000 129200 32100
rect 129100 32100 129200 32200
rect 129100 32200 129200 32300
rect 129100 32300 129200 32400
rect 129100 32400 129200 32500
rect 129100 32500 129200 32600
rect 129100 32600 129200 32700
rect 129100 32700 129200 32800
rect 129100 32800 129200 32900
rect 129100 32900 129200 33000
rect 129100 33000 129200 33100
rect 129100 33100 129200 33200
rect 129100 33200 129200 33300
rect 129100 33300 129200 33400
rect 129100 33400 129200 33500
rect 129100 33500 129200 33600
rect 129100 33600 129200 33700
rect 129100 33700 129200 33800
rect 129100 33800 129200 33900
rect 129100 33900 129200 34000
rect 129100 34000 129200 34100
rect 129100 34100 129200 34200
rect 129100 34200 129200 34300
rect 129100 34300 129200 34400
rect 129100 34400 129200 34500
rect 129100 34500 129200 34600
rect 129100 34600 129200 34700
rect 129100 34700 129200 34800
rect 129100 34800 129200 34900
rect 129100 34900 129200 35000
rect 129100 35000 129200 35100
rect 129100 35100 129200 35200
rect 129100 35200 129200 35300
rect 129100 35300 129200 35400
rect 129100 35400 129200 35500
rect 129100 35500 129200 35600
rect 129100 35600 129200 35700
rect 129100 35700 129200 35800
rect 129100 35800 129200 35900
rect 129100 35900 129200 36000
rect 129100 36000 129200 36100
rect 129100 36100 129200 36200
rect 129100 36200 129200 36300
rect 129100 36300 129200 36400
rect 129100 36400 129200 36500
rect 129100 36500 129200 36600
rect 129100 36600 129200 36700
rect 129100 36700 129200 36800
rect 129100 36800 129200 36900
rect 129100 36900 129200 37000
rect 129100 37000 129200 37100
rect 129100 37100 129200 37200
rect 129100 37200 129200 37300
rect 129100 37300 129200 37400
rect 129100 37400 129200 37500
rect 129100 37500 129200 37600
rect 129100 37600 129200 37700
rect 129100 37700 129200 37800
rect 129100 37800 129200 37900
rect 129100 37900 129200 38000
rect 129100 38000 129200 38100
rect 129100 38100 129200 38200
rect 129100 38200 129200 38300
rect 129100 38300 129200 38400
rect 129100 38400 129200 38500
rect 129100 38500 129200 38600
rect 129100 38600 129200 38700
rect 129100 38700 129200 38800
rect 129200 29900 129300 30000
rect 129200 30000 129300 30100
rect 129200 30100 129300 30200
rect 129200 30200 129300 30300
rect 129200 30300 129300 30400
rect 129200 30400 129300 30500
rect 129200 30500 129300 30600
rect 129200 30600 129300 30700
rect 129200 30700 129300 30800
rect 129200 30800 129300 30900
rect 129200 30900 129300 31000
rect 129200 31000 129300 31100
rect 129200 31100 129300 31200
rect 129200 31200 129300 31300
rect 129200 31300 129300 31400
rect 129200 31400 129300 31500
rect 129200 31500 129300 31600
rect 129200 31600 129300 31700
rect 129200 31700 129300 31800
rect 129200 31800 129300 31900
rect 129200 31900 129300 32000
rect 129200 32000 129300 32100
rect 129200 32100 129300 32200
rect 129200 32200 129300 32300
rect 129200 32300 129300 32400
rect 129200 32400 129300 32500
rect 129200 32500 129300 32600
rect 129200 32600 129300 32700
rect 129200 32700 129300 32800
rect 129200 32800 129300 32900
rect 129200 32900 129300 33000
rect 129200 33000 129300 33100
rect 129200 33100 129300 33200
rect 129200 33200 129300 33300
rect 129200 33300 129300 33400
rect 129200 33400 129300 33500
rect 129200 33500 129300 33600
rect 129200 33600 129300 33700
rect 129200 33700 129300 33800
rect 129200 33800 129300 33900
rect 129200 33900 129300 34000
rect 129200 34000 129300 34100
rect 129200 34100 129300 34200
rect 129200 34200 129300 34300
rect 129200 34300 129300 34400
rect 129200 34400 129300 34500
rect 129200 34500 129300 34600
rect 129200 34600 129300 34700
rect 129200 34700 129300 34800
rect 129200 34800 129300 34900
rect 129200 34900 129300 35000
rect 129200 35000 129300 35100
rect 129200 35100 129300 35200
rect 129200 35200 129300 35300
rect 129200 35300 129300 35400
rect 129200 35400 129300 35500
rect 129200 35500 129300 35600
rect 129200 35600 129300 35700
rect 129200 35700 129300 35800
rect 129200 35800 129300 35900
rect 129200 35900 129300 36000
rect 129200 36000 129300 36100
rect 129200 36100 129300 36200
rect 129200 36200 129300 36300
rect 129200 36300 129300 36400
rect 129200 36400 129300 36500
rect 129200 36500 129300 36600
rect 129200 36600 129300 36700
rect 129200 36700 129300 36800
rect 129200 36800 129300 36900
rect 129200 36900 129300 37000
rect 129200 37000 129300 37100
rect 129200 37100 129300 37200
rect 129200 37200 129300 37300
rect 129200 37300 129300 37400
rect 129200 37400 129300 37500
rect 129200 37500 129300 37600
rect 129200 37600 129300 37700
rect 129200 37700 129300 37800
rect 129200 37800 129300 37900
rect 129200 37900 129300 38000
rect 129200 38000 129300 38100
rect 129200 38100 129300 38200
rect 129200 38200 129300 38300
rect 129200 38300 129300 38400
rect 129200 38400 129300 38500
rect 129200 38500 129300 38600
rect 129200 38600 129300 38700
rect 129200 38700 129300 38800
rect 129200 38800 129300 38900
rect 129300 30100 129400 30200
rect 129300 30200 129400 30300
rect 129300 30300 129400 30400
rect 129300 30400 129400 30500
rect 129300 30500 129400 30600
rect 129300 30600 129400 30700
rect 129300 30700 129400 30800
rect 129300 30800 129400 30900
rect 129300 30900 129400 31000
rect 129300 31000 129400 31100
rect 129300 31100 129400 31200
rect 129300 31200 129400 31300
rect 129300 31300 129400 31400
rect 129300 31400 129400 31500
rect 129300 31500 129400 31600
rect 129300 31600 129400 31700
rect 129300 31700 129400 31800
rect 129300 31800 129400 31900
rect 129300 31900 129400 32000
rect 129300 32000 129400 32100
rect 129300 32100 129400 32200
rect 129300 32200 129400 32300
rect 129300 32300 129400 32400
rect 129300 32400 129400 32500
rect 129300 32500 129400 32600
rect 129300 32600 129400 32700
rect 129300 32700 129400 32800
rect 129300 32800 129400 32900
rect 129300 32900 129400 33000
rect 129300 33000 129400 33100
rect 129300 33100 129400 33200
rect 129300 33200 129400 33300
rect 129300 33300 129400 33400
rect 129300 33400 129400 33500
rect 129300 33500 129400 33600
rect 129300 33600 129400 33700
rect 129300 33700 129400 33800
rect 129300 33800 129400 33900
rect 129300 33900 129400 34000
rect 129300 34000 129400 34100
rect 129300 34100 129400 34200
rect 129300 34200 129400 34300
rect 129300 34300 129400 34400
rect 129300 34400 129400 34500
rect 129300 34500 129400 34600
rect 129300 34600 129400 34700
rect 129300 34700 129400 34800
rect 129300 34800 129400 34900
rect 129300 34900 129400 35000
rect 129300 35000 129400 35100
rect 129300 35100 129400 35200
rect 129300 35200 129400 35300
rect 129300 35300 129400 35400
rect 129300 35400 129400 35500
rect 129300 35500 129400 35600
rect 129300 35600 129400 35700
rect 129300 35700 129400 35800
rect 129300 35800 129400 35900
rect 129300 35900 129400 36000
rect 129300 36000 129400 36100
rect 129300 36100 129400 36200
rect 129300 36200 129400 36300
rect 129300 36300 129400 36400
rect 129300 36400 129400 36500
rect 129300 36500 129400 36600
rect 129300 36600 129400 36700
rect 129300 36700 129400 36800
rect 129300 36800 129400 36900
rect 129300 36900 129400 37000
rect 129300 37000 129400 37100
rect 129300 37100 129400 37200
rect 129300 37200 129400 37300
rect 129300 37300 129400 37400
rect 129300 37400 129400 37500
rect 129300 37500 129400 37600
rect 129300 37600 129400 37700
rect 129300 37700 129400 37800
rect 129300 37800 129400 37900
rect 129300 37900 129400 38000
rect 129300 38000 129400 38100
rect 129300 38100 129400 38200
rect 129300 38200 129400 38300
rect 129300 38300 129400 38400
rect 129300 38400 129400 38500
rect 129300 38500 129400 38600
rect 129300 38600 129400 38700
rect 129300 38700 129400 38800
rect 129300 38800 129400 38900
rect 129300 38900 129400 39000
rect 129400 30400 129500 30500
rect 129400 30500 129500 30600
rect 129400 30600 129500 30700
rect 129400 30700 129500 30800
rect 129400 30800 129500 30900
rect 129400 30900 129500 31000
rect 129400 31000 129500 31100
rect 129400 31100 129500 31200
rect 129400 31200 129500 31300
rect 129400 31300 129500 31400
rect 129400 31400 129500 31500
rect 129400 31500 129500 31600
rect 129400 31600 129500 31700
rect 129400 31700 129500 31800
rect 129400 31800 129500 31900
rect 129400 31900 129500 32000
rect 129400 32000 129500 32100
rect 129400 32100 129500 32200
rect 129400 32200 129500 32300
rect 129400 32300 129500 32400
rect 129400 32400 129500 32500
rect 129400 32500 129500 32600
rect 129400 32600 129500 32700
rect 129400 32700 129500 32800
rect 129400 32800 129500 32900
rect 129400 32900 129500 33000
rect 129400 33000 129500 33100
rect 129400 33100 129500 33200
rect 129400 33200 129500 33300
rect 129400 33300 129500 33400
rect 129400 33400 129500 33500
rect 129400 33500 129500 33600
rect 129400 33600 129500 33700
rect 129400 33700 129500 33800
rect 129400 33800 129500 33900
rect 129400 33900 129500 34000
rect 129400 34000 129500 34100
rect 129400 34100 129500 34200
rect 129400 34200 129500 34300
rect 129400 34300 129500 34400
rect 129400 34400 129500 34500
rect 129400 34500 129500 34600
rect 129400 34600 129500 34700
rect 129400 34700 129500 34800
rect 129400 34800 129500 34900
rect 129400 34900 129500 35000
rect 129400 35000 129500 35100
rect 129400 35100 129500 35200
rect 129400 35200 129500 35300
rect 129400 35300 129500 35400
rect 129400 35400 129500 35500
rect 129400 35500 129500 35600
rect 129400 35600 129500 35700
rect 129400 35700 129500 35800
rect 129400 35800 129500 35900
rect 129400 35900 129500 36000
rect 129400 36000 129500 36100
rect 129400 36100 129500 36200
rect 129400 36200 129500 36300
rect 129400 36300 129500 36400
rect 129400 36400 129500 36500
rect 129400 36500 129500 36600
rect 129400 36600 129500 36700
rect 129400 36700 129500 36800
rect 129400 36800 129500 36900
rect 129400 36900 129500 37000
rect 129400 37000 129500 37100
rect 129400 37100 129500 37200
rect 129400 37200 129500 37300
rect 129400 37300 129500 37400
rect 129400 37400 129500 37500
rect 129400 37500 129500 37600
rect 129400 37600 129500 37700
rect 129400 37700 129500 37800
rect 129400 37800 129500 37900
rect 129400 37900 129500 38000
rect 129400 38000 129500 38100
rect 129400 38100 129500 38200
rect 129400 38200 129500 38300
rect 129400 38300 129500 38400
rect 129400 38400 129500 38500
rect 129400 38500 129500 38600
rect 129400 38600 129500 38700
rect 129400 38700 129500 38800
rect 129400 38800 129500 38900
rect 129400 38900 129500 39000
rect 129500 30700 129600 30800
rect 129500 30800 129600 30900
rect 129500 30900 129600 31000
rect 129500 31000 129600 31100
rect 129500 31100 129600 31200
rect 129500 31200 129600 31300
rect 129500 31300 129600 31400
rect 129500 31400 129600 31500
rect 129500 31500 129600 31600
rect 129500 31600 129600 31700
rect 129500 31700 129600 31800
rect 129500 31800 129600 31900
rect 129500 31900 129600 32000
rect 129500 32000 129600 32100
rect 129500 32100 129600 32200
rect 129500 32200 129600 32300
rect 129500 32300 129600 32400
rect 129500 32400 129600 32500
rect 129500 32500 129600 32600
rect 129500 32600 129600 32700
rect 129500 32700 129600 32800
rect 129500 32800 129600 32900
rect 129500 32900 129600 33000
rect 129500 33000 129600 33100
rect 129500 33100 129600 33200
rect 129500 33200 129600 33300
rect 129500 33300 129600 33400
rect 129500 33400 129600 33500
rect 129500 33500 129600 33600
rect 129500 33600 129600 33700
rect 129500 33700 129600 33800
rect 129500 33800 129600 33900
rect 129500 33900 129600 34000
rect 129500 34000 129600 34100
rect 129500 34100 129600 34200
rect 129500 34200 129600 34300
rect 129500 34300 129600 34400
rect 129500 34400 129600 34500
rect 129500 34500 129600 34600
rect 129500 34600 129600 34700
rect 129500 34700 129600 34800
rect 129500 34800 129600 34900
rect 129500 34900 129600 35000
rect 129500 35000 129600 35100
rect 129500 35100 129600 35200
rect 129500 35200 129600 35300
rect 129500 35300 129600 35400
rect 129500 35400 129600 35500
rect 129500 35500 129600 35600
rect 129500 35600 129600 35700
rect 129500 35700 129600 35800
rect 129500 35800 129600 35900
rect 129500 35900 129600 36000
rect 129500 36000 129600 36100
rect 129500 36100 129600 36200
rect 129500 36200 129600 36300
rect 129500 36300 129600 36400
rect 129500 36400 129600 36500
rect 129500 36500 129600 36600
rect 129500 36600 129600 36700
rect 129500 36700 129600 36800
rect 129500 36800 129600 36900
rect 129500 36900 129600 37000
rect 129500 37000 129600 37100
rect 129500 37100 129600 37200
rect 129500 37200 129600 37300
rect 129500 37300 129600 37400
rect 129500 37400 129600 37500
rect 129500 37500 129600 37600
rect 129500 37600 129600 37700
rect 129500 37700 129600 37800
rect 129500 37800 129600 37900
rect 129500 37900 129600 38000
rect 129500 38000 129600 38100
rect 129500 38100 129600 38200
rect 129500 38200 129600 38300
rect 129500 38300 129600 38400
rect 129500 38400 129600 38500
rect 129500 38500 129600 38600
rect 129500 38600 129600 38700
rect 129500 38700 129600 38800
rect 129500 38800 129600 38900
rect 129500 38900 129600 39000
rect 129500 39000 129600 39100
rect 129600 30900 129700 31000
rect 129600 31000 129700 31100
rect 129600 31100 129700 31200
rect 129600 31200 129700 31300
rect 129600 31300 129700 31400
rect 129600 31400 129700 31500
rect 129600 31500 129700 31600
rect 129600 31600 129700 31700
rect 129600 31700 129700 31800
rect 129600 31800 129700 31900
rect 129600 31900 129700 32000
rect 129600 32000 129700 32100
rect 129600 32100 129700 32200
rect 129600 32200 129700 32300
rect 129600 32300 129700 32400
rect 129600 32400 129700 32500
rect 129600 32500 129700 32600
rect 129600 32600 129700 32700
rect 129600 32700 129700 32800
rect 129600 32800 129700 32900
rect 129600 32900 129700 33000
rect 129600 33000 129700 33100
rect 129600 33100 129700 33200
rect 129600 33200 129700 33300
rect 129600 33300 129700 33400
rect 129600 33400 129700 33500
rect 129600 33500 129700 33600
rect 129600 33600 129700 33700
rect 129600 33700 129700 33800
rect 129600 33800 129700 33900
rect 129600 33900 129700 34000
rect 129600 34000 129700 34100
rect 129600 34100 129700 34200
rect 129600 34200 129700 34300
rect 129600 34300 129700 34400
rect 129600 34400 129700 34500
rect 129600 34500 129700 34600
rect 129600 34600 129700 34700
rect 129600 34700 129700 34800
rect 129600 34800 129700 34900
rect 129600 34900 129700 35000
rect 129600 35000 129700 35100
rect 129600 35100 129700 35200
rect 129600 35200 129700 35300
rect 129600 35300 129700 35400
rect 129600 35400 129700 35500
rect 129600 35500 129700 35600
rect 129600 35600 129700 35700
rect 129600 35700 129700 35800
rect 129600 35800 129700 35900
rect 129600 35900 129700 36000
rect 129600 36000 129700 36100
rect 129600 36100 129700 36200
rect 129600 36200 129700 36300
rect 129600 36300 129700 36400
rect 129600 36400 129700 36500
rect 129600 36500 129700 36600
rect 129600 36600 129700 36700
rect 129600 36700 129700 36800
rect 129600 36800 129700 36900
rect 129600 36900 129700 37000
rect 129600 37000 129700 37100
rect 129600 37100 129700 37200
rect 129600 37200 129700 37300
rect 129600 37300 129700 37400
rect 129600 37400 129700 37500
rect 129600 37500 129700 37600
rect 129600 37600 129700 37700
rect 129600 37700 129700 37800
rect 129600 37800 129700 37900
rect 129600 37900 129700 38000
rect 129600 38000 129700 38100
rect 129600 38100 129700 38200
rect 129600 38200 129700 38300
rect 129600 38300 129700 38400
rect 129600 38400 129700 38500
rect 129600 38500 129700 38600
rect 129600 38600 129700 38700
rect 129600 38700 129700 38800
rect 129600 38800 129700 38900
rect 129600 38900 129700 39000
rect 129600 39000 129700 39100
rect 129600 39100 129700 39200
rect 129700 31200 129800 31300
rect 129700 31300 129800 31400
rect 129700 31400 129800 31500
rect 129700 31500 129800 31600
rect 129700 31600 129800 31700
rect 129700 31700 129800 31800
rect 129700 31800 129800 31900
rect 129700 31900 129800 32000
rect 129700 32000 129800 32100
rect 129700 32100 129800 32200
rect 129700 32200 129800 32300
rect 129700 32300 129800 32400
rect 129700 32400 129800 32500
rect 129700 32500 129800 32600
rect 129700 32600 129800 32700
rect 129700 32700 129800 32800
rect 129700 32800 129800 32900
rect 129700 32900 129800 33000
rect 129700 33000 129800 33100
rect 129700 33100 129800 33200
rect 129700 33200 129800 33300
rect 129700 33300 129800 33400
rect 129700 33400 129800 33500
rect 129700 33500 129800 33600
rect 129700 33600 129800 33700
rect 129700 33700 129800 33800
rect 129700 33800 129800 33900
rect 129700 33900 129800 34000
rect 129700 34000 129800 34100
rect 129700 34100 129800 34200
rect 129700 34200 129800 34300
rect 129700 34300 129800 34400
rect 129700 34400 129800 34500
rect 129700 34500 129800 34600
rect 129700 34600 129800 34700
rect 129700 34700 129800 34800
rect 129700 34800 129800 34900
rect 129700 34900 129800 35000
rect 129700 35000 129800 35100
rect 129700 35100 129800 35200
rect 129700 35200 129800 35300
rect 129700 35300 129800 35400
rect 129700 35400 129800 35500
rect 129700 35500 129800 35600
rect 129700 35600 129800 35700
rect 129700 35700 129800 35800
rect 129700 35800 129800 35900
rect 129700 35900 129800 36000
rect 129700 36000 129800 36100
rect 129700 36100 129800 36200
rect 129700 36200 129800 36300
rect 129700 36300 129800 36400
rect 129700 36400 129800 36500
rect 129700 36500 129800 36600
rect 129700 36600 129800 36700
rect 129700 36700 129800 36800
rect 129700 36800 129800 36900
rect 129700 36900 129800 37000
rect 129700 37000 129800 37100
rect 129700 37100 129800 37200
rect 129700 37200 129800 37300
rect 129700 37300 129800 37400
rect 129700 37400 129800 37500
rect 129700 37500 129800 37600
rect 129700 37600 129800 37700
rect 129700 37700 129800 37800
rect 129700 37800 129800 37900
rect 129700 37900 129800 38000
rect 129700 38000 129800 38100
rect 129700 38100 129800 38200
rect 129700 38200 129800 38300
rect 129700 38300 129800 38400
rect 129700 38400 129800 38500
rect 129700 38500 129800 38600
rect 129700 38600 129800 38700
rect 129700 38700 129800 38800
rect 129700 38800 129800 38900
rect 129700 38900 129800 39000
rect 129700 39000 129800 39100
rect 129700 39100 129800 39200
rect 129800 31500 129900 31600
rect 129800 31600 129900 31700
rect 129800 31700 129900 31800
rect 129800 31800 129900 31900
rect 129800 31900 129900 32000
rect 129800 32000 129900 32100
rect 129800 32100 129900 32200
rect 129800 32200 129900 32300
rect 129800 32300 129900 32400
rect 129800 32400 129900 32500
rect 129800 32500 129900 32600
rect 129800 32600 129900 32700
rect 129800 32700 129900 32800
rect 129800 32800 129900 32900
rect 129800 32900 129900 33000
rect 129800 33000 129900 33100
rect 129800 33100 129900 33200
rect 129800 33200 129900 33300
rect 129800 33300 129900 33400
rect 129800 33400 129900 33500
rect 129800 33500 129900 33600
rect 129800 33600 129900 33700
rect 129800 33700 129900 33800
rect 129800 33800 129900 33900
rect 129800 33900 129900 34000
rect 129800 34000 129900 34100
rect 129800 34100 129900 34200
rect 129800 34200 129900 34300
rect 129800 34300 129900 34400
rect 129800 34400 129900 34500
rect 129800 34500 129900 34600
rect 129800 34600 129900 34700
rect 129800 34700 129900 34800
rect 129800 34800 129900 34900
rect 129800 34900 129900 35000
rect 129800 35000 129900 35100
rect 129800 35100 129900 35200
rect 129800 35200 129900 35300
rect 129800 35300 129900 35400
rect 129800 35400 129900 35500
rect 129800 35500 129900 35600
rect 129800 35600 129900 35700
rect 129800 35700 129900 35800
rect 129800 35800 129900 35900
rect 129800 35900 129900 36000
rect 129800 36000 129900 36100
rect 129800 36100 129900 36200
rect 129800 36200 129900 36300
rect 129800 36300 129900 36400
rect 129800 36400 129900 36500
rect 129800 36500 129900 36600
rect 129800 36600 129900 36700
rect 129800 36700 129900 36800
rect 129800 36800 129900 36900
rect 129800 36900 129900 37000
rect 129800 37000 129900 37100
rect 129800 37100 129900 37200
rect 129800 37200 129900 37300
rect 129800 37300 129900 37400
rect 129800 37400 129900 37500
rect 129800 37500 129900 37600
rect 129800 37600 129900 37700
rect 129800 37700 129900 37800
rect 129800 37800 129900 37900
rect 129800 37900 129900 38000
rect 129800 38000 129900 38100
rect 129800 38100 129900 38200
rect 129800 38200 129900 38300
rect 129800 38300 129900 38400
rect 129800 38400 129900 38500
rect 129800 38500 129900 38600
rect 129800 38600 129900 38700
rect 129800 38700 129900 38800
rect 129800 38800 129900 38900
rect 129800 38900 129900 39000
rect 129800 39000 129900 39100
rect 129800 39100 129900 39200
rect 129800 39200 129900 39300
rect 129900 31700 130000 31800
rect 129900 31800 130000 31900
rect 129900 31900 130000 32000
rect 129900 32000 130000 32100
rect 129900 32100 130000 32200
rect 129900 32200 130000 32300
rect 129900 32300 130000 32400
rect 129900 32400 130000 32500
rect 129900 32500 130000 32600
rect 129900 32600 130000 32700
rect 129900 32700 130000 32800
rect 129900 32800 130000 32900
rect 129900 32900 130000 33000
rect 129900 33000 130000 33100
rect 129900 33100 130000 33200
rect 129900 33200 130000 33300
rect 129900 33300 130000 33400
rect 129900 33400 130000 33500
rect 129900 33500 130000 33600
rect 129900 33600 130000 33700
rect 129900 33700 130000 33800
rect 129900 33800 130000 33900
rect 129900 33900 130000 34000
rect 129900 34000 130000 34100
rect 129900 34100 130000 34200
rect 129900 34200 130000 34300
rect 129900 34300 130000 34400
rect 129900 34400 130000 34500
rect 129900 34500 130000 34600
rect 129900 34600 130000 34700
rect 129900 34700 130000 34800
rect 129900 34800 130000 34900
rect 129900 34900 130000 35000
rect 129900 35000 130000 35100
rect 129900 35100 130000 35200
rect 129900 35200 130000 35300
rect 129900 35300 130000 35400
rect 129900 35400 130000 35500
rect 129900 35500 130000 35600
rect 129900 35600 130000 35700
rect 129900 35700 130000 35800
rect 129900 35800 130000 35900
rect 129900 35900 130000 36000
rect 129900 36000 130000 36100
rect 129900 36100 130000 36200
rect 129900 36200 130000 36300
rect 129900 36300 130000 36400
rect 129900 36400 130000 36500
rect 129900 36500 130000 36600
rect 129900 36600 130000 36700
rect 129900 36700 130000 36800
rect 129900 36800 130000 36900
rect 129900 36900 130000 37000
rect 129900 37000 130000 37100
rect 129900 37100 130000 37200
rect 129900 37200 130000 37300
rect 129900 37300 130000 37400
rect 129900 37400 130000 37500
rect 129900 37500 130000 37600
rect 129900 37600 130000 37700
rect 129900 37700 130000 37800
rect 129900 37800 130000 37900
rect 129900 37900 130000 38000
rect 129900 38000 130000 38100
rect 129900 38100 130000 38200
rect 129900 38200 130000 38300
rect 129900 38300 130000 38400
rect 129900 38400 130000 38500
rect 129900 38500 130000 38600
rect 129900 38600 130000 38700
rect 129900 38700 130000 38800
rect 129900 38800 130000 38900
rect 129900 38900 130000 39000
rect 129900 39000 130000 39100
rect 129900 39100 130000 39200
rect 129900 39200 130000 39300
rect 130000 32000 130100 32100
rect 130000 32100 130100 32200
rect 130000 32200 130100 32300
rect 130000 32300 130100 32400
rect 130000 32400 130100 32500
rect 130000 32500 130100 32600
rect 130000 32600 130100 32700
rect 130000 32700 130100 32800
rect 130000 32800 130100 32900
rect 130000 32900 130100 33000
rect 130000 33000 130100 33100
rect 130000 33100 130100 33200
rect 130000 33200 130100 33300
rect 130000 33300 130100 33400
rect 130000 33400 130100 33500
rect 130000 33500 130100 33600
rect 130000 33600 130100 33700
rect 130000 33700 130100 33800
rect 130000 33800 130100 33900
rect 130000 33900 130100 34000
rect 130000 34000 130100 34100
rect 130000 34100 130100 34200
rect 130000 34200 130100 34300
rect 130000 34300 130100 34400
rect 130000 34400 130100 34500
rect 130000 34500 130100 34600
rect 130000 34600 130100 34700
rect 130000 34700 130100 34800
rect 130000 34800 130100 34900
rect 130000 34900 130100 35000
rect 130000 35000 130100 35100
rect 130000 35100 130100 35200
rect 130000 35200 130100 35300
rect 130000 35300 130100 35400
rect 130000 35400 130100 35500
rect 130000 35500 130100 35600
rect 130000 35600 130100 35700
rect 130000 35700 130100 35800
rect 130000 35800 130100 35900
rect 130000 35900 130100 36000
rect 130000 36000 130100 36100
rect 130000 36100 130100 36200
rect 130000 36200 130100 36300
rect 130000 36300 130100 36400
rect 130000 36400 130100 36500
rect 130000 36500 130100 36600
rect 130000 36600 130100 36700
rect 130000 36700 130100 36800
rect 130000 36800 130100 36900
rect 130000 36900 130100 37000
rect 130000 37000 130100 37100
rect 130000 37100 130100 37200
rect 130000 37200 130100 37300
rect 130000 37300 130100 37400
rect 130000 37400 130100 37500
rect 130000 37500 130100 37600
rect 130000 37600 130100 37700
rect 130000 37700 130100 37800
rect 130000 37800 130100 37900
rect 130000 37900 130100 38000
rect 130000 38000 130100 38100
rect 130000 38100 130100 38200
rect 130000 38200 130100 38300
rect 130000 38300 130100 38400
rect 130000 38400 130100 38500
rect 130000 38500 130100 38600
rect 130000 38600 130100 38700
rect 130000 38700 130100 38800
rect 130000 38800 130100 38900
rect 130000 38900 130100 39000
rect 130000 39000 130100 39100
rect 130000 39100 130100 39200
rect 130000 39200 130100 39300
rect 130100 32200 130200 32300
rect 130100 32300 130200 32400
rect 130100 32400 130200 32500
rect 130100 32500 130200 32600
rect 130100 32600 130200 32700
rect 130100 32700 130200 32800
rect 130100 32800 130200 32900
rect 130100 32900 130200 33000
rect 130100 33000 130200 33100
rect 130100 33100 130200 33200
rect 130100 33200 130200 33300
rect 130100 33300 130200 33400
rect 130100 33400 130200 33500
rect 130100 33500 130200 33600
rect 130100 33600 130200 33700
rect 130100 33700 130200 33800
rect 130100 33800 130200 33900
rect 130100 33900 130200 34000
rect 130100 34000 130200 34100
rect 130100 34100 130200 34200
rect 130100 34200 130200 34300
rect 130100 34300 130200 34400
rect 130100 34400 130200 34500
rect 130100 34500 130200 34600
rect 130100 34600 130200 34700
rect 130100 34700 130200 34800
rect 130100 34800 130200 34900
rect 130100 34900 130200 35000
rect 130100 35000 130200 35100
rect 130100 35100 130200 35200
rect 130100 35200 130200 35300
rect 130100 35300 130200 35400
rect 130100 35400 130200 35500
rect 130100 35500 130200 35600
rect 130100 35600 130200 35700
rect 130100 35700 130200 35800
rect 130100 35800 130200 35900
rect 130100 35900 130200 36000
rect 130100 36000 130200 36100
rect 130100 36100 130200 36200
rect 130100 36200 130200 36300
rect 130100 36300 130200 36400
rect 130100 36400 130200 36500
rect 130100 36500 130200 36600
rect 130100 36600 130200 36700
rect 130100 37300 130200 37400
rect 130100 37400 130200 37500
rect 130100 37500 130200 37600
rect 130100 37600 130200 37700
rect 130100 37700 130200 37800
rect 130100 37800 130200 37900
rect 130100 37900 130200 38000
rect 130100 38000 130200 38100
rect 130100 38100 130200 38200
rect 130100 38200 130200 38300
rect 130100 38300 130200 38400
rect 130100 38400 130200 38500
rect 130100 38500 130200 38600
rect 130100 38600 130200 38700
rect 130100 38700 130200 38800
rect 130100 38800 130200 38900
rect 130100 38900 130200 39000
rect 130100 39000 130200 39100
rect 130100 39100 130200 39200
rect 130100 39200 130200 39300
rect 130100 39300 130200 39400
rect 130200 32500 130300 32600
rect 130200 32600 130300 32700
rect 130200 32700 130300 32800
rect 130200 32800 130300 32900
rect 130200 32900 130300 33000
rect 130200 33000 130300 33100
rect 130200 33100 130300 33200
rect 130200 33200 130300 33300
rect 130200 33300 130300 33400
rect 130200 33400 130300 33500
rect 130200 33500 130300 33600
rect 130200 33600 130300 33700
rect 130200 33700 130300 33800
rect 130200 33800 130300 33900
rect 130200 33900 130300 34000
rect 130200 34000 130300 34100
rect 130200 34100 130300 34200
rect 130200 34200 130300 34300
rect 130200 34300 130300 34400
rect 130200 34400 130300 34500
rect 130200 34500 130300 34600
rect 130200 34600 130300 34700
rect 130200 34700 130300 34800
rect 130200 34800 130300 34900
rect 130200 34900 130300 35000
rect 130200 35000 130300 35100
rect 130200 35100 130300 35200
rect 130200 35200 130300 35300
rect 130200 35300 130300 35400
rect 130200 35400 130300 35500
rect 130200 35500 130300 35600
rect 130200 35600 130300 35700
rect 130200 35700 130300 35800
rect 130200 35800 130300 35900
rect 130200 35900 130300 36000
rect 130200 36000 130300 36100
rect 130200 36100 130300 36200
rect 130200 36200 130300 36300
rect 130200 36300 130300 36400
rect 130200 36400 130300 36500
rect 130200 37400 130300 37500
rect 130200 37500 130300 37600
rect 130200 37600 130300 37700
rect 130200 37700 130300 37800
rect 130200 37800 130300 37900
rect 130200 37900 130300 38000
rect 130200 38000 130300 38100
rect 130200 38100 130300 38200
rect 130200 38200 130300 38300
rect 130200 38300 130300 38400
rect 130200 38400 130300 38500
rect 130200 38500 130300 38600
rect 130200 38600 130300 38700
rect 130200 38700 130300 38800
rect 130200 38800 130300 38900
rect 130200 38900 130300 39000
rect 130200 39000 130300 39100
rect 130200 39100 130300 39200
rect 130200 39200 130300 39300
rect 130200 39300 130300 39400
rect 130300 32700 130400 32800
rect 130300 32800 130400 32900
rect 130300 32900 130400 33000
rect 130300 33000 130400 33100
rect 130300 33100 130400 33200
rect 130300 33200 130400 33300
rect 130300 33300 130400 33400
rect 130300 33400 130400 33500
rect 130300 33500 130400 33600
rect 130300 33600 130400 33700
rect 130300 33700 130400 33800
rect 130300 33800 130400 33900
rect 130300 33900 130400 34000
rect 130300 34000 130400 34100
rect 130300 34100 130400 34200
rect 130300 34200 130400 34300
rect 130300 34300 130400 34400
rect 130300 34400 130400 34500
rect 130300 34500 130400 34600
rect 130300 34600 130400 34700
rect 130300 34700 130400 34800
rect 130300 34800 130400 34900
rect 130300 34900 130400 35000
rect 130300 35000 130400 35100
rect 130300 35100 130400 35200
rect 130300 35200 130400 35300
rect 130300 35300 130400 35400
rect 130300 35400 130400 35500
rect 130300 35500 130400 35600
rect 130300 35600 130400 35700
rect 130300 35700 130400 35800
rect 130300 35800 130400 35900
rect 130300 35900 130400 36000
rect 130300 36000 130400 36100
rect 130300 36100 130400 36200
rect 130300 36200 130400 36300
rect 130300 36300 130400 36400
rect 130300 37500 130400 37600
rect 130300 37600 130400 37700
rect 130300 37700 130400 37800
rect 130300 37800 130400 37900
rect 130300 37900 130400 38000
rect 130300 38000 130400 38100
rect 130300 38100 130400 38200
rect 130300 38200 130400 38300
rect 130300 38300 130400 38400
rect 130300 38400 130400 38500
rect 130300 38500 130400 38600
rect 130300 38600 130400 38700
rect 130300 38700 130400 38800
rect 130300 38800 130400 38900
rect 130300 38900 130400 39000
rect 130300 39000 130400 39100
rect 130300 39100 130400 39200
rect 130300 39200 130400 39300
rect 130300 39300 130400 39400
rect 130400 32900 130500 33000
rect 130400 33000 130500 33100
rect 130400 33100 130500 33200
rect 130400 33200 130500 33300
rect 130400 33300 130500 33400
rect 130400 33400 130500 33500
rect 130400 33500 130500 33600
rect 130400 33600 130500 33700
rect 130400 33700 130500 33800
rect 130400 33800 130500 33900
rect 130400 33900 130500 34000
rect 130400 34000 130500 34100
rect 130400 34100 130500 34200
rect 130400 34200 130500 34300
rect 130400 34300 130500 34400
rect 130400 34400 130500 34500
rect 130400 34500 130500 34600
rect 130400 34600 130500 34700
rect 130400 34700 130500 34800
rect 130400 34800 130500 34900
rect 130400 34900 130500 35000
rect 130400 35000 130500 35100
rect 130400 35100 130500 35200
rect 130400 35200 130500 35300
rect 130400 35300 130500 35400
rect 130400 35400 130500 35500
rect 130400 35500 130500 35600
rect 130400 35600 130500 35700
rect 130400 35700 130500 35800
rect 130400 35800 130500 35900
rect 130400 35900 130500 36000
rect 130400 36000 130500 36100
rect 130400 36100 130500 36200
rect 130400 36200 130500 36300
rect 130400 36300 130500 36400
rect 130400 37500 130500 37600
rect 130400 37600 130500 37700
rect 130400 37700 130500 37800
rect 130400 37800 130500 37900
rect 130400 37900 130500 38000
rect 130400 38000 130500 38100
rect 130400 38100 130500 38200
rect 130400 38200 130500 38300
rect 130400 38300 130500 38400
rect 130400 38400 130500 38500
rect 130400 38500 130500 38600
rect 130400 38600 130500 38700
rect 130400 38700 130500 38800
rect 130400 38800 130500 38900
rect 130400 38900 130500 39000
rect 130400 39000 130500 39100
rect 130400 39100 130500 39200
rect 130400 39200 130500 39300
rect 130400 39300 130500 39400
rect 130500 33200 130600 33300
rect 130500 33300 130600 33400
rect 130500 33400 130600 33500
rect 130500 33500 130600 33600
rect 130500 33600 130600 33700
rect 130500 33700 130600 33800
rect 130500 33800 130600 33900
rect 130500 33900 130600 34000
rect 130500 34000 130600 34100
rect 130500 34100 130600 34200
rect 130500 34200 130600 34300
rect 130500 34300 130600 34400
rect 130500 34400 130600 34500
rect 130500 34500 130600 34600
rect 130500 34600 130600 34700
rect 130500 34700 130600 34800
rect 130500 34800 130600 34900
rect 130500 34900 130600 35000
rect 130500 35000 130600 35100
rect 130500 35100 130600 35200
rect 130500 35200 130600 35300
rect 130500 35300 130600 35400
rect 130500 35400 130600 35500
rect 130500 35500 130600 35600
rect 130500 35600 130600 35700
rect 130500 35700 130600 35800
rect 130500 35800 130600 35900
rect 130500 35900 130600 36000
rect 130500 36000 130600 36100
rect 130500 36100 130600 36200
rect 130500 36200 130600 36300
rect 130500 37600 130600 37700
rect 130500 37700 130600 37800
rect 130500 37800 130600 37900
rect 130500 37900 130600 38000
rect 130500 38000 130600 38100
rect 130500 38100 130600 38200
rect 130500 38200 130600 38300
rect 130500 38300 130600 38400
rect 130500 38400 130600 38500
rect 130500 38500 130600 38600
rect 130500 38600 130600 38700
rect 130500 38700 130600 38800
rect 130500 38800 130600 38900
rect 130500 38900 130600 39000
rect 130500 39000 130600 39100
rect 130500 39100 130600 39200
rect 130500 39200 130600 39300
rect 130500 39300 130600 39400
rect 130500 39400 130600 39500
rect 130600 33400 130700 33500
rect 130600 33500 130700 33600
rect 130600 33600 130700 33700
rect 130600 33700 130700 33800
rect 130600 33800 130700 33900
rect 130600 33900 130700 34000
rect 130600 34000 130700 34100
rect 130600 34100 130700 34200
rect 130600 34200 130700 34300
rect 130600 34300 130700 34400
rect 130600 34400 130700 34500
rect 130600 34500 130700 34600
rect 130600 34600 130700 34700
rect 130600 34700 130700 34800
rect 130600 34800 130700 34900
rect 130600 34900 130700 35000
rect 130600 35000 130700 35100
rect 130600 35100 130700 35200
rect 130600 35200 130700 35300
rect 130600 35300 130700 35400
rect 130600 35400 130700 35500
rect 130600 35500 130700 35600
rect 130600 35600 130700 35700
rect 130600 35700 130700 35800
rect 130600 35800 130700 35900
rect 130600 35900 130700 36000
rect 130600 36000 130700 36100
rect 130600 36100 130700 36200
rect 130600 36200 130700 36300
rect 130600 37600 130700 37700
rect 130600 37700 130700 37800
rect 130600 37800 130700 37900
rect 130600 37900 130700 38000
rect 130600 38000 130700 38100
rect 130600 38100 130700 38200
rect 130600 38200 130700 38300
rect 130600 38300 130700 38400
rect 130600 38400 130700 38500
rect 130600 38500 130700 38600
rect 130600 38600 130700 38700
rect 130600 38700 130700 38800
rect 130600 38800 130700 38900
rect 130600 38900 130700 39000
rect 130600 39000 130700 39100
rect 130600 39100 130700 39200
rect 130600 39200 130700 39300
rect 130600 39300 130700 39400
rect 130600 39400 130700 39500
rect 130700 33600 130800 33700
rect 130700 33700 130800 33800
rect 130700 33800 130800 33900
rect 130700 33900 130800 34000
rect 130700 34000 130800 34100
rect 130700 34100 130800 34200
rect 130700 34200 130800 34300
rect 130700 34300 130800 34400
rect 130700 34400 130800 34500
rect 130700 34500 130800 34600
rect 130700 34600 130800 34700
rect 130700 34700 130800 34800
rect 130700 34800 130800 34900
rect 130700 34900 130800 35000
rect 130700 35000 130800 35100
rect 130700 35100 130800 35200
rect 130700 35200 130800 35300
rect 130700 35300 130800 35400
rect 130700 35400 130800 35500
rect 130700 35500 130800 35600
rect 130700 35600 130800 35700
rect 130700 35700 130800 35800
rect 130700 35800 130800 35900
rect 130700 35900 130800 36000
rect 130700 36000 130800 36100
rect 130700 36100 130800 36200
rect 130700 37700 130800 37800
rect 130700 37800 130800 37900
rect 130700 37900 130800 38000
rect 130700 38000 130800 38100
rect 130700 38100 130800 38200
rect 130700 38200 130800 38300
rect 130700 38300 130800 38400
rect 130700 38400 130800 38500
rect 130700 38500 130800 38600
rect 130700 38600 130800 38700
rect 130700 38700 130800 38800
rect 130700 38800 130800 38900
rect 130700 38900 130800 39000
rect 130700 39000 130800 39100
rect 130700 39100 130800 39200
rect 130700 39200 130800 39300
rect 130700 39300 130800 39400
rect 130700 39400 130800 39500
rect 130800 33800 130900 33900
rect 130800 33900 130900 34000
rect 130800 34000 130900 34100
rect 130800 34100 130900 34200
rect 130800 34200 130900 34300
rect 130800 34300 130900 34400
rect 130800 34400 130900 34500
rect 130800 34500 130900 34600
rect 130800 34600 130900 34700
rect 130800 34700 130900 34800
rect 130800 34800 130900 34900
rect 130800 34900 130900 35000
rect 130800 35000 130900 35100
rect 130800 35100 130900 35200
rect 130800 35200 130900 35300
rect 130800 35300 130900 35400
rect 130800 35400 130900 35500
rect 130800 35500 130900 35600
rect 130800 35600 130900 35700
rect 130800 35700 130900 35800
rect 130800 35800 130900 35900
rect 130800 35900 130900 36000
rect 130800 36000 130900 36100
rect 130800 36100 130900 36200
rect 130800 37700 130900 37800
rect 130800 37800 130900 37900
rect 130800 37900 130900 38000
rect 130800 38000 130900 38100
rect 130800 38100 130900 38200
rect 130800 38200 130900 38300
rect 130800 38300 130900 38400
rect 130800 38400 130900 38500
rect 130800 38500 130900 38600
rect 130800 38600 130900 38700
rect 130800 38700 130900 38800
rect 130800 38800 130900 38900
rect 130800 38900 130900 39000
rect 130800 39000 130900 39100
rect 130800 39100 130900 39200
rect 130800 39200 130900 39300
rect 130800 39300 130900 39400
rect 130800 39400 130900 39500
rect 130900 33900 131000 34000
rect 130900 34000 131000 34100
rect 130900 34100 131000 34200
rect 130900 34200 131000 34300
rect 130900 34300 131000 34400
rect 130900 34400 131000 34500
rect 130900 34500 131000 34600
rect 130900 34600 131000 34700
rect 130900 34700 131000 34800
rect 130900 34800 131000 34900
rect 130900 34900 131000 35000
rect 130900 35000 131000 35100
rect 130900 35100 131000 35200
rect 130900 35200 131000 35300
rect 130900 35300 131000 35400
rect 130900 35400 131000 35500
rect 130900 35500 131000 35600
rect 130900 35600 131000 35700
rect 130900 35700 131000 35800
rect 130900 35800 131000 35900
rect 130900 35900 131000 36000
rect 130900 36000 131000 36100
rect 130900 36100 131000 36200
rect 130900 37700 131000 37800
rect 130900 37800 131000 37900
rect 130900 37900 131000 38000
rect 130900 38000 131000 38100
rect 130900 38100 131000 38200
rect 130900 38200 131000 38300
rect 130900 38300 131000 38400
rect 130900 38400 131000 38500
rect 130900 38500 131000 38600
rect 130900 38600 131000 38700
rect 130900 38700 131000 38800
rect 130900 38800 131000 38900
rect 130900 38900 131000 39000
rect 130900 39000 131000 39100
rect 130900 39100 131000 39200
rect 130900 39200 131000 39300
rect 130900 39300 131000 39400
rect 130900 39400 131000 39500
rect 131000 34100 131100 34200
rect 131000 34200 131100 34300
rect 131000 34300 131100 34400
rect 131000 34400 131100 34500
rect 131000 34500 131100 34600
rect 131000 34600 131100 34700
rect 131000 34700 131100 34800
rect 131000 34800 131100 34900
rect 131000 34900 131100 35000
rect 131000 35000 131100 35100
rect 131000 35100 131100 35200
rect 131000 35200 131100 35300
rect 131000 35300 131100 35400
rect 131000 35400 131100 35500
rect 131000 35500 131100 35600
rect 131000 35600 131100 35700
rect 131000 35700 131100 35800
rect 131000 35800 131100 35900
rect 131000 35900 131100 36000
rect 131000 36000 131100 36100
rect 131000 36100 131100 36200
rect 131000 37700 131100 37800
rect 131000 37800 131100 37900
rect 131000 37900 131100 38000
rect 131000 38000 131100 38100
rect 131000 38100 131100 38200
rect 131000 38200 131100 38300
rect 131000 38300 131100 38400
rect 131000 38400 131100 38500
rect 131000 38500 131100 38600
rect 131000 38600 131100 38700
rect 131000 38700 131100 38800
rect 131000 38800 131100 38900
rect 131000 38900 131100 39000
rect 131000 39000 131100 39100
rect 131000 39100 131100 39200
rect 131000 39200 131100 39300
rect 131000 39300 131100 39400
rect 131000 39400 131100 39500
rect 131100 34200 131200 34300
rect 131100 34300 131200 34400
rect 131100 34400 131200 34500
rect 131100 34500 131200 34600
rect 131100 34600 131200 34700
rect 131100 34700 131200 34800
rect 131100 34800 131200 34900
rect 131100 34900 131200 35000
rect 131100 35000 131200 35100
rect 131100 35100 131200 35200
rect 131100 35200 131200 35300
rect 131100 35300 131200 35400
rect 131100 35400 131200 35500
rect 131100 35500 131200 35600
rect 131100 35600 131200 35700
rect 131100 35700 131200 35800
rect 131100 35800 131200 35900
rect 131100 35900 131200 36000
rect 131100 36000 131200 36100
rect 131100 36100 131200 36200
rect 131100 37700 131200 37800
rect 131100 37800 131200 37900
rect 131100 37900 131200 38000
rect 131100 38000 131200 38100
rect 131100 38100 131200 38200
rect 131100 38200 131200 38300
rect 131100 38300 131200 38400
rect 131100 38400 131200 38500
rect 131100 38500 131200 38600
rect 131100 38600 131200 38700
rect 131100 38700 131200 38800
rect 131100 38800 131200 38900
rect 131100 38900 131200 39000
rect 131100 39000 131200 39100
rect 131100 39100 131200 39200
rect 131100 39200 131200 39300
rect 131100 39300 131200 39400
rect 131200 34400 131300 34500
rect 131200 34500 131300 34600
rect 131200 34600 131300 34700
rect 131200 34700 131300 34800
rect 131200 34800 131300 34900
rect 131200 34900 131300 35000
rect 131200 35000 131300 35100
rect 131200 35100 131300 35200
rect 131200 35200 131300 35300
rect 131200 35300 131300 35400
rect 131200 35400 131300 35500
rect 131200 35500 131300 35600
rect 131200 35600 131300 35700
rect 131200 35700 131300 35800
rect 131200 35800 131300 35900
rect 131200 35900 131300 36000
rect 131200 36000 131300 36100
rect 131200 36100 131300 36200
rect 131200 36200 131300 36300
rect 131200 37700 131300 37800
rect 131200 37800 131300 37900
rect 131200 37900 131300 38000
rect 131200 38000 131300 38100
rect 131200 38100 131300 38200
rect 131200 38200 131300 38300
rect 131200 38300 131300 38400
rect 131200 38400 131300 38500
rect 131200 38500 131300 38600
rect 131200 38600 131300 38700
rect 131200 38700 131300 38800
rect 131200 38800 131300 38900
rect 131200 38900 131300 39000
rect 131200 39000 131300 39100
rect 131200 39100 131300 39200
rect 131200 39200 131300 39300
rect 131200 39300 131300 39400
rect 131300 34500 131400 34600
rect 131300 34600 131400 34700
rect 131300 34700 131400 34800
rect 131300 34800 131400 34900
rect 131300 34900 131400 35000
rect 131300 35000 131400 35100
rect 131300 35100 131400 35200
rect 131300 35200 131400 35300
rect 131300 35300 131400 35400
rect 131300 35400 131400 35500
rect 131300 35500 131400 35600
rect 131300 35600 131400 35700
rect 131300 35700 131400 35800
rect 131300 35800 131400 35900
rect 131300 35900 131400 36000
rect 131300 36000 131400 36100
rect 131300 36100 131400 36200
rect 131300 36200 131400 36300
rect 131300 37700 131400 37800
rect 131300 37800 131400 37900
rect 131300 37900 131400 38000
rect 131300 38000 131400 38100
rect 131300 38100 131400 38200
rect 131300 38200 131400 38300
rect 131300 38300 131400 38400
rect 131300 38400 131400 38500
rect 131300 38500 131400 38600
rect 131300 38600 131400 38700
rect 131300 38700 131400 38800
rect 131300 38800 131400 38900
rect 131300 38900 131400 39000
rect 131300 39000 131400 39100
rect 131300 39100 131400 39200
rect 131300 39200 131400 39300
rect 131300 39300 131400 39400
rect 131400 34500 131500 34600
rect 131400 34600 131500 34700
rect 131400 34700 131500 34800
rect 131400 34800 131500 34900
rect 131400 34900 131500 35000
rect 131400 35000 131500 35100
rect 131400 35100 131500 35200
rect 131400 35200 131500 35300
rect 131400 35300 131500 35400
rect 131400 35400 131500 35500
rect 131400 35500 131500 35600
rect 131400 35600 131500 35700
rect 131400 35700 131500 35800
rect 131400 35800 131500 35900
rect 131400 35900 131500 36000
rect 131400 36000 131500 36100
rect 131400 36100 131500 36200
rect 131400 36200 131500 36300
rect 131400 36300 131500 36400
rect 131400 37600 131500 37700
rect 131400 37700 131500 37800
rect 131400 37800 131500 37900
rect 131400 37900 131500 38000
rect 131400 38000 131500 38100
rect 131400 38100 131500 38200
rect 131400 38200 131500 38300
rect 131400 38300 131500 38400
rect 131400 38400 131500 38500
rect 131400 38500 131500 38600
rect 131400 38600 131500 38700
rect 131400 38700 131500 38800
rect 131400 38800 131500 38900
rect 131400 38900 131500 39000
rect 131400 39000 131500 39100
rect 131400 39100 131500 39200
rect 131400 39200 131500 39300
rect 131400 39300 131500 39400
rect 131500 34600 131600 34700
rect 131500 34700 131600 34800
rect 131500 34800 131600 34900
rect 131500 34900 131600 35000
rect 131500 35000 131600 35100
rect 131500 35100 131600 35200
rect 131500 35200 131600 35300
rect 131500 35300 131600 35400
rect 131500 35400 131600 35500
rect 131500 35500 131600 35600
rect 131500 35600 131600 35700
rect 131500 35700 131600 35800
rect 131500 35800 131600 35900
rect 131500 35900 131600 36000
rect 131500 36000 131600 36100
rect 131500 36100 131600 36200
rect 131500 36200 131600 36300
rect 131500 36300 131600 36400
rect 131500 36400 131600 36500
rect 131500 37500 131600 37600
rect 131500 37600 131600 37700
rect 131500 37700 131600 37800
rect 131500 37800 131600 37900
rect 131500 37900 131600 38000
rect 131500 38000 131600 38100
rect 131500 38100 131600 38200
rect 131500 38200 131600 38300
rect 131500 38300 131600 38400
rect 131500 38400 131600 38500
rect 131500 38500 131600 38600
rect 131500 38600 131600 38700
rect 131500 38700 131600 38800
rect 131500 38800 131600 38900
rect 131500 38900 131600 39000
rect 131500 39000 131600 39100
rect 131500 39100 131600 39200
rect 131500 39200 131600 39300
rect 131500 39300 131600 39400
rect 131600 34700 131700 34800
rect 131600 34800 131700 34900
rect 131600 34900 131700 35000
rect 131600 35000 131700 35100
rect 131600 35100 131700 35200
rect 131600 35200 131700 35300
rect 131600 35300 131700 35400
rect 131600 35400 131700 35500
rect 131600 35500 131700 35600
rect 131600 35600 131700 35700
rect 131600 35700 131700 35800
rect 131600 35800 131700 35900
rect 131600 35900 131700 36000
rect 131600 36000 131700 36100
rect 131600 36100 131700 36200
rect 131600 36200 131700 36300
rect 131600 36300 131700 36400
rect 131600 36400 131700 36500
rect 131600 36500 131700 36600
rect 131600 36600 131700 36700
rect 131600 37200 131700 37300
rect 131600 37300 131700 37400
rect 131600 37400 131700 37500
rect 131600 37500 131700 37600
rect 131600 37600 131700 37700
rect 131600 37700 131700 37800
rect 131600 37800 131700 37900
rect 131600 37900 131700 38000
rect 131600 38000 131700 38100
rect 131600 38100 131700 38200
rect 131600 38200 131700 38300
rect 131600 38300 131700 38400
rect 131600 38400 131700 38500
rect 131600 38500 131700 38600
rect 131600 38600 131700 38700
rect 131600 38700 131700 38800
rect 131600 38800 131700 38900
rect 131600 38900 131700 39000
rect 131600 39000 131700 39100
rect 131600 39100 131700 39200
rect 131600 39200 131700 39300
rect 131700 34700 131800 34800
rect 131700 34800 131800 34900
rect 131700 34900 131800 35000
rect 131700 35000 131800 35100
rect 131700 35100 131800 35200
rect 131700 35200 131800 35300
rect 131700 35300 131800 35400
rect 131700 35400 131800 35500
rect 131700 35500 131800 35600
rect 131700 35600 131800 35700
rect 131700 35700 131800 35800
rect 131700 35800 131800 35900
rect 131700 35900 131800 36000
rect 131700 36000 131800 36100
rect 131700 36100 131800 36200
rect 131700 36200 131800 36300
rect 131700 36300 131800 36400
rect 131700 36400 131800 36500
rect 131700 36500 131800 36600
rect 131700 36600 131800 36700
rect 131700 36700 131800 36800
rect 131700 36800 131800 36900
rect 131700 36900 131800 37000
rect 131700 37000 131800 37100
rect 131700 37100 131800 37200
rect 131700 37200 131800 37300
rect 131700 37300 131800 37400
rect 131700 37400 131800 37500
rect 131700 37500 131800 37600
rect 131700 37600 131800 37700
rect 131700 37700 131800 37800
rect 131700 37800 131800 37900
rect 131700 37900 131800 38000
rect 131700 38000 131800 38100
rect 131700 38100 131800 38200
rect 131700 38200 131800 38300
rect 131700 38300 131800 38400
rect 131700 38400 131800 38500
rect 131700 38500 131800 38600
rect 131700 38600 131800 38700
rect 131700 38700 131800 38800
rect 131700 38800 131800 38900
rect 131700 38900 131800 39000
rect 131700 39000 131800 39100
rect 131700 39100 131800 39200
rect 131700 39200 131800 39300
rect 131800 34800 131900 34900
rect 131800 34900 131900 35000
rect 131800 35000 131900 35100
rect 131800 35100 131900 35200
rect 131800 35200 131900 35300
rect 131800 35300 131900 35400
rect 131800 35400 131900 35500
rect 131800 35500 131900 35600
rect 131800 35600 131900 35700
rect 131800 35700 131900 35800
rect 131800 35800 131900 35900
rect 131800 35900 131900 36000
rect 131800 36000 131900 36100
rect 131800 36100 131900 36200
rect 131800 36200 131900 36300
rect 131800 36300 131900 36400
rect 131800 36400 131900 36500
rect 131800 36500 131900 36600
rect 131800 36600 131900 36700
rect 131800 36700 131900 36800
rect 131800 36800 131900 36900
rect 131800 36900 131900 37000
rect 131800 37000 131900 37100
rect 131800 37100 131900 37200
rect 131800 37200 131900 37300
rect 131800 37300 131900 37400
rect 131800 37400 131900 37500
rect 131800 37500 131900 37600
rect 131800 37600 131900 37700
rect 131800 37700 131900 37800
rect 131800 37800 131900 37900
rect 131800 37900 131900 38000
rect 131800 38000 131900 38100
rect 131800 38100 131900 38200
rect 131800 38200 131900 38300
rect 131800 38300 131900 38400
rect 131800 38400 131900 38500
rect 131800 38500 131900 38600
rect 131800 38600 131900 38700
rect 131800 38700 131900 38800
rect 131800 38800 131900 38900
rect 131800 38900 131900 39000
rect 131800 39000 131900 39100
rect 131800 39100 131900 39200
rect 131900 34800 132000 34900
rect 131900 34900 132000 35000
rect 131900 35000 132000 35100
rect 131900 35100 132000 35200
rect 131900 35200 132000 35300
rect 131900 35300 132000 35400
rect 131900 35400 132000 35500
rect 131900 35500 132000 35600
rect 131900 35600 132000 35700
rect 131900 35700 132000 35800
rect 131900 35800 132000 35900
rect 131900 35900 132000 36000
rect 131900 36000 132000 36100
rect 131900 36100 132000 36200
rect 131900 36200 132000 36300
rect 131900 36300 132000 36400
rect 131900 36400 132000 36500
rect 131900 36500 132000 36600
rect 131900 36600 132000 36700
rect 131900 36700 132000 36800
rect 131900 36800 132000 36900
rect 131900 36900 132000 37000
rect 131900 37000 132000 37100
rect 131900 37100 132000 37200
rect 131900 37200 132000 37300
rect 131900 37300 132000 37400
rect 131900 37400 132000 37500
rect 131900 37500 132000 37600
rect 131900 37600 132000 37700
rect 131900 37700 132000 37800
rect 131900 37800 132000 37900
rect 131900 37900 132000 38000
rect 131900 38000 132000 38100
rect 131900 38100 132000 38200
rect 131900 38200 132000 38300
rect 131900 38300 132000 38400
rect 131900 38400 132000 38500
rect 131900 38500 132000 38600
rect 131900 38600 132000 38700
rect 131900 38700 132000 38800
rect 131900 38800 132000 38900
rect 131900 38900 132000 39000
rect 131900 39000 132000 39100
rect 131900 39100 132000 39200
rect 132000 34900 132100 35000
rect 132000 35000 132100 35100
rect 132000 35100 132100 35200
rect 132000 35200 132100 35300
rect 132000 35300 132100 35400
rect 132000 35400 132100 35500
rect 132000 35500 132100 35600
rect 132000 35600 132100 35700
rect 132000 35700 132100 35800
rect 132000 35800 132100 35900
rect 132000 35900 132100 36000
rect 132000 36000 132100 36100
rect 132000 36100 132100 36200
rect 132000 36200 132100 36300
rect 132000 36300 132100 36400
rect 132000 36400 132100 36500
rect 132000 36500 132100 36600
rect 132000 36600 132100 36700
rect 132000 36700 132100 36800
rect 132000 36800 132100 36900
rect 132000 36900 132100 37000
rect 132000 37000 132100 37100
rect 132000 37100 132100 37200
rect 132000 37200 132100 37300
rect 132000 37300 132100 37400
rect 132000 37400 132100 37500
rect 132000 37500 132100 37600
rect 132000 37600 132100 37700
rect 132000 37700 132100 37800
rect 132000 37800 132100 37900
rect 132000 37900 132100 38000
rect 132000 38000 132100 38100
rect 132000 38100 132100 38200
rect 132000 38200 132100 38300
rect 132000 38300 132100 38400
rect 132000 38400 132100 38500
rect 132000 38500 132100 38600
rect 132000 38600 132100 38700
rect 132000 38700 132100 38800
rect 132000 38800 132100 38900
rect 132000 38900 132100 39000
rect 132000 39000 132100 39100
rect 132100 34900 132200 35000
rect 132100 35000 132200 35100
rect 132100 35100 132200 35200
rect 132100 35200 132200 35300
rect 132100 35300 132200 35400
rect 132100 35400 132200 35500
rect 132100 35500 132200 35600
rect 132100 35600 132200 35700
rect 132100 35700 132200 35800
rect 132100 35800 132200 35900
rect 132100 35900 132200 36000
rect 132100 36000 132200 36100
rect 132100 36100 132200 36200
rect 132100 36200 132200 36300
rect 132100 36300 132200 36400
rect 132100 36400 132200 36500
rect 132100 36500 132200 36600
rect 132100 36600 132200 36700
rect 132100 36700 132200 36800
rect 132100 36800 132200 36900
rect 132100 36900 132200 37000
rect 132100 37000 132200 37100
rect 132100 37100 132200 37200
rect 132100 37200 132200 37300
rect 132100 37300 132200 37400
rect 132100 37400 132200 37500
rect 132100 37500 132200 37600
rect 132100 37600 132200 37700
rect 132100 37700 132200 37800
rect 132100 37800 132200 37900
rect 132100 37900 132200 38000
rect 132100 38000 132200 38100
rect 132100 38100 132200 38200
rect 132100 38200 132200 38300
rect 132100 38300 132200 38400
rect 132100 38400 132200 38500
rect 132100 38500 132200 38600
rect 132100 38600 132200 38700
rect 132100 38700 132200 38800
rect 132100 38800 132200 38900
rect 132100 38900 132200 39000
rect 132100 39000 132200 39100
rect 132200 35000 132300 35100
rect 132200 35100 132300 35200
rect 132200 35200 132300 35300
rect 132200 35300 132300 35400
rect 132200 35400 132300 35500
rect 132200 35500 132300 35600
rect 132200 35600 132300 35700
rect 132200 35700 132300 35800
rect 132200 35800 132300 35900
rect 132200 35900 132300 36000
rect 132200 36000 132300 36100
rect 132200 36100 132300 36200
rect 132200 36200 132300 36300
rect 132200 36300 132300 36400
rect 132200 36400 132300 36500
rect 132200 36500 132300 36600
rect 132200 36600 132300 36700
rect 132200 36700 132300 36800
rect 132200 36800 132300 36900
rect 132200 36900 132300 37000
rect 132200 37000 132300 37100
rect 132200 37100 132300 37200
rect 132200 37200 132300 37300
rect 132200 37300 132300 37400
rect 132200 37400 132300 37500
rect 132200 37500 132300 37600
rect 132200 37600 132300 37700
rect 132200 37700 132300 37800
rect 132200 37800 132300 37900
rect 132200 37900 132300 38000
rect 132200 38000 132300 38100
rect 132200 38100 132300 38200
rect 132200 38200 132300 38300
rect 132200 38300 132300 38400
rect 132200 38400 132300 38500
rect 132200 38500 132300 38600
rect 132200 38600 132300 38700
rect 132200 38700 132300 38800
rect 132200 38800 132300 38900
rect 132200 38900 132300 39000
rect 132300 35100 132400 35200
rect 132300 35200 132400 35300
rect 132300 35300 132400 35400
rect 132300 35400 132400 35500
rect 132300 35500 132400 35600
rect 132300 35600 132400 35700
rect 132300 35700 132400 35800
rect 132300 35800 132400 35900
rect 132300 35900 132400 36000
rect 132300 36000 132400 36100
rect 132300 36100 132400 36200
rect 132300 36200 132400 36300
rect 132300 36300 132400 36400
rect 132300 36400 132400 36500
rect 132300 36500 132400 36600
rect 132300 36600 132400 36700
rect 132300 36700 132400 36800
rect 132300 36800 132400 36900
rect 132300 36900 132400 37000
rect 132300 37000 132400 37100
rect 132300 37100 132400 37200
rect 132300 37200 132400 37300
rect 132300 37300 132400 37400
rect 132300 37400 132400 37500
rect 132300 37500 132400 37600
rect 132300 37600 132400 37700
rect 132300 37700 132400 37800
rect 132300 37800 132400 37900
rect 132300 37900 132400 38000
rect 132300 38000 132400 38100
rect 132300 38100 132400 38200
rect 132300 38200 132400 38300
rect 132300 38300 132400 38400
rect 132300 38400 132400 38500
rect 132300 38500 132400 38600
rect 132300 38600 132400 38700
rect 132300 38700 132400 38800
rect 132300 38800 132400 38900
rect 132300 38900 132400 39000
rect 132400 35200 132500 35300
rect 132400 35300 132500 35400
rect 132400 35400 132500 35500
rect 132400 35500 132500 35600
rect 132400 35600 132500 35700
rect 132400 35700 132500 35800
rect 132400 35800 132500 35900
rect 132400 35900 132500 36000
rect 132400 36000 132500 36100
rect 132400 36100 132500 36200
rect 132400 36200 132500 36300
rect 132400 36300 132500 36400
rect 132400 36400 132500 36500
rect 132400 36500 132500 36600
rect 132400 36600 132500 36700
rect 132400 36700 132500 36800
rect 132400 36800 132500 36900
rect 132400 36900 132500 37000
rect 132400 37000 132500 37100
rect 132400 37100 132500 37200
rect 132400 37200 132500 37300
rect 132400 37300 132500 37400
rect 132400 37400 132500 37500
rect 132400 37500 132500 37600
rect 132400 37600 132500 37700
rect 132400 37700 132500 37800
rect 132400 37800 132500 37900
rect 132400 37900 132500 38000
rect 132400 38000 132500 38100
rect 132400 38100 132500 38200
rect 132400 38200 132500 38300
rect 132400 38300 132500 38400
rect 132400 38400 132500 38500
rect 132400 38500 132500 38600
rect 132400 38600 132500 38700
rect 132400 38700 132500 38800
rect 132400 38800 132500 38900
rect 132500 35200 132600 35300
rect 132500 35300 132600 35400
rect 132500 35400 132600 35500
rect 132500 35500 132600 35600
rect 132500 35600 132600 35700
rect 132500 35700 132600 35800
rect 132500 35800 132600 35900
rect 132500 35900 132600 36000
rect 132500 36000 132600 36100
rect 132500 36100 132600 36200
rect 132500 36200 132600 36300
rect 132500 36300 132600 36400
rect 132500 36400 132600 36500
rect 132500 36500 132600 36600
rect 132500 36600 132600 36700
rect 132500 36700 132600 36800
rect 132500 36800 132600 36900
rect 132500 36900 132600 37000
rect 132500 37000 132600 37100
rect 132500 37100 132600 37200
rect 132500 37200 132600 37300
rect 132500 37300 132600 37400
rect 132500 37400 132600 37500
rect 132500 37500 132600 37600
rect 132500 37600 132600 37700
rect 132500 37700 132600 37800
rect 132500 37800 132600 37900
rect 132500 37900 132600 38000
rect 132500 38000 132600 38100
rect 132500 38100 132600 38200
rect 132500 38200 132600 38300
rect 132500 38300 132600 38400
rect 132500 38400 132600 38500
rect 132500 38500 132600 38600
rect 132500 38600 132600 38700
rect 132500 38700 132600 38800
rect 132600 35300 132700 35400
rect 132600 35400 132700 35500
rect 132600 35500 132700 35600
rect 132600 35600 132700 35700
rect 132600 35700 132700 35800
rect 132600 35800 132700 35900
rect 132600 35900 132700 36000
rect 132600 36000 132700 36100
rect 132600 36100 132700 36200
rect 132600 36200 132700 36300
rect 132600 36300 132700 36400
rect 132600 36400 132700 36500
rect 132600 36500 132700 36600
rect 132600 36600 132700 36700
rect 132600 36700 132700 36800
rect 132600 36800 132700 36900
rect 132600 36900 132700 37000
rect 132600 37000 132700 37100
rect 132600 37100 132700 37200
rect 132600 37200 132700 37300
rect 132600 37300 132700 37400
rect 132600 37400 132700 37500
rect 132600 37500 132700 37600
rect 132600 37600 132700 37700
rect 132600 37700 132700 37800
rect 132600 37800 132700 37900
rect 132600 37900 132700 38000
rect 132600 38000 132700 38100
rect 132600 38100 132700 38200
rect 132600 38200 132700 38300
rect 132600 38300 132700 38400
rect 132600 38400 132700 38500
rect 132600 38500 132700 38600
rect 132600 38600 132700 38700
rect 132700 35400 132800 35500
rect 132700 35500 132800 35600
rect 132700 35600 132800 35700
rect 132700 35700 132800 35800
rect 132700 35800 132800 35900
rect 132700 35900 132800 36000
rect 132700 36000 132800 36100
rect 132700 36100 132800 36200
rect 132700 36200 132800 36300
rect 132700 36300 132800 36400
rect 132700 36400 132800 36500
rect 132700 36500 132800 36600
rect 132700 36600 132800 36700
rect 132700 36700 132800 36800
rect 132700 36800 132800 36900
rect 132700 36900 132800 37000
rect 132700 37000 132800 37100
rect 132700 37100 132800 37200
rect 132700 37200 132800 37300
rect 132700 37300 132800 37400
rect 132700 37400 132800 37500
rect 132700 37500 132800 37600
rect 132700 37600 132800 37700
rect 132700 37700 132800 37800
rect 132700 37800 132800 37900
rect 132700 37900 132800 38000
rect 132700 38000 132800 38100
rect 132700 38100 132800 38200
rect 132700 38200 132800 38300
rect 132700 38300 132800 38400
rect 132700 38400 132800 38500
rect 132700 38500 132800 38600
rect 132800 35500 132900 35600
rect 132800 35600 132900 35700
rect 132800 35700 132900 35800
rect 132800 35800 132900 35900
rect 132800 35900 132900 36000
rect 132800 36000 132900 36100
rect 132800 36100 132900 36200
rect 132800 36200 132900 36300
rect 132800 36300 132900 36400
rect 132800 36400 132900 36500
rect 132800 36500 132900 36600
rect 132800 36600 132900 36700
rect 132800 36700 132900 36800
rect 132800 36800 132900 36900
rect 132800 36900 132900 37000
rect 132800 37000 132900 37100
rect 132800 37100 132900 37200
rect 132800 37200 132900 37300
rect 132800 37300 132900 37400
rect 132800 37400 132900 37500
rect 132800 37500 132900 37600
rect 132800 37600 132900 37700
rect 132800 37700 132900 37800
rect 132800 37800 132900 37900
rect 132800 37900 132900 38000
rect 132800 38000 132900 38100
rect 132800 38100 132900 38200
rect 132800 38200 132900 38300
rect 132800 38300 132900 38400
rect 132900 35600 133000 35700
rect 132900 35700 133000 35800
rect 132900 35800 133000 35900
rect 132900 35900 133000 36000
rect 132900 36000 133000 36100
rect 132900 36100 133000 36200
rect 132900 36200 133000 36300
rect 132900 36300 133000 36400
rect 132900 36400 133000 36500
rect 132900 36500 133000 36600
rect 132900 36600 133000 36700
rect 132900 36700 133000 36800
rect 132900 36800 133000 36900
rect 132900 36900 133000 37000
rect 132900 37000 133000 37100
rect 132900 37100 133000 37200
rect 132900 37200 133000 37300
rect 132900 37300 133000 37400
rect 132900 37400 133000 37500
rect 132900 37500 133000 37600
rect 132900 37600 133000 37700
rect 132900 37700 133000 37800
rect 132900 37800 133000 37900
rect 132900 37900 133000 38000
rect 132900 38000 133000 38100
rect 132900 38100 133000 38200
rect 132900 38200 133000 38300
rect 133000 35700 133100 35800
rect 133000 35800 133100 35900
rect 133000 35900 133100 36000
rect 133000 36000 133100 36100
rect 133000 36100 133100 36200
rect 133000 36200 133100 36300
rect 133000 36300 133100 36400
rect 133000 36400 133100 36500
rect 133000 36500 133100 36600
rect 133000 36600 133100 36700
rect 133000 36700 133100 36800
rect 133000 36800 133100 36900
rect 133000 36900 133100 37000
rect 133000 37000 133100 37100
rect 133000 37100 133100 37200
rect 133000 37200 133100 37300
rect 133000 37300 133100 37400
rect 133000 37400 133100 37500
rect 133000 37500 133100 37600
rect 133000 37600 133100 37700
rect 133000 37700 133100 37800
rect 133000 37800 133100 37900
rect 133000 37900 133100 38000
rect 133100 35800 133200 35900
rect 133100 35900 133200 36000
rect 133100 36000 133200 36100
rect 133100 36100 133200 36200
rect 133100 36200 133200 36300
rect 133100 36300 133200 36400
rect 133100 36400 133200 36500
rect 133100 36500 133200 36600
rect 133100 36600 133200 36700
rect 133100 36700 133200 36800
rect 133100 36800 133200 36900
rect 133100 36900 133200 37000
rect 133100 37000 133200 37100
rect 133100 37100 133200 37200
rect 133100 37200 133200 37300
rect 133100 37300 133200 37400
rect 133100 37400 133200 37500
rect 133100 37500 133200 37600
rect 133100 37600 133200 37700
rect 133100 37700 133200 37800
rect 133200 35900 133300 36000
rect 133200 36000 133300 36100
rect 133200 36100 133300 36200
rect 133200 36200 133300 36300
rect 133200 36300 133300 36400
rect 133200 36400 133300 36500
rect 133200 36500 133300 36600
rect 133200 36600 133300 36700
rect 133200 36700 133300 36800
rect 133200 36800 133300 36900
rect 133200 36900 133300 37000
rect 133200 37000 133300 37100
rect 133200 37100 133300 37200
rect 133200 37200 133300 37300
rect 133200 37300 133300 37400
rect 133200 37400 133300 37500
rect 133300 36000 133400 36100
rect 133300 36100 133400 36200
rect 133300 36200 133400 36300
rect 133300 36300 133400 36400
rect 133300 36400 133400 36500
rect 133300 36500 133400 36600
rect 133300 36600 133400 36700
rect 133300 36700 133400 36800
rect 133300 36800 133400 36900
rect 133300 36900 133400 37000
rect 133300 37000 133400 37100
rect 133300 37100 133400 37200
rect 133400 27700 133500 27800
rect 133400 27800 133500 27900
rect 133400 27900 133500 28000
rect 133400 28000 133500 28100
rect 133400 28100 133500 28200
rect 133400 28200 133500 28300
rect 133400 28300 133500 28400
rect 133400 28400 133500 28500
rect 133400 28500 133500 28600
rect 133400 28600 133500 28700
rect 133400 28700 133500 28800
rect 133400 28800 133500 28900
rect 133400 28900 133500 29000
rect 133400 29000 133500 29100
rect 133400 29100 133500 29200
rect 133400 29200 133500 29300
rect 133400 29300 133500 29400
rect 133400 29400 133500 29500
rect 133400 29500 133500 29600
rect 133400 29600 133500 29700
rect 133400 29700 133500 29800
rect 133400 29800 133500 29900
rect 133400 30000 133500 30100
rect 133400 36300 133500 36400
rect 133400 36400 133500 36500
rect 133400 36500 133500 36600
rect 133400 36600 133500 36700
rect 133400 36700 133500 36800
rect 133500 26900 133600 27000
rect 133500 27000 133600 27100
rect 133500 27100 133600 27200
rect 133500 27200 133600 27300
rect 133500 27300 133600 27400
rect 133500 27400 133600 27500
rect 133500 27500 133600 27600
rect 133500 27600 133600 27700
rect 133500 27700 133600 27800
rect 133500 27800 133600 27900
rect 133500 27900 133600 28000
rect 133500 28000 133600 28100
rect 133500 28100 133600 28200
rect 133500 28200 133600 28300
rect 133500 28300 133600 28400
rect 133500 28400 133600 28500
rect 133500 28500 133600 28600
rect 133500 28600 133600 28700
rect 133500 28700 133600 28800
rect 133500 28800 133600 28900
rect 133500 28900 133600 29000
rect 133500 29000 133600 29100
rect 133500 29100 133600 29200
rect 133500 29200 133600 29300
rect 133500 29300 133600 29400
rect 133500 29400 133600 29500
rect 133500 29500 133600 29600
rect 133500 29600 133600 29700
rect 133500 29700 133600 29800
rect 133500 29800 133600 29900
rect 133500 29900 133600 30000
rect 133500 30000 133600 30100
rect 133500 30100 133600 30200
rect 133500 30200 133600 30300
rect 133500 30300 133600 30400
rect 133500 30400 133600 30500
rect 133500 30500 133600 30600
rect 133500 30600 133600 30700
rect 133500 30700 133600 30800
rect 133600 26500 133700 26600
rect 133600 26600 133700 26700
rect 133600 26700 133700 26800
rect 133600 26800 133700 26900
rect 133600 26900 133700 27000
rect 133600 27000 133700 27100
rect 133600 27100 133700 27200
rect 133600 27200 133700 27300
rect 133600 27300 133700 27400
rect 133600 27400 133700 27500
rect 133600 27500 133700 27600
rect 133600 27600 133700 27700
rect 133600 27700 133700 27800
rect 133600 27800 133700 27900
rect 133600 27900 133700 28000
rect 133600 28000 133700 28100
rect 133600 28100 133700 28200
rect 133600 28200 133700 28300
rect 133600 28300 133700 28400
rect 133600 28400 133700 28500
rect 133600 28500 133700 28600
rect 133600 28600 133700 28700
rect 133600 28700 133700 28800
rect 133600 28800 133700 28900
rect 133600 28900 133700 29000
rect 133600 29000 133700 29100
rect 133600 29100 133700 29200
rect 133600 29200 133700 29300
rect 133600 29300 133700 29400
rect 133600 29400 133700 29500
rect 133600 29500 133700 29600
rect 133600 29600 133700 29700
rect 133600 29700 133700 29800
rect 133600 29800 133700 29900
rect 133600 29900 133700 30000
rect 133600 30000 133700 30100
rect 133600 30100 133700 30200
rect 133600 30200 133700 30300
rect 133600 30300 133700 30400
rect 133600 30400 133700 30500
rect 133600 30500 133700 30600
rect 133600 30600 133700 30700
rect 133600 30700 133700 30800
rect 133600 30800 133700 30900
rect 133600 30900 133700 31000
rect 133600 31000 133700 31100
rect 133600 31100 133700 31200
rect 133600 31200 133700 31300
rect 133700 26100 133800 26200
rect 133700 26200 133800 26300
rect 133700 26300 133800 26400
rect 133700 26400 133800 26500
rect 133700 26500 133800 26600
rect 133700 26600 133800 26700
rect 133700 26700 133800 26800
rect 133700 26800 133800 26900
rect 133700 26900 133800 27000
rect 133700 27000 133800 27100
rect 133700 27100 133800 27200
rect 133700 27200 133800 27300
rect 133700 27300 133800 27400
rect 133700 27400 133800 27500
rect 133700 27500 133800 27600
rect 133700 27600 133800 27700
rect 133700 27700 133800 27800
rect 133700 27800 133800 27900
rect 133700 27900 133800 28000
rect 133700 28000 133800 28100
rect 133700 28100 133800 28200
rect 133700 28200 133800 28300
rect 133700 28300 133800 28400
rect 133700 28400 133800 28500
rect 133700 28500 133800 28600
rect 133700 28600 133800 28700
rect 133700 28700 133800 28800
rect 133700 28800 133800 28900
rect 133700 28900 133800 29000
rect 133700 29000 133800 29100
rect 133700 29100 133800 29200
rect 133700 29200 133800 29300
rect 133700 29300 133800 29400
rect 133700 29400 133800 29500
rect 133700 29500 133800 29600
rect 133700 29600 133800 29700
rect 133700 29700 133800 29800
rect 133700 29800 133800 29900
rect 133700 29900 133800 30000
rect 133700 30000 133800 30100
rect 133700 30100 133800 30200
rect 133700 30200 133800 30300
rect 133700 30300 133800 30400
rect 133700 30400 133800 30500
rect 133700 30500 133800 30600
rect 133700 30600 133800 30700
rect 133700 30700 133800 30800
rect 133700 30800 133800 30900
rect 133700 30900 133800 31000
rect 133700 31000 133800 31100
rect 133700 31100 133800 31200
rect 133700 31200 133800 31300
rect 133700 31300 133800 31400
rect 133700 31400 133800 31500
rect 133700 31500 133800 31600
rect 133700 31600 133800 31700
rect 133800 25800 133900 25900
rect 133800 25900 133900 26000
rect 133800 26000 133900 26100
rect 133800 26100 133900 26200
rect 133800 26200 133900 26300
rect 133800 26300 133900 26400
rect 133800 26400 133900 26500
rect 133800 26500 133900 26600
rect 133800 26600 133900 26700
rect 133800 26700 133900 26800
rect 133800 26800 133900 26900
rect 133800 26900 133900 27000
rect 133800 27000 133900 27100
rect 133800 27100 133900 27200
rect 133800 27200 133900 27300
rect 133800 27300 133900 27400
rect 133800 27400 133900 27500
rect 133800 27500 133900 27600
rect 133800 27600 133900 27700
rect 133800 27700 133900 27800
rect 133800 27800 133900 27900
rect 133800 27900 133900 28000
rect 133800 28000 133900 28100
rect 133800 28100 133900 28200
rect 133800 28200 133900 28300
rect 133800 28300 133900 28400
rect 133800 28400 133900 28500
rect 133800 28500 133900 28600
rect 133800 28600 133900 28700
rect 133800 28700 133900 28800
rect 133800 28800 133900 28900
rect 133800 28900 133900 29000
rect 133800 29000 133900 29100
rect 133800 29100 133900 29200
rect 133800 29200 133900 29300
rect 133800 29300 133900 29400
rect 133800 29400 133900 29500
rect 133800 29500 133900 29600
rect 133800 29600 133900 29700
rect 133800 29700 133900 29800
rect 133800 29800 133900 29900
rect 133800 29900 133900 30000
rect 133800 30000 133900 30100
rect 133800 30100 133900 30200
rect 133800 30200 133900 30300
rect 133800 30300 133900 30400
rect 133800 30400 133900 30500
rect 133800 30500 133900 30600
rect 133800 30600 133900 30700
rect 133800 30700 133900 30800
rect 133800 30800 133900 30900
rect 133800 30900 133900 31000
rect 133800 31000 133900 31100
rect 133800 31100 133900 31200
rect 133800 31200 133900 31300
rect 133800 31300 133900 31400
rect 133800 31400 133900 31500
rect 133800 31500 133900 31600
rect 133800 31600 133900 31700
rect 133800 31700 133900 31800
rect 133800 31800 133900 31900
rect 133800 31900 133900 32000
rect 133800 32000 133900 32100
rect 133900 25500 134000 25600
rect 133900 25600 134000 25700
rect 133900 25700 134000 25800
rect 133900 25800 134000 25900
rect 133900 25900 134000 26000
rect 133900 26000 134000 26100
rect 133900 26100 134000 26200
rect 133900 26200 134000 26300
rect 133900 26300 134000 26400
rect 133900 26400 134000 26500
rect 133900 26500 134000 26600
rect 133900 26600 134000 26700
rect 133900 26700 134000 26800
rect 133900 26800 134000 26900
rect 133900 26900 134000 27000
rect 133900 27000 134000 27100
rect 133900 27100 134000 27200
rect 133900 27200 134000 27300
rect 133900 27300 134000 27400
rect 133900 27400 134000 27500
rect 133900 27500 134000 27600
rect 133900 27600 134000 27700
rect 133900 27700 134000 27800
rect 133900 27800 134000 27900
rect 133900 27900 134000 28000
rect 133900 28000 134000 28100
rect 133900 28100 134000 28200
rect 133900 28200 134000 28300
rect 133900 28300 134000 28400
rect 133900 28400 134000 28500
rect 133900 28500 134000 28600
rect 133900 28600 134000 28700
rect 133900 28700 134000 28800
rect 133900 28800 134000 28900
rect 133900 28900 134000 29000
rect 133900 29000 134000 29100
rect 133900 29100 134000 29200
rect 133900 29200 134000 29300
rect 133900 29300 134000 29400
rect 133900 29400 134000 29500
rect 133900 29500 134000 29600
rect 133900 29600 134000 29700
rect 133900 29700 134000 29800
rect 133900 29800 134000 29900
rect 133900 29900 134000 30000
rect 133900 30000 134000 30100
rect 133900 30100 134000 30200
rect 133900 30200 134000 30300
rect 133900 30300 134000 30400
rect 133900 30400 134000 30500
rect 133900 30500 134000 30600
rect 133900 30600 134000 30700
rect 133900 30700 134000 30800
rect 133900 30800 134000 30900
rect 133900 30900 134000 31000
rect 133900 31000 134000 31100
rect 133900 31100 134000 31200
rect 133900 31200 134000 31300
rect 133900 31300 134000 31400
rect 133900 31400 134000 31500
rect 133900 31500 134000 31600
rect 133900 31600 134000 31700
rect 133900 31700 134000 31800
rect 133900 31800 134000 31900
rect 133900 31900 134000 32000
rect 133900 32000 134000 32100
rect 133900 32100 134000 32200
rect 133900 32200 134000 32300
rect 133900 32300 134000 32400
rect 134000 25300 134100 25400
rect 134000 25400 134100 25500
rect 134000 25500 134100 25600
rect 134000 25600 134100 25700
rect 134000 25700 134100 25800
rect 134000 25800 134100 25900
rect 134000 25900 134100 26000
rect 134000 26000 134100 26100
rect 134000 26100 134100 26200
rect 134000 26200 134100 26300
rect 134000 26300 134100 26400
rect 134000 26400 134100 26500
rect 134000 26500 134100 26600
rect 134000 26600 134100 26700
rect 134000 26700 134100 26800
rect 134000 26800 134100 26900
rect 134000 26900 134100 27000
rect 134000 27000 134100 27100
rect 134000 27100 134100 27200
rect 134000 27200 134100 27300
rect 134000 27300 134100 27400
rect 134000 27400 134100 27500
rect 134000 27500 134100 27600
rect 134000 27600 134100 27700
rect 134000 27700 134100 27800
rect 134000 27800 134100 27900
rect 134000 27900 134100 28000
rect 134000 28000 134100 28100
rect 134000 28100 134100 28200
rect 134000 28200 134100 28300
rect 134000 28300 134100 28400
rect 134000 28400 134100 28500
rect 134000 28500 134100 28600
rect 134000 28600 134100 28700
rect 134000 28700 134100 28800
rect 134000 28800 134100 28900
rect 134000 28900 134100 29000
rect 134000 29000 134100 29100
rect 134000 29100 134100 29200
rect 134000 29200 134100 29300
rect 134000 29300 134100 29400
rect 134000 29400 134100 29500
rect 134000 29500 134100 29600
rect 134000 29600 134100 29700
rect 134000 29700 134100 29800
rect 134000 29800 134100 29900
rect 134000 29900 134100 30000
rect 134000 30000 134100 30100
rect 134000 30100 134100 30200
rect 134000 30200 134100 30300
rect 134000 30300 134100 30400
rect 134000 30400 134100 30500
rect 134000 30500 134100 30600
rect 134000 30600 134100 30700
rect 134000 30700 134100 30800
rect 134000 30800 134100 30900
rect 134000 30900 134100 31000
rect 134000 31000 134100 31100
rect 134000 31100 134100 31200
rect 134000 31200 134100 31300
rect 134000 31300 134100 31400
rect 134000 31400 134100 31500
rect 134000 31500 134100 31600
rect 134000 31600 134100 31700
rect 134000 31700 134100 31800
rect 134000 31800 134100 31900
rect 134000 31900 134100 32000
rect 134000 32000 134100 32100
rect 134000 32100 134100 32200
rect 134000 32200 134100 32300
rect 134000 32300 134100 32400
rect 134000 32400 134100 32500
rect 134000 32500 134100 32600
rect 134000 32600 134100 32700
rect 134100 25000 134200 25100
rect 134100 25100 134200 25200
rect 134100 25200 134200 25300
rect 134100 25300 134200 25400
rect 134100 25400 134200 25500
rect 134100 25500 134200 25600
rect 134100 25600 134200 25700
rect 134100 25700 134200 25800
rect 134100 25800 134200 25900
rect 134100 25900 134200 26000
rect 134100 26000 134200 26100
rect 134100 26100 134200 26200
rect 134100 26200 134200 26300
rect 134100 26300 134200 26400
rect 134100 26400 134200 26500
rect 134100 26500 134200 26600
rect 134100 26600 134200 26700
rect 134100 26700 134200 26800
rect 134100 26800 134200 26900
rect 134100 26900 134200 27000
rect 134100 27000 134200 27100
rect 134100 27100 134200 27200
rect 134100 27200 134200 27300
rect 134100 27300 134200 27400
rect 134100 27400 134200 27500
rect 134100 27500 134200 27600
rect 134100 27600 134200 27700
rect 134100 27700 134200 27800
rect 134100 27800 134200 27900
rect 134100 27900 134200 28000
rect 134100 28000 134200 28100
rect 134100 28100 134200 28200
rect 134100 28200 134200 28300
rect 134100 28300 134200 28400
rect 134100 28400 134200 28500
rect 134100 28500 134200 28600
rect 134100 28600 134200 28700
rect 134100 28700 134200 28800
rect 134100 28800 134200 28900
rect 134100 28900 134200 29000
rect 134100 29000 134200 29100
rect 134100 29100 134200 29200
rect 134100 29200 134200 29300
rect 134100 29300 134200 29400
rect 134100 29400 134200 29500
rect 134100 29500 134200 29600
rect 134100 29600 134200 29700
rect 134100 29700 134200 29800
rect 134100 29800 134200 29900
rect 134100 29900 134200 30000
rect 134100 30000 134200 30100
rect 134100 30100 134200 30200
rect 134100 30200 134200 30300
rect 134100 30300 134200 30400
rect 134100 30400 134200 30500
rect 134100 30500 134200 30600
rect 134100 30600 134200 30700
rect 134100 30700 134200 30800
rect 134100 30800 134200 30900
rect 134100 30900 134200 31000
rect 134100 31000 134200 31100
rect 134100 31100 134200 31200
rect 134100 31200 134200 31300
rect 134100 31300 134200 31400
rect 134100 31400 134200 31500
rect 134100 31500 134200 31600
rect 134100 31600 134200 31700
rect 134100 31700 134200 31800
rect 134100 31800 134200 31900
rect 134100 31900 134200 32000
rect 134100 32000 134200 32100
rect 134100 32100 134200 32200
rect 134100 32200 134200 32300
rect 134100 32300 134200 32400
rect 134100 32400 134200 32500
rect 134100 32500 134200 32600
rect 134100 32600 134200 32700
rect 134100 32700 134200 32800
rect 134100 32800 134200 32900
rect 134100 32900 134200 33000
rect 134200 24800 134300 24900
rect 134200 24900 134300 25000
rect 134200 25000 134300 25100
rect 134200 25100 134300 25200
rect 134200 25200 134300 25300
rect 134200 25300 134300 25400
rect 134200 25400 134300 25500
rect 134200 25500 134300 25600
rect 134200 25600 134300 25700
rect 134200 25700 134300 25800
rect 134200 25800 134300 25900
rect 134200 25900 134300 26000
rect 134200 26000 134300 26100
rect 134200 26100 134300 26200
rect 134200 26200 134300 26300
rect 134200 26300 134300 26400
rect 134200 26400 134300 26500
rect 134200 26500 134300 26600
rect 134200 26600 134300 26700
rect 134200 26700 134300 26800
rect 134200 26800 134300 26900
rect 134200 26900 134300 27000
rect 134200 27000 134300 27100
rect 134200 27100 134300 27200
rect 134200 27200 134300 27300
rect 134200 27300 134300 27400
rect 134200 27400 134300 27500
rect 134200 27500 134300 27600
rect 134200 27600 134300 27700
rect 134200 27700 134300 27800
rect 134200 27800 134300 27900
rect 134200 27900 134300 28000
rect 134200 28000 134300 28100
rect 134200 28100 134300 28200
rect 134200 28200 134300 28300
rect 134200 28300 134300 28400
rect 134200 28400 134300 28500
rect 134200 28500 134300 28600
rect 134200 28600 134300 28700
rect 134200 28700 134300 28800
rect 134200 28800 134300 28900
rect 134200 28900 134300 29000
rect 134200 29000 134300 29100
rect 134200 29100 134300 29200
rect 134200 29200 134300 29300
rect 134200 29300 134300 29400
rect 134200 29400 134300 29500
rect 134200 29500 134300 29600
rect 134200 29600 134300 29700
rect 134200 29700 134300 29800
rect 134200 29800 134300 29900
rect 134200 29900 134300 30000
rect 134200 30000 134300 30100
rect 134200 30100 134300 30200
rect 134200 30200 134300 30300
rect 134200 30300 134300 30400
rect 134200 30400 134300 30500
rect 134200 30500 134300 30600
rect 134200 30600 134300 30700
rect 134200 30700 134300 30800
rect 134200 30800 134300 30900
rect 134200 30900 134300 31000
rect 134200 31000 134300 31100
rect 134200 31100 134300 31200
rect 134200 31200 134300 31300
rect 134200 31300 134300 31400
rect 134200 31400 134300 31500
rect 134200 31500 134300 31600
rect 134200 31600 134300 31700
rect 134200 31700 134300 31800
rect 134200 31800 134300 31900
rect 134200 31900 134300 32000
rect 134200 32000 134300 32100
rect 134200 32100 134300 32200
rect 134200 32200 134300 32300
rect 134200 32300 134300 32400
rect 134200 32400 134300 32500
rect 134200 32500 134300 32600
rect 134200 32600 134300 32700
rect 134200 32700 134300 32800
rect 134200 32800 134300 32900
rect 134200 32900 134300 33000
rect 134200 33000 134300 33100
rect 134200 33100 134300 33200
rect 134200 33200 134300 33300
rect 134300 24700 134400 24800
rect 134300 24800 134400 24900
rect 134300 24900 134400 25000
rect 134300 25000 134400 25100
rect 134300 25100 134400 25200
rect 134300 25200 134400 25300
rect 134300 25300 134400 25400
rect 134300 25400 134400 25500
rect 134300 25500 134400 25600
rect 134300 25600 134400 25700
rect 134300 25700 134400 25800
rect 134300 25800 134400 25900
rect 134300 25900 134400 26000
rect 134300 26000 134400 26100
rect 134300 26100 134400 26200
rect 134300 26200 134400 26300
rect 134300 26300 134400 26400
rect 134300 26400 134400 26500
rect 134300 26500 134400 26600
rect 134300 26600 134400 26700
rect 134300 26700 134400 26800
rect 134300 26800 134400 26900
rect 134300 26900 134400 27000
rect 134300 27000 134400 27100
rect 134300 27100 134400 27200
rect 134300 27200 134400 27300
rect 134300 27300 134400 27400
rect 134300 27400 134400 27500
rect 134300 27500 134400 27600
rect 134300 27600 134400 27700
rect 134300 27700 134400 27800
rect 134300 27800 134400 27900
rect 134300 27900 134400 28000
rect 134300 28000 134400 28100
rect 134300 28100 134400 28200
rect 134300 28200 134400 28300
rect 134300 28300 134400 28400
rect 134300 28400 134400 28500
rect 134300 28500 134400 28600
rect 134300 28600 134400 28700
rect 134300 28700 134400 28800
rect 134300 28800 134400 28900
rect 134300 28900 134400 29000
rect 134300 29000 134400 29100
rect 134300 29100 134400 29200
rect 134300 29200 134400 29300
rect 134300 29300 134400 29400
rect 134300 29400 134400 29500
rect 134300 29500 134400 29600
rect 134300 29600 134400 29700
rect 134300 29700 134400 29800
rect 134300 29800 134400 29900
rect 134300 29900 134400 30000
rect 134300 30000 134400 30100
rect 134300 30100 134400 30200
rect 134300 30200 134400 30300
rect 134300 30300 134400 30400
rect 134300 30400 134400 30500
rect 134300 30500 134400 30600
rect 134300 30600 134400 30700
rect 134300 30700 134400 30800
rect 134300 30800 134400 30900
rect 134300 30900 134400 31000
rect 134300 31000 134400 31100
rect 134300 31100 134400 31200
rect 134300 31200 134400 31300
rect 134300 31300 134400 31400
rect 134300 31400 134400 31500
rect 134300 31500 134400 31600
rect 134300 31600 134400 31700
rect 134300 31700 134400 31800
rect 134300 31800 134400 31900
rect 134300 31900 134400 32000
rect 134300 32000 134400 32100
rect 134300 32100 134400 32200
rect 134300 32200 134400 32300
rect 134300 32300 134400 32400
rect 134300 32400 134400 32500
rect 134300 32500 134400 32600
rect 134300 32600 134400 32700
rect 134300 32700 134400 32800
rect 134300 32800 134400 32900
rect 134300 32900 134400 33000
rect 134300 33000 134400 33100
rect 134300 33100 134400 33200
rect 134300 33200 134400 33300
rect 134300 33300 134400 33400
rect 134300 33400 134400 33500
rect 134400 24500 134500 24600
rect 134400 24600 134500 24700
rect 134400 24700 134500 24800
rect 134400 24800 134500 24900
rect 134400 24900 134500 25000
rect 134400 25000 134500 25100
rect 134400 25100 134500 25200
rect 134400 25200 134500 25300
rect 134400 25300 134500 25400
rect 134400 25400 134500 25500
rect 134400 25500 134500 25600
rect 134400 25600 134500 25700
rect 134400 25700 134500 25800
rect 134400 25800 134500 25900
rect 134400 25900 134500 26000
rect 134400 26000 134500 26100
rect 134400 26100 134500 26200
rect 134400 26200 134500 26300
rect 134400 26300 134500 26400
rect 134400 26400 134500 26500
rect 134400 26500 134500 26600
rect 134400 26600 134500 26700
rect 134400 26700 134500 26800
rect 134400 26800 134500 26900
rect 134400 26900 134500 27000
rect 134400 27000 134500 27100
rect 134400 27100 134500 27200
rect 134400 27200 134500 27300
rect 134400 27300 134500 27400
rect 134400 27400 134500 27500
rect 134400 27500 134500 27600
rect 134400 27600 134500 27700
rect 134400 27700 134500 27800
rect 134400 27800 134500 27900
rect 134400 27900 134500 28000
rect 134400 28000 134500 28100
rect 134400 28100 134500 28200
rect 134400 28200 134500 28300
rect 134400 28300 134500 28400
rect 134400 28400 134500 28500
rect 134400 28500 134500 28600
rect 134400 28600 134500 28700
rect 134400 28700 134500 28800
rect 134400 28800 134500 28900
rect 134400 28900 134500 29000
rect 134400 29000 134500 29100
rect 134400 29100 134500 29200
rect 134400 29200 134500 29300
rect 134400 29300 134500 29400
rect 134400 29400 134500 29500
rect 134400 29500 134500 29600
rect 134400 29600 134500 29700
rect 134400 29700 134500 29800
rect 134400 29800 134500 29900
rect 134400 29900 134500 30000
rect 134400 30000 134500 30100
rect 134400 30100 134500 30200
rect 134400 30200 134500 30300
rect 134400 30300 134500 30400
rect 134400 30400 134500 30500
rect 134400 30500 134500 30600
rect 134400 30600 134500 30700
rect 134400 30700 134500 30800
rect 134400 30800 134500 30900
rect 134400 30900 134500 31000
rect 134400 31000 134500 31100
rect 134400 31100 134500 31200
rect 134400 31200 134500 31300
rect 134400 31300 134500 31400
rect 134400 31400 134500 31500
rect 134400 31500 134500 31600
rect 134400 31600 134500 31700
rect 134400 31700 134500 31800
rect 134400 31800 134500 31900
rect 134400 31900 134500 32000
rect 134400 32000 134500 32100
rect 134400 32100 134500 32200
rect 134400 32200 134500 32300
rect 134400 32300 134500 32400
rect 134400 32400 134500 32500
rect 134400 32500 134500 32600
rect 134400 32600 134500 32700
rect 134400 32700 134500 32800
rect 134400 32800 134500 32900
rect 134400 32900 134500 33000
rect 134400 33000 134500 33100
rect 134400 33100 134500 33200
rect 134400 33200 134500 33300
rect 134400 33300 134500 33400
rect 134400 33400 134500 33500
rect 134400 33500 134500 33600
rect 134400 33600 134500 33700
rect 134500 24300 134600 24400
rect 134500 24400 134600 24500
rect 134500 24500 134600 24600
rect 134500 24600 134600 24700
rect 134500 24700 134600 24800
rect 134500 24800 134600 24900
rect 134500 24900 134600 25000
rect 134500 25000 134600 25100
rect 134500 25100 134600 25200
rect 134500 25200 134600 25300
rect 134500 25300 134600 25400
rect 134500 25400 134600 25500
rect 134500 25500 134600 25600
rect 134500 25600 134600 25700
rect 134500 25700 134600 25800
rect 134500 25800 134600 25900
rect 134500 25900 134600 26000
rect 134500 26000 134600 26100
rect 134500 26100 134600 26200
rect 134500 26200 134600 26300
rect 134500 26300 134600 26400
rect 134500 26400 134600 26500
rect 134500 26500 134600 26600
rect 134500 26600 134600 26700
rect 134500 26700 134600 26800
rect 134500 26800 134600 26900
rect 134500 26900 134600 27000
rect 134500 27000 134600 27100
rect 134500 27100 134600 27200
rect 134500 27200 134600 27300
rect 134500 27300 134600 27400
rect 134500 27400 134600 27500
rect 134500 27500 134600 27600
rect 134500 27600 134600 27700
rect 134500 27700 134600 27800
rect 134500 27800 134600 27900
rect 134500 27900 134600 28000
rect 134500 28000 134600 28100
rect 134500 28100 134600 28200
rect 134500 28200 134600 28300
rect 134500 28300 134600 28400
rect 134500 28400 134600 28500
rect 134500 28500 134600 28600
rect 134500 28600 134600 28700
rect 134500 28700 134600 28800
rect 134500 28800 134600 28900
rect 134500 28900 134600 29000
rect 134500 29000 134600 29100
rect 134500 29100 134600 29200
rect 134500 29200 134600 29300
rect 134500 29300 134600 29400
rect 134500 29400 134600 29500
rect 134500 29500 134600 29600
rect 134500 29600 134600 29700
rect 134500 29700 134600 29800
rect 134500 29800 134600 29900
rect 134500 29900 134600 30000
rect 134500 30000 134600 30100
rect 134500 30100 134600 30200
rect 134500 30200 134600 30300
rect 134500 30300 134600 30400
rect 134500 30400 134600 30500
rect 134500 30500 134600 30600
rect 134500 30600 134600 30700
rect 134500 30700 134600 30800
rect 134500 30800 134600 30900
rect 134500 30900 134600 31000
rect 134500 31000 134600 31100
rect 134500 31100 134600 31200
rect 134500 31200 134600 31300
rect 134500 31300 134600 31400
rect 134500 31400 134600 31500
rect 134500 31500 134600 31600
rect 134500 31600 134600 31700
rect 134500 31700 134600 31800
rect 134500 31800 134600 31900
rect 134500 31900 134600 32000
rect 134500 32000 134600 32100
rect 134500 32100 134600 32200
rect 134500 32200 134600 32300
rect 134500 32300 134600 32400
rect 134500 32400 134600 32500
rect 134500 32500 134600 32600
rect 134500 32600 134600 32700
rect 134500 32700 134600 32800
rect 134500 32800 134600 32900
rect 134500 32900 134600 33000
rect 134500 33000 134600 33100
rect 134500 33100 134600 33200
rect 134500 33200 134600 33300
rect 134500 33300 134600 33400
rect 134500 33400 134600 33500
rect 134500 33500 134600 33600
rect 134500 33600 134600 33700
rect 134500 33700 134600 33800
rect 134500 33800 134600 33900
rect 134600 24200 134700 24300
rect 134600 24300 134700 24400
rect 134600 24400 134700 24500
rect 134600 24500 134700 24600
rect 134600 24600 134700 24700
rect 134600 24700 134700 24800
rect 134600 24800 134700 24900
rect 134600 24900 134700 25000
rect 134600 25000 134700 25100
rect 134600 25100 134700 25200
rect 134600 25200 134700 25300
rect 134600 25300 134700 25400
rect 134600 25400 134700 25500
rect 134600 25500 134700 25600
rect 134600 25600 134700 25700
rect 134600 25700 134700 25800
rect 134600 25800 134700 25900
rect 134600 25900 134700 26000
rect 134600 26000 134700 26100
rect 134600 26100 134700 26200
rect 134600 26200 134700 26300
rect 134600 26300 134700 26400
rect 134600 26400 134700 26500
rect 134600 26500 134700 26600
rect 134600 26600 134700 26700
rect 134600 26700 134700 26800
rect 134600 26800 134700 26900
rect 134600 26900 134700 27000
rect 134600 27000 134700 27100
rect 134600 27100 134700 27200
rect 134600 27200 134700 27300
rect 134600 27300 134700 27400
rect 134600 27400 134700 27500
rect 134600 27500 134700 27600
rect 134600 27600 134700 27700
rect 134600 27700 134700 27800
rect 134600 27800 134700 27900
rect 134600 27900 134700 28000
rect 134600 28000 134700 28100
rect 134600 28100 134700 28200
rect 134600 28200 134700 28300
rect 134600 28300 134700 28400
rect 134600 28400 134700 28500
rect 134600 28500 134700 28600
rect 134600 28600 134700 28700
rect 134600 28700 134700 28800
rect 134600 28800 134700 28900
rect 134600 28900 134700 29000
rect 134600 29000 134700 29100
rect 134600 29100 134700 29200
rect 134600 29200 134700 29300
rect 134600 29300 134700 29400
rect 134600 29400 134700 29500
rect 134600 29500 134700 29600
rect 134600 29600 134700 29700
rect 134600 29700 134700 29800
rect 134600 29800 134700 29900
rect 134600 29900 134700 30000
rect 134600 30000 134700 30100
rect 134600 30100 134700 30200
rect 134600 30200 134700 30300
rect 134600 30300 134700 30400
rect 134600 30400 134700 30500
rect 134600 30500 134700 30600
rect 134600 30600 134700 30700
rect 134600 30700 134700 30800
rect 134600 30800 134700 30900
rect 134600 30900 134700 31000
rect 134600 31000 134700 31100
rect 134600 31100 134700 31200
rect 134600 31200 134700 31300
rect 134600 31300 134700 31400
rect 134600 31400 134700 31500
rect 134600 31500 134700 31600
rect 134600 31600 134700 31700
rect 134600 31700 134700 31800
rect 134600 31800 134700 31900
rect 134600 31900 134700 32000
rect 134600 32000 134700 32100
rect 134600 32100 134700 32200
rect 134600 32200 134700 32300
rect 134600 32300 134700 32400
rect 134600 32400 134700 32500
rect 134600 32500 134700 32600
rect 134600 32600 134700 32700
rect 134600 32700 134700 32800
rect 134600 32800 134700 32900
rect 134600 32900 134700 33000
rect 134600 33000 134700 33100
rect 134600 33100 134700 33200
rect 134600 33200 134700 33300
rect 134600 33300 134700 33400
rect 134600 33400 134700 33500
rect 134600 33500 134700 33600
rect 134600 33600 134700 33700
rect 134600 33700 134700 33800
rect 134600 33800 134700 33900
rect 134600 33900 134700 34000
rect 134600 34000 134700 34100
rect 134700 24100 134800 24200
rect 134700 24200 134800 24300
rect 134700 24300 134800 24400
rect 134700 24400 134800 24500
rect 134700 24500 134800 24600
rect 134700 24600 134800 24700
rect 134700 24700 134800 24800
rect 134700 24800 134800 24900
rect 134700 24900 134800 25000
rect 134700 25000 134800 25100
rect 134700 25100 134800 25200
rect 134700 25200 134800 25300
rect 134700 25300 134800 25400
rect 134700 25400 134800 25500
rect 134700 25500 134800 25600
rect 134700 25600 134800 25700
rect 134700 25700 134800 25800
rect 134700 25800 134800 25900
rect 134700 25900 134800 26000
rect 134700 26000 134800 26100
rect 134700 26100 134800 26200
rect 134700 26200 134800 26300
rect 134700 26300 134800 26400
rect 134700 26400 134800 26500
rect 134700 26500 134800 26600
rect 134700 26600 134800 26700
rect 134700 26700 134800 26800
rect 134700 26800 134800 26900
rect 134700 26900 134800 27000
rect 134700 27000 134800 27100
rect 134700 27100 134800 27200
rect 134700 27200 134800 27300
rect 134700 27300 134800 27400
rect 134700 27400 134800 27500
rect 134700 27500 134800 27600
rect 134700 27600 134800 27700
rect 134700 27700 134800 27800
rect 134700 27800 134800 27900
rect 134700 27900 134800 28000
rect 134700 28000 134800 28100
rect 134700 28100 134800 28200
rect 134700 28200 134800 28300
rect 134700 28300 134800 28400
rect 134700 28400 134800 28500
rect 134700 28500 134800 28600
rect 134700 28600 134800 28700
rect 134700 28700 134800 28800
rect 134700 28800 134800 28900
rect 134700 28900 134800 29000
rect 134700 29000 134800 29100
rect 134700 29100 134800 29200
rect 134700 29200 134800 29300
rect 134700 29300 134800 29400
rect 134700 29400 134800 29500
rect 134700 29500 134800 29600
rect 134700 29600 134800 29700
rect 134700 29700 134800 29800
rect 134700 29800 134800 29900
rect 134700 29900 134800 30000
rect 134700 30000 134800 30100
rect 134700 30100 134800 30200
rect 134700 30200 134800 30300
rect 134700 30300 134800 30400
rect 134700 30400 134800 30500
rect 134700 30500 134800 30600
rect 134700 30600 134800 30700
rect 134700 30700 134800 30800
rect 134700 30800 134800 30900
rect 134700 30900 134800 31000
rect 134700 31000 134800 31100
rect 134700 31100 134800 31200
rect 134700 31200 134800 31300
rect 134700 31300 134800 31400
rect 134700 31400 134800 31500
rect 134700 31500 134800 31600
rect 134700 31600 134800 31700
rect 134700 31700 134800 31800
rect 134700 31800 134800 31900
rect 134700 31900 134800 32000
rect 134700 32000 134800 32100
rect 134700 32100 134800 32200
rect 134700 32200 134800 32300
rect 134700 32300 134800 32400
rect 134700 32400 134800 32500
rect 134700 32500 134800 32600
rect 134700 32600 134800 32700
rect 134700 32700 134800 32800
rect 134700 32800 134800 32900
rect 134700 32900 134800 33000
rect 134700 33000 134800 33100
rect 134700 33100 134800 33200
rect 134700 33200 134800 33300
rect 134700 33300 134800 33400
rect 134700 33400 134800 33500
rect 134700 33500 134800 33600
rect 134700 33600 134800 33700
rect 134700 33700 134800 33800
rect 134700 33800 134800 33900
rect 134700 33900 134800 34000
rect 134700 34000 134800 34100
rect 134700 34100 134800 34200
rect 134700 34200 134800 34300
rect 134800 23900 134900 24000
rect 134800 24000 134900 24100
rect 134800 24100 134900 24200
rect 134800 24200 134900 24300
rect 134800 24300 134900 24400
rect 134800 24400 134900 24500
rect 134800 24500 134900 24600
rect 134800 24600 134900 24700
rect 134800 24700 134900 24800
rect 134800 24800 134900 24900
rect 134800 24900 134900 25000
rect 134800 25000 134900 25100
rect 134800 25100 134900 25200
rect 134800 25200 134900 25300
rect 134800 25300 134900 25400
rect 134800 25400 134900 25500
rect 134800 25500 134900 25600
rect 134800 25600 134900 25700
rect 134800 25700 134900 25800
rect 134800 25800 134900 25900
rect 134800 25900 134900 26000
rect 134800 26000 134900 26100
rect 134800 26100 134900 26200
rect 134800 26200 134900 26300
rect 134800 26300 134900 26400
rect 134800 26400 134900 26500
rect 134800 26500 134900 26600
rect 134800 26600 134900 26700
rect 134800 26700 134900 26800
rect 134800 26800 134900 26900
rect 134800 26900 134900 27000
rect 134800 27000 134900 27100
rect 134800 27100 134900 27200
rect 134800 27200 134900 27300
rect 134800 27300 134900 27400
rect 134800 27400 134900 27500
rect 134800 27500 134900 27600
rect 134800 27600 134900 27700
rect 134800 27700 134900 27800
rect 134800 27800 134900 27900
rect 134800 27900 134900 28000
rect 134800 28000 134900 28100
rect 134800 28100 134900 28200
rect 134800 28200 134900 28300
rect 134800 28300 134900 28400
rect 134800 28400 134900 28500
rect 134800 28500 134900 28600
rect 134800 28600 134900 28700
rect 134800 28700 134900 28800
rect 134800 28800 134900 28900
rect 134800 28900 134900 29000
rect 134800 29000 134900 29100
rect 134800 29100 134900 29200
rect 134800 29200 134900 29300
rect 134800 29300 134900 29400
rect 134800 29400 134900 29500
rect 134800 29500 134900 29600
rect 134800 29600 134900 29700
rect 134800 29700 134900 29800
rect 134800 29800 134900 29900
rect 134800 29900 134900 30000
rect 134800 30000 134900 30100
rect 134800 30100 134900 30200
rect 134800 30200 134900 30300
rect 134800 30300 134900 30400
rect 134800 30400 134900 30500
rect 134800 30500 134900 30600
rect 134800 30600 134900 30700
rect 134800 30700 134900 30800
rect 134800 30800 134900 30900
rect 134800 30900 134900 31000
rect 134800 31000 134900 31100
rect 134800 31100 134900 31200
rect 134800 31200 134900 31300
rect 134800 31300 134900 31400
rect 134800 31400 134900 31500
rect 134800 31500 134900 31600
rect 134800 31600 134900 31700
rect 134800 31700 134900 31800
rect 134800 31800 134900 31900
rect 134800 31900 134900 32000
rect 134800 32000 134900 32100
rect 134800 32100 134900 32200
rect 134800 32200 134900 32300
rect 134800 32300 134900 32400
rect 134800 32400 134900 32500
rect 134800 32500 134900 32600
rect 134800 32600 134900 32700
rect 134800 32700 134900 32800
rect 134800 32800 134900 32900
rect 134800 32900 134900 33000
rect 134800 33000 134900 33100
rect 134800 33100 134900 33200
rect 134800 33200 134900 33300
rect 134800 33300 134900 33400
rect 134800 33400 134900 33500
rect 134800 33500 134900 33600
rect 134800 33600 134900 33700
rect 134800 33700 134900 33800
rect 134800 33800 134900 33900
rect 134800 33900 134900 34000
rect 134800 34000 134900 34100
rect 134800 34100 134900 34200
rect 134800 34200 134900 34300
rect 134800 34300 134900 34400
rect 134800 34400 134900 34500
rect 134900 23800 135000 23900
rect 134900 23900 135000 24000
rect 134900 24000 135000 24100
rect 134900 24100 135000 24200
rect 134900 24200 135000 24300
rect 134900 24300 135000 24400
rect 134900 24400 135000 24500
rect 134900 24500 135000 24600
rect 134900 24600 135000 24700
rect 134900 24700 135000 24800
rect 134900 24800 135000 24900
rect 134900 24900 135000 25000
rect 134900 25000 135000 25100
rect 134900 25100 135000 25200
rect 134900 25200 135000 25300
rect 134900 25300 135000 25400
rect 134900 25400 135000 25500
rect 134900 25500 135000 25600
rect 134900 25600 135000 25700
rect 134900 25700 135000 25800
rect 134900 25800 135000 25900
rect 134900 25900 135000 26000
rect 134900 26000 135000 26100
rect 134900 26100 135000 26200
rect 134900 26200 135000 26300
rect 134900 26300 135000 26400
rect 134900 26400 135000 26500
rect 134900 26500 135000 26600
rect 134900 26600 135000 26700
rect 134900 26700 135000 26800
rect 134900 26800 135000 26900
rect 134900 26900 135000 27000
rect 134900 27000 135000 27100
rect 134900 27100 135000 27200
rect 134900 27200 135000 27300
rect 134900 27300 135000 27400
rect 134900 27400 135000 27500
rect 134900 27500 135000 27600
rect 134900 27600 135000 27700
rect 134900 27700 135000 27800
rect 134900 27800 135000 27900
rect 134900 27900 135000 28000
rect 134900 28000 135000 28100
rect 134900 28100 135000 28200
rect 134900 28200 135000 28300
rect 134900 28300 135000 28400
rect 134900 28400 135000 28500
rect 134900 28500 135000 28600
rect 134900 28600 135000 28700
rect 134900 28700 135000 28800
rect 134900 28800 135000 28900
rect 134900 28900 135000 29000
rect 134900 29000 135000 29100
rect 134900 29100 135000 29200
rect 134900 29200 135000 29300
rect 134900 29300 135000 29400
rect 134900 29400 135000 29500
rect 134900 29500 135000 29600
rect 134900 29600 135000 29700
rect 134900 29700 135000 29800
rect 134900 29800 135000 29900
rect 134900 29900 135000 30000
rect 134900 30000 135000 30100
rect 134900 30100 135000 30200
rect 134900 30200 135000 30300
rect 134900 30300 135000 30400
rect 134900 30400 135000 30500
rect 134900 30500 135000 30600
rect 134900 30600 135000 30700
rect 134900 30700 135000 30800
rect 134900 30800 135000 30900
rect 134900 30900 135000 31000
rect 134900 31000 135000 31100
rect 134900 31100 135000 31200
rect 134900 31200 135000 31300
rect 134900 31300 135000 31400
rect 134900 31400 135000 31500
rect 134900 31500 135000 31600
rect 134900 31600 135000 31700
rect 134900 31700 135000 31800
rect 134900 31800 135000 31900
rect 134900 31900 135000 32000
rect 134900 32000 135000 32100
rect 134900 32100 135000 32200
rect 134900 32200 135000 32300
rect 134900 32300 135000 32400
rect 134900 32400 135000 32500
rect 134900 32500 135000 32600
rect 134900 32600 135000 32700
rect 134900 32700 135000 32800
rect 134900 32800 135000 32900
rect 134900 32900 135000 33000
rect 134900 33000 135000 33100
rect 134900 33100 135000 33200
rect 134900 33200 135000 33300
rect 134900 33300 135000 33400
rect 134900 33400 135000 33500
rect 134900 33500 135000 33600
rect 134900 33600 135000 33700
rect 134900 33700 135000 33800
rect 134900 33800 135000 33900
rect 134900 33900 135000 34000
rect 134900 34000 135000 34100
rect 134900 34100 135000 34200
rect 134900 34200 135000 34300
rect 134900 34300 135000 34400
rect 134900 34400 135000 34500
rect 134900 34500 135000 34600
rect 134900 34600 135000 34700
rect 135000 23700 135100 23800
rect 135000 23800 135100 23900
rect 135000 23900 135100 24000
rect 135000 24000 135100 24100
rect 135000 24100 135100 24200
rect 135000 24200 135100 24300
rect 135000 24300 135100 24400
rect 135000 24400 135100 24500
rect 135000 24500 135100 24600
rect 135000 24600 135100 24700
rect 135000 24700 135100 24800
rect 135000 24800 135100 24900
rect 135000 24900 135100 25000
rect 135000 25000 135100 25100
rect 135000 25100 135100 25200
rect 135000 25200 135100 25300
rect 135000 25300 135100 25400
rect 135000 25400 135100 25500
rect 135000 25500 135100 25600
rect 135000 25600 135100 25700
rect 135000 25700 135100 25800
rect 135000 25800 135100 25900
rect 135000 25900 135100 26000
rect 135000 26000 135100 26100
rect 135000 26100 135100 26200
rect 135000 26200 135100 26300
rect 135000 26300 135100 26400
rect 135000 26400 135100 26500
rect 135000 26500 135100 26600
rect 135000 26600 135100 26700
rect 135000 26700 135100 26800
rect 135000 26800 135100 26900
rect 135000 26900 135100 27000
rect 135000 27000 135100 27100
rect 135000 27100 135100 27200
rect 135000 27200 135100 27300
rect 135000 27300 135100 27400
rect 135000 27400 135100 27500
rect 135000 27500 135100 27600
rect 135000 27600 135100 27700
rect 135000 27700 135100 27800
rect 135000 27800 135100 27900
rect 135000 27900 135100 28000
rect 135000 28000 135100 28100
rect 135000 28100 135100 28200
rect 135000 28200 135100 28300
rect 135000 28300 135100 28400
rect 135000 28400 135100 28500
rect 135000 28500 135100 28600
rect 135000 28600 135100 28700
rect 135000 28700 135100 28800
rect 135000 28800 135100 28900
rect 135000 28900 135100 29000
rect 135000 29000 135100 29100
rect 135000 29100 135100 29200
rect 135000 29200 135100 29300
rect 135000 29300 135100 29400
rect 135000 29400 135100 29500
rect 135000 29500 135100 29600
rect 135000 29600 135100 29700
rect 135000 29700 135100 29800
rect 135000 29800 135100 29900
rect 135000 29900 135100 30000
rect 135000 30000 135100 30100
rect 135000 30100 135100 30200
rect 135000 30200 135100 30300
rect 135000 30300 135100 30400
rect 135000 30400 135100 30500
rect 135000 30500 135100 30600
rect 135000 30600 135100 30700
rect 135000 30700 135100 30800
rect 135000 30800 135100 30900
rect 135000 30900 135100 31000
rect 135000 31000 135100 31100
rect 135000 31100 135100 31200
rect 135000 31200 135100 31300
rect 135000 31300 135100 31400
rect 135000 31400 135100 31500
rect 135000 31500 135100 31600
rect 135000 31600 135100 31700
rect 135000 31700 135100 31800
rect 135000 31800 135100 31900
rect 135000 31900 135100 32000
rect 135000 32000 135100 32100
rect 135000 32100 135100 32200
rect 135000 32200 135100 32300
rect 135000 32300 135100 32400
rect 135000 32400 135100 32500
rect 135000 32500 135100 32600
rect 135000 32600 135100 32700
rect 135000 32700 135100 32800
rect 135000 32800 135100 32900
rect 135000 32900 135100 33000
rect 135000 33000 135100 33100
rect 135000 33100 135100 33200
rect 135000 33200 135100 33300
rect 135000 33300 135100 33400
rect 135000 33400 135100 33500
rect 135000 33500 135100 33600
rect 135000 33600 135100 33700
rect 135000 33700 135100 33800
rect 135000 33800 135100 33900
rect 135000 33900 135100 34000
rect 135000 34000 135100 34100
rect 135000 34100 135100 34200
rect 135000 34200 135100 34300
rect 135000 34300 135100 34400
rect 135000 34400 135100 34500
rect 135000 34500 135100 34600
rect 135000 34600 135100 34700
rect 135000 34700 135100 34800
rect 135000 34800 135100 34900
rect 135100 23600 135200 23700
rect 135100 23700 135200 23800
rect 135100 23800 135200 23900
rect 135100 23900 135200 24000
rect 135100 24000 135200 24100
rect 135100 24100 135200 24200
rect 135100 24200 135200 24300
rect 135100 24300 135200 24400
rect 135100 24400 135200 24500
rect 135100 24500 135200 24600
rect 135100 24600 135200 24700
rect 135100 24700 135200 24800
rect 135100 24800 135200 24900
rect 135100 24900 135200 25000
rect 135100 25000 135200 25100
rect 135100 25100 135200 25200
rect 135100 25200 135200 25300
rect 135100 25300 135200 25400
rect 135100 25400 135200 25500
rect 135100 25500 135200 25600
rect 135100 25600 135200 25700
rect 135100 25700 135200 25800
rect 135100 25800 135200 25900
rect 135100 25900 135200 26000
rect 135100 26000 135200 26100
rect 135100 26100 135200 26200
rect 135100 26200 135200 26300
rect 135100 26300 135200 26400
rect 135100 26400 135200 26500
rect 135100 26500 135200 26600
rect 135100 26600 135200 26700
rect 135100 26700 135200 26800
rect 135100 26800 135200 26900
rect 135100 26900 135200 27000
rect 135100 27000 135200 27100
rect 135100 27100 135200 27200
rect 135100 27200 135200 27300
rect 135100 27300 135200 27400
rect 135100 27400 135200 27500
rect 135100 27500 135200 27600
rect 135100 27600 135200 27700
rect 135100 27700 135200 27800
rect 135100 27800 135200 27900
rect 135100 27900 135200 28000
rect 135100 28000 135200 28100
rect 135100 28100 135200 28200
rect 135100 28200 135200 28300
rect 135100 28300 135200 28400
rect 135100 28400 135200 28500
rect 135100 28500 135200 28600
rect 135100 28600 135200 28700
rect 135100 28700 135200 28800
rect 135100 28800 135200 28900
rect 135100 28900 135200 29000
rect 135100 29000 135200 29100
rect 135100 29100 135200 29200
rect 135100 29200 135200 29300
rect 135100 29300 135200 29400
rect 135100 29400 135200 29500
rect 135100 29500 135200 29600
rect 135100 29600 135200 29700
rect 135100 29700 135200 29800
rect 135100 29800 135200 29900
rect 135100 29900 135200 30000
rect 135100 30000 135200 30100
rect 135100 30100 135200 30200
rect 135100 30200 135200 30300
rect 135100 30300 135200 30400
rect 135100 30400 135200 30500
rect 135100 30500 135200 30600
rect 135100 30600 135200 30700
rect 135100 30700 135200 30800
rect 135100 30800 135200 30900
rect 135100 30900 135200 31000
rect 135100 31000 135200 31100
rect 135100 31100 135200 31200
rect 135100 31200 135200 31300
rect 135100 31300 135200 31400
rect 135100 31400 135200 31500
rect 135100 31500 135200 31600
rect 135100 31600 135200 31700
rect 135100 31700 135200 31800
rect 135100 31800 135200 31900
rect 135100 31900 135200 32000
rect 135100 32000 135200 32100
rect 135100 32100 135200 32200
rect 135100 32200 135200 32300
rect 135100 32300 135200 32400
rect 135100 32400 135200 32500
rect 135100 32500 135200 32600
rect 135100 32600 135200 32700
rect 135100 32700 135200 32800
rect 135100 32800 135200 32900
rect 135100 32900 135200 33000
rect 135100 33000 135200 33100
rect 135100 33100 135200 33200
rect 135100 33200 135200 33300
rect 135100 33300 135200 33400
rect 135100 33400 135200 33500
rect 135100 33500 135200 33600
rect 135100 33600 135200 33700
rect 135100 33700 135200 33800
rect 135100 33800 135200 33900
rect 135100 33900 135200 34000
rect 135100 34000 135200 34100
rect 135100 34100 135200 34200
rect 135100 34200 135200 34300
rect 135100 34300 135200 34400
rect 135100 34400 135200 34500
rect 135100 34500 135200 34600
rect 135100 34600 135200 34700
rect 135100 34700 135200 34800
rect 135100 34800 135200 34900
rect 135100 34900 135200 35000
rect 135200 23500 135300 23600
rect 135200 23600 135300 23700
rect 135200 23700 135300 23800
rect 135200 23800 135300 23900
rect 135200 23900 135300 24000
rect 135200 24000 135300 24100
rect 135200 24100 135300 24200
rect 135200 24200 135300 24300
rect 135200 24300 135300 24400
rect 135200 24400 135300 24500
rect 135200 24500 135300 24600
rect 135200 24600 135300 24700
rect 135200 24700 135300 24800
rect 135200 24800 135300 24900
rect 135200 24900 135300 25000
rect 135200 25000 135300 25100
rect 135200 25100 135300 25200
rect 135200 25200 135300 25300
rect 135200 25300 135300 25400
rect 135200 25400 135300 25500
rect 135200 25500 135300 25600
rect 135200 25600 135300 25700
rect 135200 25700 135300 25800
rect 135200 25800 135300 25900
rect 135200 25900 135300 26000
rect 135200 26000 135300 26100
rect 135200 26100 135300 26200
rect 135200 26200 135300 26300
rect 135200 26300 135300 26400
rect 135200 26400 135300 26500
rect 135200 26500 135300 26600
rect 135200 26600 135300 26700
rect 135200 26700 135300 26800
rect 135200 26800 135300 26900
rect 135200 26900 135300 27000
rect 135200 27000 135300 27100
rect 135200 27100 135300 27200
rect 135200 27200 135300 27300
rect 135200 27300 135300 27400
rect 135200 27400 135300 27500
rect 135200 27500 135300 27600
rect 135200 27600 135300 27700
rect 135200 27700 135300 27800
rect 135200 27800 135300 27900
rect 135200 27900 135300 28000
rect 135200 28000 135300 28100
rect 135200 28100 135300 28200
rect 135200 28200 135300 28300
rect 135200 28300 135300 28400
rect 135200 28400 135300 28500
rect 135200 28500 135300 28600
rect 135200 28600 135300 28700
rect 135200 28700 135300 28800
rect 135200 28800 135300 28900
rect 135200 28900 135300 29000
rect 135200 29000 135300 29100
rect 135200 29100 135300 29200
rect 135200 29200 135300 29300
rect 135200 29300 135300 29400
rect 135200 29400 135300 29500
rect 135200 29500 135300 29600
rect 135200 29600 135300 29700
rect 135200 29700 135300 29800
rect 135200 29800 135300 29900
rect 135200 29900 135300 30000
rect 135200 30000 135300 30100
rect 135200 30100 135300 30200
rect 135200 30200 135300 30300
rect 135200 30300 135300 30400
rect 135200 30400 135300 30500
rect 135200 30500 135300 30600
rect 135200 30600 135300 30700
rect 135200 30700 135300 30800
rect 135200 30800 135300 30900
rect 135200 30900 135300 31000
rect 135200 31000 135300 31100
rect 135200 31100 135300 31200
rect 135200 31200 135300 31300
rect 135200 31300 135300 31400
rect 135200 31400 135300 31500
rect 135200 31500 135300 31600
rect 135200 31600 135300 31700
rect 135200 31700 135300 31800
rect 135200 31800 135300 31900
rect 135200 31900 135300 32000
rect 135200 32000 135300 32100
rect 135200 32100 135300 32200
rect 135200 32200 135300 32300
rect 135200 32300 135300 32400
rect 135200 32400 135300 32500
rect 135200 32500 135300 32600
rect 135200 32600 135300 32700
rect 135200 32700 135300 32800
rect 135200 32800 135300 32900
rect 135200 32900 135300 33000
rect 135200 33000 135300 33100
rect 135200 33100 135300 33200
rect 135200 33200 135300 33300
rect 135200 33300 135300 33400
rect 135200 33400 135300 33500
rect 135200 33500 135300 33600
rect 135200 33600 135300 33700
rect 135200 33700 135300 33800
rect 135200 33800 135300 33900
rect 135200 33900 135300 34000
rect 135200 34000 135300 34100
rect 135200 34100 135300 34200
rect 135200 34200 135300 34300
rect 135200 34300 135300 34400
rect 135200 34400 135300 34500
rect 135200 34500 135300 34600
rect 135200 34600 135300 34700
rect 135200 34700 135300 34800
rect 135200 34800 135300 34900
rect 135200 34900 135300 35000
rect 135200 35000 135300 35100
rect 135200 35100 135300 35200
rect 135300 23400 135400 23500
rect 135300 23500 135400 23600
rect 135300 23600 135400 23700
rect 135300 23700 135400 23800
rect 135300 23800 135400 23900
rect 135300 23900 135400 24000
rect 135300 24000 135400 24100
rect 135300 24100 135400 24200
rect 135300 24200 135400 24300
rect 135300 24300 135400 24400
rect 135300 24400 135400 24500
rect 135300 24500 135400 24600
rect 135300 24600 135400 24700
rect 135300 24700 135400 24800
rect 135300 24800 135400 24900
rect 135300 24900 135400 25000
rect 135300 25000 135400 25100
rect 135300 25100 135400 25200
rect 135300 25200 135400 25300
rect 135300 25300 135400 25400
rect 135300 25400 135400 25500
rect 135300 25500 135400 25600
rect 135300 25600 135400 25700
rect 135300 25700 135400 25800
rect 135300 25800 135400 25900
rect 135300 25900 135400 26000
rect 135300 26000 135400 26100
rect 135300 26100 135400 26200
rect 135300 26200 135400 26300
rect 135300 26300 135400 26400
rect 135300 26400 135400 26500
rect 135300 26500 135400 26600
rect 135300 26600 135400 26700
rect 135300 26700 135400 26800
rect 135300 26800 135400 26900
rect 135300 26900 135400 27000
rect 135300 27000 135400 27100
rect 135300 27100 135400 27200
rect 135300 27200 135400 27300
rect 135300 27300 135400 27400
rect 135300 27400 135400 27500
rect 135300 27500 135400 27600
rect 135300 27600 135400 27700
rect 135300 27700 135400 27800
rect 135300 27800 135400 27900
rect 135300 27900 135400 28000
rect 135300 28000 135400 28100
rect 135300 28100 135400 28200
rect 135300 28200 135400 28300
rect 135300 28300 135400 28400
rect 135300 28400 135400 28500
rect 135300 28500 135400 28600
rect 135300 28600 135400 28700
rect 135300 28700 135400 28800
rect 135300 28800 135400 28900
rect 135300 28900 135400 29000
rect 135300 29000 135400 29100
rect 135300 29100 135400 29200
rect 135300 29200 135400 29300
rect 135300 29300 135400 29400
rect 135300 29400 135400 29500
rect 135300 29500 135400 29600
rect 135300 29600 135400 29700
rect 135300 29700 135400 29800
rect 135300 29800 135400 29900
rect 135300 29900 135400 30000
rect 135300 30000 135400 30100
rect 135300 30100 135400 30200
rect 135300 30200 135400 30300
rect 135300 30300 135400 30400
rect 135300 30400 135400 30500
rect 135300 30500 135400 30600
rect 135300 30600 135400 30700
rect 135300 30700 135400 30800
rect 135300 30800 135400 30900
rect 135300 30900 135400 31000
rect 135300 31000 135400 31100
rect 135300 31100 135400 31200
rect 135300 31200 135400 31300
rect 135300 31300 135400 31400
rect 135300 31400 135400 31500
rect 135300 31500 135400 31600
rect 135300 31600 135400 31700
rect 135300 31700 135400 31800
rect 135300 31800 135400 31900
rect 135300 31900 135400 32000
rect 135300 32000 135400 32100
rect 135300 32100 135400 32200
rect 135300 32200 135400 32300
rect 135300 32300 135400 32400
rect 135300 32400 135400 32500
rect 135300 32500 135400 32600
rect 135300 32600 135400 32700
rect 135300 32700 135400 32800
rect 135300 32800 135400 32900
rect 135300 32900 135400 33000
rect 135300 33000 135400 33100
rect 135300 33100 135400 33200
rect 135300 33200 135400 33300
rect 135300 33300 135400 33400
rect 135300 33400 135400 33500
rect 135300 33500 135400 33600
rect 135300 33600 135400 33700
rect 135300 33700 135400 33800
rect 135300 33800 135400 33900
rect 135300 33900 135400 34000
rect 135300 34000 135400 34100
rect 135300 34100 135400 34200
rect 135300 34200 135400 34300
rect 135300 34300 135400 34400
rect 135300 34400 135400 34500
rect 135300 34500 135400 34600
rect 135300 34600 135400 34700
rect 135300 34700 135400 34800
rect 135300 34800 135400 34900
rect 135300 34900 135400 35000
rect 135300 35000 135400 35100
rect 135300 35100 135400 35200
rect 135300 35200 135400 35300
rect 135400 23300 135500 23400
rect 135400 23400 135500 23500
rect 135400 23500 135500 23600
rect 135400 23600 135500 23700
rect 135400 23700 135500 23800
rect 135400 23800 135500 23900
rect 135400 23900 135500 24000
rect 135400 24000 135500 24100
rect 135400 24100 135500 24200
rect 135400 24200 135500 24300
rect 135400 24300 135500 24400
rect 135400 24400 135500 24500
rect 135400 24500 135500 24600
rect 135400 24600 135500 24700
rect 135400 24700 135500 24800
rect 135400 24800 135500 24900
rect 135400 24900 135500 25000
rect 135400 25000 135500 25100
rect 135400 25100 135500 25200
rect 135400 25200 135500 25300
rect 135400 25300 135500 25400
rect 135400 25400 135500 25500
rect 135400 25500 135500 25600
rect 135400 25600 135500 25700
rect 135400 25700 135500 25800
rect 135400 25800 135500 25900
rect 135400 25900 135500 26000
rect 135400 26000 135500 26100
rect 135400 26100 135500 26200
rect 135400 26200 135500 26300
rect 135400 26300 135500 26400
rect 135400 26400 135500 26500
rect 135400 26500 135500 26600
rect 135400 26600 135500 26700
rect 135400 26700 135500 26800
rect 135400 26800 135500 26900
rect 135400 26900 135500 27000
rect 135400 27000 135500 27100
rect 135400 27100 135500 27200
rect 135400 27200 135500 27300
rect 135400 27300 135500 27400
rect 135400 27400 135500 27500
rect 135400 27500 135500 27600
rect 135400 27600 135500 27700
rect 135400 27700 135500 27800
rect 135400 27800 135500 27900
rect 135400 27900 135500 28000
rect 135400 28100 135500 28200
rect 135400 29600 135500 29700
rect 135400 29700 135500 29800
rect 135400 29800 135500 29900
rect 135400 29900 135500 30000
rect 135400 30000 135500 30100
rect 135400 30100 135500 30200
rect 135400 30200 135500 30300
rect 135400 30300 135500 30400
rect 135400 30400 135500 30500
rect 135400 30500 135500 30600
rect 135400 30600 135500 30700
rect 135400 30700 135500 30800
rect 135400 30800 135500 30900
rect 135400 30900 135500 31000
rect 135400 31000 135500 31100
rect 135400 31100 135500 31200
rect 135400 31200 135500 31300
rect 135400 31300 135500 31400
rect 135400 31400 135500 31500
rect 135400 31500 135500 31600
rect 135400 31600 135500 31700
rect 135400 31700 135500 31800
rect 135400 31800 135500 31900
rect 135400 31900 135500 32000
rect 135400 32000 135500 32100
rect 135400 32100 135500 32200
rect 135400 32200 135500 32300
rect 135400 32300 135500 32400
rect 135400 32400 135500 32500
rect 135400 32500 135500 32600
rect 135400 32600 135500 32700
rect 135400 32700 135500 32800
rect 135400 32800 135500 32900
rect 135400 32900 135500 33000
rect 135400 33000 135500 33100
rect 135400 33100 135500 33200
rect 135400 33200 135500 33300
rect 135400 33300 135500 33400
rect 135400 33400 135500 33500
rect 135400 33500 135500 33600
rect 135400 33600 135500 33700
rect 135400 33700 135500 33800
rect 135400 33800 135500 33900
rect 135400 33900 135500 34000
rect 135400 34000 135500 34100
rect 135400 34100 135500 34200
rect 135400 34200 135500 34300
rect 135400 34300 135500 34400
rect 135400 34400 135500 34500
rect 135400 34500 135500 34600
rect 135400 34600 135500 34700
rect 135400 34700 135500 34800
rect 135400 34800 135500 34900
rect 135400 34900 135500 35000
rect 135400 35000 135500 35100
rect 135400 35100 135500 35200
rect 135400 35200 135500 35300
rect 135400 35300 135500 35400
rect 135400 35400 135500 35500
rect 135500 23200 135600 23300
rect 135500 23300 135600 23400
rect 135500 23400 135600 23500
rect 135500 23500 135600 23600
rect 135500 23600 135600 23700
rect 135500 23700 135600 23800
rect 135500 23800 135600 23900
rect 135500 23900 135600 24000
rect 135500 24000 135600 24100
rect 135500 24100 135600 24200
rect 135500 24200 135600 24300
rect 135500 24300 135600 24400
rect 135500 24400 135600 24500
rect 135500 24500 135600 24600
rect 135500 24600 135600 24700
rect 135500 24700 135600 24800
rect 135500 24800 135600 24900
rect 135500 24900 135600 25000
rect 135500 25000 135600 25100
rect 135500 25100 135600 25200
rect 135500 25200 135600 25300
rect 135500 25300 135600 25400
rect 135500 25400 135600 25500
rect 135500 25500 135600 25600
rect 135500 25600 135600 25700
rect 135500 25700 135600 25800
rect 135500 25800 135600 25900
rect 135500 25900 135600 26000
rect 135500 26000 135600 26100
rect 135500 26100 135600 26200
rect 135500 26200 135600 26300
rect 135500 26300 135600 26400
rect 135500 26400 135600 26500
rect 135500 26500 135600 26600
rect 135500 26600 135600 26700
rect 135500 26700 135600 26800
rect 135500 26800 135600 26900
rect 135500 26900 135600 27000
rect 135500 27000 135600 27100
rect 135500 27100 135600 27200
rect 135500 27200 135600 27300
rect 135500 30400 135600 30500
rect 135500 30500 135600 30600
rect 135500 30600 135600 30700
rect 135500 30700 135600 30800
rect 135500 30800 135600 30900
rect 135500 30900 135600 31000
rect 135500 31000 135600 31100
rect 135500 31100 135600 31200
rect 135500 31200 135600 31300
rect 135500 31300 135600 31400
rect 135500 31400 135600 31500
rect 135500 31500 135600 31600
rect 135500 31600 135600 31700
rect 135500 31700 135600 31800
rect 135500 31800 135600 31900
rect 135500 31900 135600 32000
rect 135500 32000 135600 32100
rect 135500 32100 135600 32200
rect 135500 32200 135600 32300
rect 135500 32300 135600 32400
rect 135500 32400 135600 32500
rect 135500 32500 135600 32600
rect 135500 32600 135600 32700
rect 135500 32700 135600 32800
rect 135500 32800 135600 32900
rect 135500 32900 135600 33000
rect 135500 33000 135600 33100
rect 135500 33100 135600 33200
rect 135500 33200 135600 33300
rect 135500 33300 135600 33400
rect 135500 33400 135600 33500
rect 135500 33500 135600 33600
rect 135500 33600 135600 33700
rect 135500 33700 135600 33800
rect 135500 33800 135600 33900
rect 135500 33900 135600 34000
rect 135500 34000 135600 34100
rect 135500 34100 135600 34200
rect 135500 34200 135600 34300
rect 135500 34300 135600 34400
rect 135500 34400 135600 34500
rect 135500 34500 135600 34600
rect 135500 34600 135600 34700
rect 135500 34700 135600 34800
rect 135500 34800 135600 34900
rect 135500 34900 135600 35000
rect 135500 35000 135600 35100
rect 135500 35100 135600 35200
rect 135500 35200 135600 35300
rect 135500 35300 135600 35400
rect 135500 35400 135600 35500
rect 135500 35500 135600 35600
rect 135600 23100 135700 23200
rect 135600 23200 135700 23300
rect 135600 23300 135700 23400
rect 135600 23400 135700 23500
rect 135600 23500 135700 23600
rect 135600 23600 135700 23700
rect 135600 23700 135700 23800
rect 135600 23800 135700 23900
rect 135600 23900 135700 24000
rect 135600 24000 135700 24100
rect 135600 24100 135700 24200
rect 135600 24200 135700 24300
rect 135600 24300 135700 24400
rect 135600 24400 135700 24500
rect 135600 24500 135700 24600
rect 135600 24600 135700 24700
rect 135600 24700 135700 24800
rect 135600 24800 135700 24900
rect 135600 24900 135700 25000
rect 135600 25000 135700 25100
rect 135600 25100 135700 25200
rect 135600 25200 135700 25300
rect 135600 25300 135700 25400
rect 135600 25400 135700 25500
rect 135600 25500 135700 25600
rect 135600 25600 135700 25700
rect 135600 25700 135700 25800
rect 135600 25800 135700 25900
rect 135600 25900 135700 26000
rect 135600 26000 135700 26100
rect 135600 26100 135700 26200
rect 135600 26200 135700 26300
rect 135600 26300 135700 26400
rect 135600 26400 135700 26500
rect 135600 26500 135700 26600
rect 135600 26600 135700 26700
rect 135600 26700 135700 26800
rect 135600 30900 135700 31000
rect 135600 31000 135700 31100
rect 135600 31100 135700 31200
rect 135600 31200 135700 31300
rect 135600 31300 135700 31400
rect 135600 31400 135700 31500
rect 135600 31500 135700 31600
rect 135600 31600 135700 31700
rect 135600 31700 135700 31800
rect 135600 31800 135700 31900
rect 135600 31900 135700 32000
rect 135600 32000 135700 32100
rect 135600 32100 135700 32200
rect 135600 32200 135700 32300
rect 135600 32300 135700 32400
rect 135600 32400 135700 32500
rect 135600 32500 135700 32600
rect 135600 32600 135700 32700
rect 135600 32700 135700 32800
rect 135600 32800 135700 32900
rect 135600 32900 135700 33000
rect 135600 33000 135700 33100
rect 135600 33100 135700 33200
rect 135600 33200 135700 33300
rect 135600 33300 135700 33400
rect 135600 33400 135700 33500
rect 135600 33500 135700 33600
rect 135600 33600 135700 33700
rect 135600 33700 135700 33800
rect 135600 33800 135700 33900
rect 135600 33900 135700 34000
rect 135600 34000 135700 34100
rect 135600 34100 135700 34200
rect 135600 34200 135700 34300
rect 135600 34300 135700 34400
rect 135600 34400 135700 34500
rect 135600 34500 135700 34600
rect 135600 34600 135700 34700
rect 135600 34700 135700 34800
rect 135600 34800 135700 34900
rect 135600 34900 135700 35000
rect 135600 35000 135700 35100
rect 135600 35100 135700 35200
rect 135600 35200 135700 35300
rect 135600 35300 135700 35400
rect 135600 35400 135700 35500
rect 135600 35500 135700 35600
rect 135600 35600 135700 35700
rect 135600 35700 135700 35800
rect 135700 23000 135800 23100
rect 135700 23100 135800 23200
rect 135700 23200 135800 23300
rect 135700 23300 135800 23400
rect 135700 23400 135800 23500
rect 135700 23500 135800 23600
rect 135700 23600 135800 23700
rect 135700 23700 135800 23800
rect 135700 23800 135800 23900
rect 135700 23900 135800 24000
rect 135700 24000 135800 24100
rect 135700 24100 135800 24200
rect 135700 24200 135800 24300
rect 135700 24300 135800 24400
rect 135700 24400 135800 24500
rect 135700 24500 135800 24600
rect 135700 24600 135800 24700
rect 135700 24700 135800 24800
rect 135700 24800 135800 24900
rect 135700 24900 135800 25000
rect 135700 25000 135800 25100
rect 135700 25100 135800 25200
rect 135700 25200 135800 25300
rect 135700 25300 135800 25400
rect 135700 25400 135800 25500
rect 135700 25500 135800 25600
rect 135700 25600 135800 25700
rect 135700 25700 135800 25800
rect 135700 25800 135800 25900
rect 135700 25900 135800 26000
rect 135700 26000 135800 26100
rect 135700 26100 135800 26200
rect 135700 26200 135800 26300
rect 135700 26300 135800 26400
rect 135700 26400 135800 26500
rect 135700 31300 135800 31400
rect 135700 31400 135800 31500
rect 135700 31500 135800 31600
rect 135700 31600 135800 31700
rect 135700 31700 135800 31800
rect 135700 31800 135800 31900
rect 135700 31900 135800 32000
rect 135700 32000 135800 32100
rect 135700 32100 135800 32200
rect 135700 32200 135800 32300
rect 135700 32300 135800 32400
rect 135700 32400 135800 32500
rect 135700 32500 135800 32600
rect 135700 32600 135800 32700
rect 135700 32700 135800 32800
rect 135700 32800 135800 32900
rect 135700 32900 135800 33000
rect 135700 33000 135800 33100
rect 135700 33100 135800 33200
rect 135700 33200 135800 33300
rect 135700 33300 135800 33400
rect 135700 33400 135800 33500
rect 135700 33500 135800 33600
rect 135700 33600 135800 33700
rect 135700 33700 135800 33800
rect 135700 33800 135800 33900
rect 135700 33900 135800 34000
rect 135700 34000 135800 34100
rect 135700 34100 135800 34200
rect 135700 34200 135800 34300
rect 135700 34300 135800 34400
rect 135700 34400 135800 34500
rect 135700 34500 135800 34600
rect 135700 34600 135800 34700
rect 135700 34700 135800 34800
rect 135700 34800 135800 34900
rect 135700 34900 135800 35000
rect 135700 35000 135800 35100
rect 135700 35100 135800 35200
rect 135700 35200 135800 35300
rect 135700 35300 135800 35400
rect 135700 35400 135800 35500
rect 135700 35500 135800 35600
rect 135700 35600 135800 35700
rect 135700 35700 135800 35800
rect 135700 35800 135800 35900
rect 135800 23000 135900 23100
rect 135800 23100 135900 23200
rect 135800 23200 135900 23300
rect 135800 23300 135900 23400
rect 135800 23400 135900 23500
rect 135800 23500 135900 23600
rect 135800 23600 135900 23700
rect 135800 23700 135900 23800
rect 135800 23800 135900 23900
rect 135800 23900 135900 24000
rect 135800 24000 135900 24100
rect 135800 24100 135900 24200
rect 135800 24200 135900 24300
rect 135800 24300 135900 24400
rect 135800 24400 135900 24500
rect 135800 24500 135900 24600
rect 135800 24600 135900 24700
rect 135800 24700 135900 24800
rect 135800 24800 135900 24900
rect 135800 24900 135900 25000
rect 135800 25000 135900 25100
rect 135800 25100 135900 25200
rect 135800 25200 135900 25300
rect 135800 25300 135900 25400
rect 135800 25400 135900 25500
rect 135800 25500 135900 25600
rect 135800 25600 135900 25700
rect 135800 25700 135900 25800
rect 135800 25800 135900 25900
rect 135800 25900 135900 26000
rect 135800 26000 135900 26100
rect 135800 26100 135900 26200
rect 135800 26200 135900 26300
rect 135800 31700 135900 31800
rect 135800 31800 135900 31900
rect 135800 31900 135900 32000
rect 135800 32000 135900 32100
rect 135800 32100 135900 32200
rect 135800 32200 135900 32300
rect 135800 32300 135900 32400
rect 135800 32400 135900 32500
rect 135800 32500 135900 32600
rect 135800 32600 135900 32700
rect 135800 32700 135900 32800
rect 135800 32800 135900 32900
rect 135800 32900 135900 33000
rect 135800 33000 135900 33100
rect 135800 33100 135900 33200
rect 135800 33200 135900 33300
rect 135800 33300 135900 33400
rect 135800 33400 135900 33500
rect 135800 33500 135900 33600
rect 135800 33600 135900 33700
rect 135800 33700 135900 33800
rect 135800 33800 135900 33900
rect 135800 33900 135900 34000
rect 135800 34000 135900 34100
rect 135800 34100 135900 34200
rect 135800 34200 135900 34300
rect 135800 34300 135900 34400
rect 135800 34400 135900 34500
rect 135800 34500 135900 34600
rect 135800 34600 135900 34700
rect 135800 34700 135900 34800
rect 135800 34800 135900 34900
rect 135800 34900 135900 35000
rect 135800 35000 135900 35100
rect 135800 35100 135900 35200
rect 135800 35200 135900 35300
rect 135800 35300 135900 35400
rect 135800 35400 135900 35500
rect 135800 35500 135900 35600
rect 135800 35600 135900 35700
rect 135800 35700 135900 35800
rect 135800 35800 135900 35900
rect 135800 35900 135900 36000
rect 135900 22900 136000 23000
rect 135900 23000 136000 23100
rect 135900 23100 136000 23200
rect 135900 23200 136000 23300
rect 135900 23300 136000 23400
rect 135900 23400 136000 23500
rect 135900 23500 136000 23600
rect 135900 23600 136000 23700
rect 135900 23700 136000 23800
rect 135900 23800 136000 23900
rect 135900 23900 136000 24000
rect 135900 24000 136000 24100
rect 135900 24100 136000 24200
rect 135900 24200 136000 24300
rect 135900 24300 136000 24400
rect 135900 24400 136000 24500
rect 135900 24500 136000 24600
rect 135900 24600 136000 24700
rect 135900 24700 136000 24800
rect 135900 24800 136000 24900
rect 135900 24900 136000 25000
rect 135900 25000 136000 25100
rect 135900 25100 136000 25200
rect 135900 25200 136000 25300
rect 135900 25300 136000 25400
rect 135900 25400 136000 25500
rect 135900 25500 136000 25600
rect 135900 25600 136000 25700
rect 135900 25700 136000 25800
rect 135900 25800 136000 25900
rect 135900 25900 136000 26000
rect 135900 31900 136000 32000
rect 135900 32000 136000 32100
rect 135900 32100 136000 32200
rect 135900 32200 136000 32300
rect 135900 32300 136000 32400
rect 135900 32400 136000 32500
rect 135900 32500 136000 32600
rect 135900 32600 136000 32700
rect 135900 32700 136000 32800
rect 135900 32800 136000 32900
rect 135900 32900 136000 33000
rect 135900 33000 136000 33100
rect 135900 33100 136000 33200
rect 135900 33200 136000 33300
rect 135900 33300 136000 33400
rect 135900 33400 136000 33500
rect 135900 33500 136000 33600
rect 135900 33600 136000 33700
rect 135900 33700 136000 33800
rect 135900 33800 136000 33900
rect 135900 33900 136000 34000
rect 135900 34000 136000 34100
rect 135900 34100 136000 34200
rect 135900 34200 136000 34300
rect 135900 34300 136000 34400
rect 135900 34400 136000 34500
rect 135900 34500 136000 34600
rect 135900 34600 136000 34700
rect 135900 34700 136000 34800
rect 135900 34800 136000 34900
rect 135900 34900 136000 35000
rect 135900 35000 136000 35100
rect 135900 35100 136000 35200
rect 135900 35200 136000 35300
rect 135900 35300 136000 35400
rect 135900 35400 136000 35500
rect 135900 35500 136000 35600
rect 135900 35600 136000 35700
rect 135900 35700 136000 35800
rect 135900 35800 136000 35900
rect 135900 35900 136000 36000
rect 135900 36000 136000 36100
rect 136000 22800 136100 22900
rect 136000 22900 136100 23000
rect 136000 23000 136100 23100
rect 136000 23100 136100 23200
rect 136000 23200 136100 23300
rect 136000 23300 136100 23400
rect 136000 23400 136100 23500
rect 136000 23500 136100 23600
rect 136000 23600 136100 23700
rect 136000 23700 136100 23800
rect 136000 23800 136100 23900
rect 136000 23900 136100 24000
rect 136000 24000 136100 24100
rect 136000 24100 136100 24200
rect 136000 24200 136100 24300
rect 136000 24300 136100 24400
rect 136000 24400 136100 24500
rect 136000 24500 136100 24600
rect 136000 24600 136100 24700
rect 136000 24700 136100 24800
rect 136000 24800 136100 24900
rect 136000 24900 136100 25000
rect 136000 25000 136100 25100
rect 136000 25100 136100 25200
rect 136000 25200 136100 25300
rect 136000 25300 136100 25400
rect 136000 25400 136100 25500
rect 136000 25500 136100 25600
rect 136000 25600 136100 25700
rect 136000 25700 136100 25800
rect 136000 25800 136100 25900
rect 136000 32200 136100 32300
rect 136000 32300 136100 32400
rect 136000 32400 136100 32500
rect 136000 32500 136100 32600
rect 136000 32600 136100 32700
rect 136000 32700 136100 32800
rect 136000 32800 136100 32900
rect 136000 32900 136100 33000
rect 136000 33000 136100 33100
rect 136000 33100 136100 33200
rect 136000 33200 136100 33300
rect 136000 33300 136100 33400
rect 136000 33400 136100 33500
rect 136000 33500 136100 33600
rect 136000 33600 136100 33700
rect 136000 33700 136100 33800
rect 136000 33800 136100 33900
rect 136000 33900 136100 34000
rect 136000 34000 136100 34100
rect 136000 34100 136100 34200
rect 136000 34200 136100 34300
rect 136000 34300 136100 34400
rect 136000 34400 136100 34500
rect 136000 34500 136100 34600
rect 136000 34600 136100 34700
rect 136000 34700 136100 34800
rect 136000 34800 136100 34900
rect 136000 34900 136100 35000
rect 136000 35000 136100 35100
rect 136000 35100 136100 35200
rect 136000 35200 136100 35300
rect 136000 35300 136100 35400
rect 136000 35400 136100 35500
rect 136000 35500 136100 35600
rect 136000 35600 136100 35700
rect 136000 35700 136100 35800
rect 136000 35800 136100 35900
rect 136000 35900 136100 36000
rect 136000 36000 136100 36100
rect 136000 36100 136100 36200
rect 136100 22700 136200 22800
rect 136100 22800 136200 22900
rect 136100 22900 136200 23000
rect 136100 23000 136200 23100
rect 136100 23100 136200 23200
rect 136100 23200 136200 23300
rect 136100 23300 136200 23400
rect 136100 23400 136200 23500
rect 136100 23500 136200 23600
rect 136100 23600 136200 23700
rect 136100 23700 136200 23800
rect 136100 23800 136200 23900
rect 136100 23900 136200 24000
rect 136100 24000 136200 24100
rect 136100 24100 136200 24200
rect 136100 24200 136200 24300
rect 136100 24300 136200 24400
rect 136100 24400 136200 24500
rect 136100 24500 136200 24600
rect 136100 24600 136200 24700
rect 136100 24700 136200 24800
rect 136100 24800 136200 24900
rect 136100 24900 136200 25000
rect 136100 25000 136200 25100
rect 136100 25100 136200 25200
rect 136100 25200 136200 25300
rect 136100 25300 136200 25400
rect 136100 25400 136200 25500
rect 136100 25500 136200 25600
rect 136100 25600 136200 25700
rect 136100 32500 136200 32600
rect 136100 32600 136200 32700
rect 136100 32700 136200 32800
rect 136100 32800 136200 32900
rect 136100 32900 136200 33000
rect 136100 33000 136200 33100
rect 136100 33100 136200 33200
rect 136100 33200 136200 33300
rect 136100 33300 136200 33400
rect 136100 33400 136200 33500
rect 136100 33500 136200 33600
rect 136100 33600 136200 33700
rect 136100 33700 136200 33800
rect 136100 33800 136200 33900
rect 136100 33900 136200 34000
rect 136100 34000 136200 34100
rect 136100 34100 136200 34200
rect 136100 34200 136200 34300
rect 136100 34300 136200 34400
rect 136100 34400 136200 34500
rect 136100 34500 136200 34600
rect 136100 34600 136200 34700
rect 136100 34700 136200 34800
rect 136100 34800 136200 34900
rect 136100 34900 136200 35000
rect 136100 35000 136200 35100
rect 136100 35100 136200 35200
rect 136100 35200 136200 35300
rect 136100 35300 136200 35400
rect 136100 35400 136200 35500
rect 136100 35500 136200 35600
rect 136100 35600 136200 35700
rect 136100 35700 136200 35800
rect 136100 35800 136200 35900
rect 136100 35900 136200 36000
rect 136100 36000 136200 36100
rect 136100 36100 136200 36200
rect 136100 36200 136200 36300
rect 136200 22700 136300 22800
rect 136200 22800 136300 22900
rect 136200 22900 136300 23000
rect 136200 23000 136300 23100
rect 136200 23100 136300 23200
rect 136200 23200 136300 23300
rect 136200 23300 136300 23400
rect 136200 23400 136300 23500
rect 136200 23500 136300 23600
rect 136200 23600 136300 23700
rect 136200 23700 136300 23800
rect 136200 23800 136300 23900
rect 136200 23900 136300 24000
rect 136200 24000 136300 24100
rect 136200 24100 136300 24200
rect 136200 24200 136300 24300
rect 136200 24300 136300 24400
rect 136200 24400 136300 24500
rect 136200 24500 136300 24600
rect 136200 24600 136300 24700
rect 136200 24700 136300 24800
rect 136200 24800 136300 24900
rect 136200 24900 136300 25000
rect 136200 25000 136300 25100
rect 136200 25100 136300 25200
rect 136200 25200 136300 25300
rect 136200 25300 136300 25400
rect 136200 25400 136300 25500
rect 136200 32700 136300 32800
rect 136200 32800 136300 32900
rect 136200 32900 136300 33000
rect 136200 33000 136300 33100
rect 136200 33100 136300 33200
rect 136200 33200 136300 33300
rect 136200 33300 136300 33400
rect 136200 33400 136300 33500
rect 136200 33500 136300 33600
rect 136200 33600 136300 33700
rect 136200 33700 136300 33800
rect 136200 33800 136300 33900
rect 136200 33900 136300 34000
rect 136200 34000 136300 34100
rect 136200 34100 136300 34200
rect 136200 34200 136300 34300
rect 136200 34300 136300 34400
rect 136200 34400 136300 34500
rect 136200 34500 136300 34600
rect 136200 34600 136300 34700
rect 136200 34700 136300 34800
rect 136200 34800 136300 34900
rect 136200 34900 136300 35000
rect 136200 35000 136300 35100
rect 136200 35100 136300 35200
rect 136200 35200 136300 35300
rect 136200 35300 136300 35400
rect 136200 35400 136300 35500
rect 136200 35500 136300 35600
rect 136200 35600 136300 35700
rect 136200 35700 136300 35800
rect 136200 35800 136300 35900
rect 136200 35900 136300 36000
rect 136200 36000 136300 36100
rect 136200 36100 136300 36200
rect 136200 36200 136300 36300
rect 136200 36300 136300 36400
rect 136300 22600 136400 22700
rect 136300 22700 136400 22800
rect 136300 22800 136400 22900
rect 136300 22900 136400 23000
rect 136300 23000 136400 23100
rect 136300 23100 136400 23200
rect 136300 23200 136400 23300
rect 136300 23300 136400 23400
rect 136300 23400 136400 23500
rect 136300 23500 136400 23600
rect 136300 23600 136400 23700
rect 136300 23700 136400 23800
rect 136300 23800 136400 23900
rect 136300 23900 136400 24000
rect 136300 24000 136400 24100
rect 136300 24100 136400 24200
rect 136300 24200 136400 24300
rect 136300 24300 136400 24400
rect 136300 24400 136400 24500
rect 136300 24500 136400 24600
rect 136300 24600 136400 24700
rect 136300 24700 136400 24800
rect 136300 24800 136400 24900
rect 136300 24900 136400 25000
rect 136300 25000 136400 25100
rect 136300 25100 136400 25200
rect 136300 25200 136400 25300
rect 136300 25300 136400 25400
rect 136300 32900 136400 33000
rect 136300 33000 136400 33100
rect 136300 33100 136400 33200
rect 136300 33200 136400 33300
rect 136300 33300 136400 33400
rect 136300 33400 136400 33500
rect 136300 33500 136400 33600
rect 136300 33600 136400 33700
rect 136300 33700 136400 33800
rect 136300 33800 136400 33900
rect 136300 33900 136400 34000
rect 136300 34000 136400 34100
rect 136300 34100 136400 34200
rect 136300 34200 136400 34300
rect 136300 34300 136400 34400
rect 136300 34400 136400 34500
rect 136300 34500 136400 34600
rect 136300 34600 136400 34700
rect 136300 34700 136400 34800
rect 136300 34800 136400 34900
rect 136300 34900 136400 35000
rect 136300 35000 136400 35100
rect 136300 35100 136400 35200
rect 136300 35200 136400 35300
rect 136300 35300 136400 35400
rect 136300 35400 136400 35500
rect 136300 35500 136400 35600
rect 136300 35600 136400 35700
rect 136300 35700 136400 35800
rect 136300 35800 136400 35900
rect 136300 35900 136400 36000
rect 136300 36000 136400 36100
rect 136300 36100 136400 36200
rect 136300 36200 136400 36300
rect 136300 36300 136400 36400
rect 136300 36400 136400 36500
rect 136400 22500 136500 22600
rect 136400 22600 136500 22700
rect 136400 22700 136500 22800
rect 136400 22800 136500 22900
rect 136400 22900 136500 23000
rect 136400 23000 136500 23100
rect 136400 23100 136500 23200
rect 136400 23200 136500 23300
rect 136400 23300 136500 23400
rect 136400 23400 136500 23500
rect 136400 23500 136500 23600
rect 136400 23600 136500 23700
rect 136400 23700 136500 23800
rect 136400 23800 136500 23900
rect 136400 23900 136500 24000
rect 136400 24000 136500 24100
rect 136400 24100 136500 24200
rect 136400 24200 136500 24300
rect 136400 24300 136500 24400
rect 136400 24400 136500 24500
rect 136400 24500 136500 24600
rect 136400 24600 136500 24700
rect 136400 24700 136500 24800
rect 136400 24800 136500 24900
rect 136400 24900 136500 25000
rect 136400 25000 136500 25100
rect 136400 25100 136500 25200
rect 136400 25200 136500 25300
rect 136400 33100 136500 33200
rect 136400 33200 136500 33300
rect 136400 33300 136500 33400
rect 136400 33400 136500 33500
rect 136400 33500 136500 33600
rect 136400 33600 136500 33700
rect 136400 33700 136500 33800
rect 136400 33800 136500 33900
rect 136400 33900 136500 34000
rect 136400 34000 136500 34100
rect 136400 34100 136500 34200
rect 136400 34200 136500 34300
rect 136400 34300 136500 34400
rect 136400 34400 136500 34500
rect 136400 34500 136500 34600
rect 136400 34600 136500 34700
rect 136400 34700 136500 34800
rect 136400 34800 136500 34900
rect 136400 34900 136500 35000
rect 136400 35000 136500 35100
rect 136400 35100 136500 35200
rect 136400 35200 136500 35300
rect 136400 35300 136500 35400
rect 136400 35400 136500 35500
rect 136400 35500 136500 35600
rect 136400 35600 136500 35700
rect 136400 35700 136500 35800
rect 136400 35800 136500 35900
rect 136400 35900 136500 36000
rect 136400 36000 136500 36100
rect 136400 36100 136500 36200
rect 136400 36200 136500 36300
rect 136400 36300 136500 36400
rect 136400 36400 136500 36500
rect 136400 36500 136500 36600
rect 136500 22500 136600 22600
rect 136500 22600 136600 22700
rect 136500 22700 136600 22800
rect 136500 22800 136600 22900
rect 136500 22900 136600 23000
rect 136500 23000 136600 23100
rect 136500 23100 136600 23200
rect 136500 23200 136600 23300
rect 136500 23300 136600 23400
rect 136500 23400 136600 23500
rect 136500 23500 136600 23600
rect 136500 23600 136600 23700
rect 136500 23700 136600 23800
rect 136500 23800 136600 23900
rect 136500 23900 136600 24000
rect 136500 24000 136600 24100
rect 136500 24100 136600 24200
rect 136500 24200 136600 24300
rect 136500 24300 136600 24400
rect 136500 24400 136600 24500
rect 136500 24500 136600 24600
rect 136500 24600 136600 24700
rect 136500 24700 136600 24800
rect 136500 24800 136600 24900
rect 136500 24900 136600 25000
rect 136500 25000 136600 25100
rect 136500 25100 136600 25200
rect 136500 33300 136600 33400
rect 136500 33400 136600 33500
rect 136500 33500 136600 33600
rect 136500 33600 136600 33700
rect 136500 33700 136600 33800
rect 136500 33800 136600 33900
rect 136500 33900 136600 34000
rect 136500 34000 136600 34100
rect 136500 34100 136600 34200
rect 136500 34200 136600 34300
rect 136500 34300 136600 34400
rect 136500 34400 136600 34500
rect 136500 34500 136600 34600
rect 136500 34600 136600 34700
rect 136500 34700 136600 34800
rect 136500 34800 136600 34900
rect 136500 34900 136600 35000
rect 136500 35000 136600 35100
rect 136500 35100 136600 35200
rect 136500 35200 136600 35300
rect 136500 35300 136600 35400
rect 136500 35400 136600 35500
rect 136500 35500 136600 35600
rect 136500 35600 136600 35700
rect 136500 35700 136600 35800
rect 136500 35800 136600 35900
rect 136500 35900 136600 36000
rect 136500 36000 136600 36100
rect 136500 36100 136600 36200
rect 136500 36200 136600 36300
rect 136500 36300 136600 36400
rect 136500 36400 136600 36500
rect 136500 36500 136600 36600
rect 136500 36600 136600 36700
rect 136600 22400 136700 22500
rect 136600 22500 136700 22600
rect 136600 22600 136700 22700
rect 136600 22700 136700 22800
rect 136600 22800 136700 22900
rect 136600 22900 136700 23000
rect 136600 23000 136700 23100
rect 136600 23100 136700 23200
rect 136600 23200 136700 23300
rect 136600 23300 136700 23400
rect 136600 23400 136700 23500
rect 136600 23500 136700 23600
rect 136600 23600 136700 23700
rect 136600 23700 136700 23800
rect 136600 23800 136700 23900
rect 136600 23900 136700 24000
rect 136600 24000 136700 24100
rect 136600 24100 136700 24200
rect 136600 24200 136700 24300
rect 136600 24300 136700 24400
rect 136600 24400 136700 24500
rect 136600 24500 136700 24600
rect 136600 24600 136700 24700
rect 136600 24700 136700 24800
rect 136600 24800 136700 24900
rect 136600 24900 136700 25000
rect 136600 25000 136700 25100
rect 136600 33500 136700 33600
rect 136600 33600 136700 33700
rect 136600 33700 136700 33800
rect 136600 33800 136700 33900
rect 136600 33900 136700 34000
rect 136600 34000 136700 34100
rect 136600 34100 136700 34200
rect 136600 34200 136700 34300
rect 136600 34300 136700 34400
rect 136600 34400 136700 34500
rect 136600 34500 136700 34600
rect 136600 34600 136700 34700
rect 136600 34700 136700 34800
rect 136600 34800 136700 34900
rect 136600 34900 136700 35000
rect 136600 35000 136700 35100
rect 136600 35100 136700 35200
rect 136600 35200 136700 35300
rect 136600 35300 136700 35400
rect 136600 35400 136700 35500
rect 136600 35500 136700 35600
rect 136600 35600 136700 35700
rect 136600 35700 136700 35800
rect 136600 35800 136700 35900
rect 136600 35900 136700 36000
rect 136600 36000 136700 36100
rect 136600 36100 136700 36200
rect 136600 36200 136700 36300
rect 136600 36300 136700 36400
rect 136600 36400 136700 36500
rect 136600 36500 136700 36600
rect 136600 36600 136700 36700
rect 136600 36700 136700 36800
rect 136700 22400 136800 22500
rect 136700 22500 136800 22600
rect 136700 22600 136800 22700
rect 136700 22700 136800 22800
rect 136700 22800 136800 22900
rect 136700 22900 136800 23000
rect 136700 23000 136800 23100
rect 136700 23100 136800 23200
rect 136700 23200 136800 23300
rect 136700 23300 136800 23400
rect 136700 23400 136800 23500
rect 136700 23500 136800 23600
rect 136700 23600 136800 23700
rect 136700 23700 136800 23800
rect 136700 23800 136800 23900
rect 136700 23900 136800 24000
rect 136700 24000 136800 24100
rect 136700 24100 136800 24200
rect 136700 24200 136800 24300
rect 136700 24300 136800 24400
rect 136700 24400 136800 24500
rect 136700 24500 136800 24600
rect 136700 24600 136800 24700
rect 136700 24700 136800 24800
rect 136700 24800 136800 24900
rect 136700 24900 136800 25000
rect 136700 33700 136800 33800
rect 136700 33800 136800 33900
rect 136700 33900 136800 34000
rect 136700 34000 136800 34100
rect 136700 34100 136800 34200
rect 136700 34200 136800 34300
rect 136700 34300 136800 34400
rect 136700 34400 136800 34500
rect 136700 34500 136800 34600
rect 136700 34600 136800 34700
rect 136700 34700 136800 34800
rect 136700 34800 136800 34900
rect 136700 34900 136800 35000
rect 136700 35000 136800 35100
rect 136700 35100 136800 35200
rect 136700 35200 136800 35300
rect 136700 35300 136800 35400
rect 136700 35400 136800 35500
rect 136700 35500 136800 35600
rect 136700 35600 136800 35700
rect 136700 35700 136800 35800
rect 136700 35800 136800 35900
rect 136700 35900 136800 36000
rect 136700 36000 136800 36100
rect 136700 36100 136800 36200
rect 136700 36200 136800 36300
rect 136700 36300 136800 36400
rect 136700 36400 136800 36500
rect 136700 36500 136800 36600
rect 136700 36600 136800 36700
rect 136700 36700 136800 36800
rect 136700 36800 136800 36900
rect 136800 22300 136900 22400
rect 136800 22400 136900 22500
rect 136800 22500 136900 22600
rect 136800 22600 136900 22700
rect 136800 22700 136900 22800
rect 136800 22800 136900 22900
rect 136800 22900 136900 23000
rect 136800 23000 136900 23100
rect 136800 23100 136900 23200
rect 136800 23200 136900 23300
rect 136800 23300 136900 23400
rect 136800 23400 136900 23500
rect 136800 23500 136900 23600
rect 136800 23600 136900 23700
rect 136800 23700 136900 23800
rect 136800 23800 136900 23900
rect 136800 23900 136900 24000
rect 136800 24000 136900 24100
rect 136800 24100 136900 24200
rect 136800 24200 136900 24300
rect 136800 24300 136900 24400
rect 136800 24400 136900 24500
rect 136800 24500 136900 24600
rect 136800 24600 136900 24700
rect 136800 24700 136900 24800
rect 136800 24800 136900 24900
rect 136800 33800 136900 33900
rect 136800 33900 136900 34000
rect 136800 34000 136900 34100
rect 136800 34100 136900 34200
rect 136800 34200 136900 34300
rect 136800 34300 136900 34400
rect 136800 34400 136900 34500
rect 136800 34500 136900 34600
rect 136800 34600 136900 34700
rect 136800 34700 136900 34800
rect 136800 34800 136900 34900
rect 136800 34900 136900 35000
rect 136800 35000 136900 35100
rect 136800 35100 136900 35200
rect 136800 35200 136900 35300
rect 136800 35300 136900 35400
rect 136800 35400 136900 35500
rect 136800 35500 136900 35600
rect 136800 35600 136900 35700
rect 136800 35700 136900 35800
rect 136800 35800 136900 35900
rect 136800 35900 136900 36000
rect 136800 36000 136900 36100
rect 136800 36100 136900 36200
rect 136800 36200 136900 36300
rect 136800 36300 136900 36400
rect 136800 36400 136900 36500
rect 136800 36500 136900 36600
rect 136800 36600 136900 36700
rect 136800 36700 136900 36800
rect 136800 36800 136900 36900
rect 136800 36900 136900 37000
rect 136900 22300 137000 22400
rect 136900 22400 137000 22500
rect 136900 22500 137000 22600
rect 136900 22600 137000 22700
rect 136900 22700 137000 22800
rect 136900 22800 137000 22900
rect 136900 22900 137000 23000
rect 136900 23000 137000 23100
rect 136900 23100 137000 23200
rect 136900 23200 137000 23300
rect 136900 23300 137000 23400
rect 136900 23400 137000 23500
rect 136900 23500 137000 23600
rect 136900 23600 137000 23700
rect 136900 23700 137000 23800
rect 136900 23800 137000 23900
rect 136900 23900 137000 24000
rect 136900 24000 137000 24100
rect 136900 24100 137000 24200
rect 136900 24200 137000 24300
rect 136900 24300 137000 24400
rect 136900 24400 137000 24500
rect 136900 24500 137000 24600
rect 136900 24600 137000 24700
rect 136900 24700 137000 24800
rect 136900 34000 137000 34100
rect 136900 34100 137000 34200
rect 136900 34200 137000 34300
rect 136900 34300 137000 34400
rect 136900 34400 137000 34500
rect 136900 34500 137000 34600
rect 136900 34600 137000 34700
rect 136900 34700 137000 34800
rect 136900 34800 137000 34900
rect 136900 34900 137000 35000
rect 136900 35000 137000 35100
rect 136900 35100 137000 35200
rect 136900 35200 137000 35300
rect 136900 35300 137000 35400
rect 136900 35400 137000 35500
rect 136900 35500 137000 35600
rect 136900 35600 137000 35700
rect 136900 35700 137000 35800
rect 136900 35800 137000 35900
rect 136900 35900 137000 36000
rect 136900 36000 137000 36100
rect 136900 36100 137000 36200
rect 136900 36200 137000 36300
rect 136900 36300 137000 36400
rect 136900 36400 137000 36500
rect 136900 36500 137000 36600
rect 136900 36600 137000 36700
rect 136900 36700 137000 36800
rect 136900 36800 137000 36900
rect 136900 36900 137000 37000
rect 137000 22200 137100 22300
rect 137000 22300 137100 22400
rect 137000 22400 137100 22500
rect 137000 22500 137100 22600
rect 137000 22600 137100 22700
rect 137000 22700 137100 22800
rect 137000 22800 137100 22900
rect 137000 22900 137100 23000
rect 137000 23000 137100 23100
rect 137000 23100 137100 23200
rect 137000 23200 137100 23300
rect 137000 23300 137100 23400
rect 137000 23400 137100 23500
rect 137000 23500 137100 23600
rect 137000 23600 137100 23700
rect 137000 23700 137100 23800
rect 137000 23800 137100 23900
rect 137000 23900 137100 24000
rect 137000 24000 137100 24100
rect 137000 24100 137100 24200
rect 137000 24200 137100 24300
rect 137000 24300 137100 24400
rect 137000 24400 137100 24500
rect 137000 24500 137100 24600
rect 137000 24600 137100 24700
rect 137000 34100 137100 34200
rect 137000 34200 137100 34300
rect 137000 34300 137100 34400
rect 137000 34400 137100 34500
rect 137000 34500 137100 34600
rect 137000 34600 137100 34700
rect 137000 34700 137100 34800
rect 137000 34800 137100 34900
rect 137000 34900 137100 35000
rect 137000 35000 137100 35100
rect 137000 35100 137100 35200
rect 137000 35200 137100 35300
rect 137000 35300 137100 35400
rect 137000 35400 137100 35500
rect 137000 35500 137100 35600
rect 137000 35600 137100 35700
rect 137000 35700 137100 35800
rect 137000 35800 137100 35900
rect 137000 35900 137100 36000
rect 137000 36000 137100 36100
rect 137000 36100 137100 36200
rect 137000 36200 137100 36300
rect 137000 36300 137100 36400
rect 137000 36400 137100 36500
rect 137000 36500 137100 36600
rect 137000 36600 137100 36700
rect 137000 36700 137100 36800
rect 137000 36800 137100 36900
rect 137000 36900 137100 37000
rect 137000 37000 137100 37100
rect 137100 22200 137200 22300
rect 137100 22300 137200 22400
rect 137100 22400 137200 22500
rect 137100 22500 137200 22600
rect 137100 22600 137200 22700
rect 137100 22700 137200 22800
rect 137100 22800 137200 22900
rect 137100 22900 137200 23000
rect 137100 23000 137200 23100
rect 137100 23100 137200 23200
rect 137100 23200 137200 23300
rect 137100 23300 137200 23400
rect 137100 23400 137200 23500
rect 137100 23500 137200 23600
rect 137100 23600 137200 23700
rect 137100 23700 137200 23800
rect 137100 23800 137200 23900
rect 137100 23900 137200 24000
rect 137100 24000 137200 24100
rect 137100 24100 137200 24200
rect 137100 24200 137200 24300
rect 137100 24300 137200 24400
rect 137100 24400 137200 24500
rect 137100 24500 137200 24600
rect 137100 34300 137200 34400
rect 137100 34400 137200 34500
rect 137100 34500 137200 34600
rect 137100 34600 137200 34700
rect 137100 34700 137200 34800
rect 137100 34800 137200 34900
rect 137100 34900 137200 35000
rect 137100 35000 137200 35100
rect 137100 35100 137200 35200
rect 137100 35200 137200 35300
rect 137100 35300 137200 35400
rect 137100 35400 137200 35500
rect 137100 35500 137200 35600
rect 137100 35600 137200 35700
rect 137100 35700 137200 35800
rect 137100 35800 137200 35900
rect 137100 35900 137200 36000
rect 137100 36000 137200 36100
rect 137100 36100 137200 36200
rect 137100 36200 137200 36300
rect 137100 36300 137200 36400
rect 137100 36400 137200 36500
rect 137100 36500 137200 36600
rect 137100 36600 137200 36700
rect 137100 36700 137200 36800
rect 137100 36800 137200 36900
rect 137100 36900 137200 37000
rect 137100 37000 137200 37100
rect 137100 37100 137200 37200
rect 137200 22100 137300 22200
rect 137200 22200 137300 22300
rect 137200 22300 137300 22400
rect 137200 22400 137300 22500
rect 137200 22500 137300 22600
rect 137200 22600 137300 22700
rect 137200 22700 137300 22800
rect 137200 22800 137300 22900
rect 137200 22900 137300 23000
rect 137200 23000 137300 23100
rect 137200 23100 137300 23200
rect 137200 23200 137300 23300
rect 137200 23300 137300 23400
rect 137200 23400 137300 23500
rect 137200 23500 137300 23600
rect 137200 23600 137300 23700
rect 137200 23700 137300 23800
rect 137200 23800 137300 23900
rect 137200 23900 137300 24000
rect 137200 24000 137300 24100
rect 137200 24100 137300 24200
rect 137200 24200 137300 24300
rect 137200 24300 137300 24400
rect 137200 24400 137300 24500
rect 137200 24500 137300 24600
rect 137200 34400 137300 34500
rect 137200 34500 137300 34600
rect 137200 34600 137300 34700
rect 137200 34700 137300 34800
rect 137200 34800 137300 34900
rect 137200 34900 137300 35000
rect 137200 35000 137300 35100
rect 137200 35100 137300 35200
rect 137200 35200 137300 35300
rect 137200 35300 137300 35400
rect 137200 35400 137300 35500
rect 137200 35500 137300 35600
rect 137200 35600 137300 35700
rect 137200 35700 137300 35800
rect 137200 35800 137300 35900
rect 137200 35900 137300 36000
rect 137200 36000 137300 36100
rect 137200 36100 137300 36200
rect 137200 36200 137300 36300
rect 137200 36300 137300 36400
rect 137200 36400 137300 36500
rect 137200 36500 137300 36600
rect 137200 36600 137300 36700
rect 137200 36700 137300 36800
rect 137200 36800 137300 36900
rect 137200 36900 137300 37000
rect 137200 37000 137300 37100
rect 137200 37100 137300 37200
rect 137200 37200 137300 37300
rect 137300 22100 137400 22200
rect 137300 22200 137400 22300
rect 137300 22300 137400 22400
rect 137300 22400 137400 22500
rect 137300 22500 137400 22600
rect 137300 22600 137400 22700
rect 137300 22700 137400 22800
rect 137300 22800 137400 22900
rect 137300 22900 137400 23000
rect 137300 23000 137400 23100
rect 137300 23100 137400 23200
rect 137300 23200 137400 23300
rect 137300 23300 137400 23400
rect 137300 23400 137400 23500
rect 137300 23500 137400 23600
rect 137300 23600 137400 23700
rect 137300 23700 137400 23800
rect 137300 23800 137400 23900
rect 137300 23900 137400 24000
rect 137300 24000 137400 24100
rect 137300 24100 137400 24200
rect 137300 24200 137400 24300
rect 137300 24300 137400 24400
rect 137300 24400 137400 24500
rect 137300 34500 137400 34600
rect 137300 34600 137400 34700
rect 137300 34700 137400 34800
rect 137300 34800 137400 34900
rect 137300 34900 137400 35000
rect 137300 35000 137400 35100
rect 137300 35100 137400 35200
rect 137300 35200 137400 35300
rect 137300 35300 137400 35400
rect 137300 35400 137400 35500
rect 137300 35500 137400 35600
rect 137300 35600 137400 35700
rect 137300 35700 137400 35800
rect 137300 35800 137400 35900
rect 137300 35900 137400 36000
rect 137300 36000 137400 36100
rect 137300 36100 137400 36200
rect 137300 36200 137400 36300
rect 137300 36300 137400 36400
rect 137300 36400 137400 36500
rect 137300 36500 137400 36600
rect 137300 36600 137400 36700
rect 137300 36700 137400 36800
rect 137300 36800 137400 36900
rect 137300 36900 137400 37000
rect 137300 37000 137400 37100
rect 137300 37100 137400 37200
rect 137300 37200 137400 37300
rect 137400 22000 137500 22100
rect 137400 22100 137500 22200
rect 137400 22200 137500 22300
rect 137400 22300 137500 22400
rect 137400 22400 137500 22500
rect 137400 22500 137500 22600
rect 137400 22600 137500 22700
rect 137400 22700 137500 22800
rect 137400 22800 137500 22900
rect 137400 22900 137500 23000
rect 137400 23000 137500 23100
rect 137400 23100 137500 23200
rect 137400 23200 137500 23300
rect 137400 23300 137500 23400
rect 137400 23400 137500 23500
rect 137400 23500 137500 23600
rect 137400 23600 137500 23700
rect 137400 23700 137500 23800
rect 137400 23800 137500 23900
rect 137400 23900 137500 24000
rect 137400 24000 137500 24100
rect 137400 24100 137500 24200
rect 137400 24200 137500 24300
rect 137400 24300 137500 24400
rect 137400 34600 137500 34700
rect 137400 34700 137500 34800
rect 137400 34800 137500 34900
rect 137400 34900 137500 35000
rect 137400 35000 137500 35100
rect 137400 35100 137500 35200
rect 137400 35200 137500 35300
rect 137400 35300 137500 35400
rect 137400 35400 137500 35500
rect 137400 35500 137500 35600
rect 137400 35600 137500 35700
rect 137400 35700 137500 35800
rect 137400 35800 137500 35900
rect 137400 35900 137500 36000
rect 137400 36000 137500 36100
rect 137400 36100 137500 36200
rect 137400 36200 137500 36300
rect 137400 36300 137500 36400
rect 137400 36400 137500 36500
rect 137400 36500 137500 36600
rect 137400 36600 137500 36700
rect 137400 36700 137500 36800
rect 137400 36800 137500 36900
rect 137400 36900 137500 37000
rect 137400 37000 137500 37100
rect 137400 37100 137500 37200
rect 137400 37200 137500 37300
rect 137400 37300 137500 37400
rect 137500 22000 137600 22100
rect 137500 22100 137600 22200
rect 137500 22200 137600 22300
rect 137500 22300 137600 22400
rect 137500 22400 137600 22500
rect 137500 22500 137600 22600
rect 137500 22600 137600 22700
rect 137500 22700 137600 22800
rect 137500 22800 137600 22900
rect 137500 22900 137600 23000
rect 137500 23000 137600 23100
rect 137500 23100 137600 23200
rect 137500 23200 137600 23300
rect 137500 23300 137600 23400
rect 137500 23400 137600 23500
rect 137500 23500 137600 23600
rect 137500 23600 137600 23700
rect 137500 23700 137600 23800
rect 137500 23800 137600 23900
rect 137500 23900 137600 24000
rect 137500 24000 137600 24100
rect 137500 24100 137600 24200
rect 137500 24200 137600 24300
rect 137500 24300 137600 24400
rect 137500 34800 137600 34900
rect 137500 34900 137600 35000
rect 137500 35000 137600 35100
rect 137500 35100 137600 35200
rect 137500 35200 137600 35300
rect 137500 35300 137600 35400
rect 137500 35400 137600 35500
rect 137500 35500 137600 35600
rect 137500 35600 137600 35700
rect 137500 35700 137600 35800
rect 137500 35800 137600 35900
rect 137500 35900 137600 36000
rect 137500 36000 137600 36100
rect 137500 36100 137600 36200
rect 137500 36200 137600 36300
rect 137500 36300 137600 36400
rect 137500 36400 137600 36500
rect 137500 36500 137600 36600
rect 137500 36600 137600 36700
rect 137500 36700 137600 36800
rect 137500 36800 137600 36900
rect 137500 36900 137600 37000
rect 137500 37000 137600 37100
rect 137500 37100 137600 37200
rect 137500 37200 137600 37300
rect 137500 37300 137600 37400
rect 137600 22000 137700 22100
rect 137600 22100 137700 22200
rect 137600 22200 137700 22300
rect 137600 22300 137700 22400
rect 137600 22400 137700 22500
rect 137600 22500 137700 22600
rect 137600 22600 137700 22700
rect 137600 22700 137700 22800
rect 137600 22800 137700 22900
rect 137600 22900 137700 23000
rect 137600 23000 137700 23100
rect 137600 23100 137700 23200
rect 137600 23200 137700 23300
rect 137600 23300 137700 23400
rect 137600 23400 137700 23500
rect 137600 23500 137700 23600
rect 137600 23600 137700 23700
rect 137600 23700 137700 23800
rect 137600 23800 137700 23900
rect 137600 23900 137700 24000
rect 137600 24000 137700 24100
rect 137600 24100 137700 24200
rect 137600 24200 137700 24300
rect 137600 34800 137700 34900
rect 137600 34900 137700 35000
rect 137600 35000 137700 35100
rect 137600 35100 137700 35200
rect 137600 35200 137700 35300
rect 137600 35300 137700 35400
rect 137600 35400 137700 35500
rect 137600 35500 137700 35600
rect 137600 35600 137700 35700
rect 137600 35700 137700 35800
rect 137600 35800 137700 35900
rect 137600 35900 137700 36000
rect 137600 36000 137700 36100
rect 137600 36100 137700 36200
rect 137600 36200 137700 36300
rect 137600 36300 137700 36400
rect 137600 36400 137700 36500
rect 137600 36500 137700 36600
rect 137600 36600 137700 36700
rect 137600 36700 137700 36800
rect 137600 36800 137700 36900
rect 137600 36900 137700 37000
rect 137600 37000 137700 37100
rect 137600 37100 137700 37200
rect 137600 37200 137700 37300
rect 137600 37300 137700 37400
rect 137600 37400 137700 37500
rect 137700 21900 137800 22000
rect 137700 22000 137800 22100
rect 137700 22100 137800 22200
rect 137700 22200 137800 22300
rect 137700 22300 137800 22400
rect 137700 22400 137800 22500
rect 137700 22500 137800 22600
rect 137700 22600 137800 22700
rect 137700 22700 137800 22800
rect 137700 22800 137800 22900
rect 137700 22900 137800 23000
rect 137700 23000 137800 23100
rect 137700 23100 137800 23200
rect 137700 23200 137800 23300
rect 137700 23300 137800 23400
rect 137700 23400 137800 23500
rect 137700 23500 137800 23600
rect 137700 23600 137800 23700
rect 137700 23700 137800 23800
rect 137700 23800 137800 23900
rect 137700 23900 137800 24000
rect 137700 24000 137800 24100
rect 137700 24100 137800 24200
rect 137700 24200 137800 24300
rect 137700 35000 137800 35100
rect 137700 35100 137800 35200
rect 137700 35200 137800 35300
rect 137700 35300 137800 35400
rect 137700 35400 137800 35500
rect 137700 35500 137800 35600
rect 137700 35600 137800 35700
rect 137700 35700 137800 35800
rect 137700 35800 137800 35900
rect 137700 35900 137800 36000
rect 137700 36000 137800 36100
rect 137700 36100 137800 36200
rect 137700 36200 137800 36300
rect 137700 36300 137800 36400
rect 137700 36400 137800 36500
rect 137700 36500 137800 36600
rect 137700 36600 137800 36700
rect 137700 36700 137800 36800
rect 137700 36800 137800 36900
rect 137700 36900 137800 37000
rect 137700 37000 137800 37100
rect 137700 37100 137800 37200
rect 137700 37200 137800 37300
rect 137700 37300 137800 37400
rect 137700 37400 137800 37500
rect 137700 37500 137800 37600
rect 137800 21900 137900 22000
rect 137800 22000 137900 22100
rect 137800 22100 137900 22200
rect 137800 22200 137900 22300
rect 137800 22300 137900 22400
rect 137800 22400 137900 22500
rect 137800 22500 137900 22600
rect 137800 22600 137900 22700
rect 137800 22700 137900 22800
rect 137800 22800 137900 22900
rect 137800 22900 137900 23000
rect 137800 23000 137900 23100
rect 137800 23100 137900 23200
rect 137800 23200 137900 23300
rect 137800 23300 137900 23400
rect 137800 23400 137900 23500
rect 137800 23500 137900 23600
rect 137800 23600 137900 23700
rect 137800 23700 137900 23800
rect 137800 23800 137900 23900
rect 137800 23900 137900 24000
rect 137800 24000 137900 24100
rect 137800 24100 137900 24200
rect 137800 35000 137900 35100
rect 137800 35100 137900 35200
rect 137800 35200 137900 35300
rect 137800 35300 137900 35400
rect 137800 35400 137900 35500
rect 137800 35500 137900 35600
rect 137800 35600 137900 35700
rect 137800 35700 137900 35800
rect 137800 35800 137900 35900
rect 137800 35900 137900 36000
rect 137800 36000 137900 36100
rect 137800 36100 137900 36200
rect 137800 36200 137900 36300
rect 137800 36300 137900 36400
rect 137800 36400 137900 36500
rect 137800 36500 137900 36600
rect 137800 36600 137900 36700
rect 137800 36700 137900 36800
rect 137800 36800 137900 36900
rect 137800 36900 137900 37000
rect 137800 37000 137900 37100
rect 137800 37100 137900 37200
rect 137800 37200 137900 37300
rect 137800 37300 137900 37400
rect 137800 37400 137900 37500
rect 137800 37500 137900 37600
rect 137900 21900 138000 22000
rect 137900 22000 138000 22100
rect 137900 22100 138000 22200
rect 137900 22200 138000 22300
rect 137900 22300 138000 22400
rect 137900 22400 138000 22500
rect 137900 22500 138000 22600
rect 137900 22600 138000 22700
rect 137900 22700 138000 22800
rect 137900 22800 138000 22900
rect 137900 22900 138000 23000
rect 137900 23000 138000 23100
rect 137900 23100 138000 23200
rect 137900 23200 138000 23300
rect 137900 23300 138000 23400
rect 137900 23400 138000 23500
rect 137900 23500 138000 23600
rect 137900 23600 138000 23700
rect 137900 23700 138000 23800
rect 137900 23800 138000 23900
rect 137900 23900 138000 24000
rect 137900 24000 138000 24100
rect 137900 24100 138000 24200
rect 137900 35100 138000 35200
rect 137900 35200 138000 35300
rect 137900 35300 138000 35400
rect 137900 35400 138000 35500
rect 137900 35500 138000 35600
rect 137900 35600 138000 35700
rect 137900 35700 138000 35800
rect 137900 35800 138000 35900
rect 137900 35900 138000 36000
rect 137900 36000 138000 36100
rect 137900 36100 138000 36200
rect 137900 36200 138000 36300
rect 137900 36300 138000 36400
rect 137900 36400 138000 36500
rect 137900 36500 138000 36600
rect 137900 36600 138000 36700
rect 137900 36700 138000 36800
rect 137900 36800 138000 36900
rect 137900 36900 138000 37000
rect 137900 37000 138000 37100
rect 137900 37100 138000 37200
rect 137900 37200 138000 37300
rect 137900 37300 138000 37400
rect 137900 37400 138000 37500
rect 137900 37500 138000 37600
rect 137900 37600 138000 37700
rect 138000 21800 138100 21900
rect 138000 21900 138100 22000
rect 138000 22000 138100 22100
rect 138000 22100 138100 22200
rect 138000 22200 138100 22300
rect 138000 22300 138100 22400
rect 138000 22400 138100 22500
rect 138000 22500 138100 22600
rect 138000 22600 138100 22700
rect 138000 22700 138100 22800
rect 138000 22800 138100 22900
rect 138000 22900 138100 23000
rect 138000 23000 138100 23100
rect 138000 23100 138100 23200
rect 138000 23200 138100 23300
rect 138000 23300 138100 23400
rect 138000 23400 138100 23500
rect 138000 23500 138100 23600
rect 138000 23600 138100 23700
rect 138000 23700 138100 23800
rect 138000 23800 138100 23900
rect 138000 23900 138100 24000
rect 138000 24000 138100 24100
rect 138000 35200 138100 35300
rect 138000 35300 138100 35400
rect 138000 35400 138100 35500
rect 138000 35500 138100 35600
rect 138000 35600 138100 35700
rect 138000 35700 138100 35800
rect 138000 35800 138100 35900
rect 138000 35900 138100 36000
rect 138000 36000 138100 36100
rect 138000 36100 138100 36200
rect 138000 36200 138100 36300
rect 138000 36300 138100 36400
rect 138000 36400 138100 36500
rect 138000 36500 138100 36600
rect 138000 36600 138100 36700
rect 138000 36700 138100 36800
rect 138000 36800 138100 36900
rect 138000 36900 138100 37000
rect 138000 37000 138100 37100
rect 138000 37100 138100 37200
rect 138000 37200 138100 37300
rect 138000 37300 138100 37400
rect 138000 37400 138100 37500
rect 138000 37500 138100 37600
rect 138000 37600 138100 37700
rect 138100 21800 138200 21900
rect 138100 21900 138200 22000
rect 138100 22000 138200 22100
rect 138100 22100 138200 22200
rect 138100 22200 138200 22300
rect 138100 22300 138200 22400
rect 138100 22400 138200 22500
rect 138100 22500 138200 22600
rect 138100 22600 138200 22700
rect 138100 22700 138200 22800
rect 138100 22800 138200 22900
rect 138100 22900 138200 23000
rect 138100 23000 138200 23100
rect 138100 23100 138200 23200
rect 138100 23200 138200 23300
rect 138100 23300 138200 23400
rect 138100 23400 138200 23500
rect 138100 23500 138200 23600
rect 138100 23600 138200 23700
rect 138100 23700 138200 23800
rect 138100 23800 138200 23900
rect 138100 23900 138200 24000
rect 138100 24000 138200 24100
rect 138100 35300 138200 35400
rect 138100 35400 138200 35500
rect 138100 35500 138200 35600
rect 138100 35600 138200 35700
rect 138100 35700 138200 35800
rect 138100 35800 138200 35900
rect 138100 35900 138200 36000
rect 138100 36000 138200 36100
rect 138100 36100 138200 36200
rect 138100 36200 138200 36300
rect 138100 36300 138200 36400
rect 138100 36400 138200 36500
rect 138100 36500 138200 36600
rect 138100 36600 138200 36700
rect 138100 36700 138200 36800
rect 138100 36800 138200 36900
rect 138100 36900 138200 37000
rect 138100 37000 138200 37100
rect 138100 37100 138200 37200
rect 138100 37200 138200 37300
rect 138100 37300 138200 37400
rect 138100 37400 138200 37500
rect 138100 37500 138200 37600
rect 138100 37600 138200 37700
rect 138100 37700 138200 37800
rect 138200 21800 138300 21900
rect 138200 21900 138300 22000
rect 138200 22000 138300 22100
rect 138200 22100 138300 22200
rect 138200 22200 138300 22300
rect 138200 22300 138300 22400
rect 138200 22400 138300 22500
rect 138200 22500 138300 22600
rect 138200 22600 138300 22700
rect 138200 22700 138300 22800
rect 138200 22800 138300 22900
rect 138200 22900 138300 23000
rect 138200 23000 138300 23100
rect 138200 23100 138300 23200
rect 138200 23200 138300 23300
rect 138200 23300 138300 23400
rect 138200 23400 138300 23500
rect 138200 23500 138300 23600
rect 138200 23600 138300 23700
rect 138200 23700 138300 23800
rect 138200 23800 138300 23900
rect 138200 23900 138300 24000
rect 138200 35400 138300 35500
rect 138200 35500 138300 35600
rect 138200 35600 138300 35700
rect 138200 35700 138300 35800
rect 138200 35800 138300 35900
rect 138200 35900 138300 36000
rect 138200 36000 138300 36100
rect 138200 36100 138300 36200
rect 138200 36200 138300 36300
rect 138200 36300 138300 36400
rect 138200 36400 138300 36500
rect 138200 36500 138300 36600
rect 138200 36600 138300 36700
rect 138200 36700 138300 36800
rect 138200 36800 138300 36900
rect 138200 36900 138300 37000
rect 138200 37000 138300 37100
rect 138200 37100 138300 37200
rect 138200 37200 138300 37300
rect 138200 37300 138300 37400
rect 138200 37400 138300 37500
rect 138200 37500 138300 37600
rect 138200 37600 138300 37700
rect 138200 37700 138300 37800
rect 138300 21700 138400 21800
rect 138300 21800 138400 21900
rect 138300 21900 138400 22000
rect 138300 22000 138400 22100
rect 138300 22100 138400 22200
rect 138300 22200 138400 22300
rect 138300 22300 138400 22400
rect 138300 22400 138400 22500
rect 138300 22500 138400 22600
rect 138300 22600 138400 22700
rect 138300 22700 138400 22800
rect 138300 22800 138400 22900
rect 138300 22900 138400 23000
rect 138300 23000 138400 23100
rect 138300 23100 138400 23200
rect 138300 23200 138400 23300
rect 138300 23300 138400 23400
rect 138300 23400 138400 23500
rect 138300 23500 138400 23600
rect 138300 23600 138400 23700
rect 138300 23700 138400 23800
rect 138300 23800 138400 23900
rect 138300 23900 138400 24000
rect 138300 35400 138400 35500
rect 138300 35500 138400 35600
rect 138300 35600 138400 35700
rect 138300 35700 138400 35800
rect 138300 35800 138400 35900
rect 138300 35900 138400 36000
rect 138300 36000 138400 36100
rect 138300 36100 138400 36200
rect 138300 36200 138400 36300
rect 138300 36300 138400 36400
rect 138300 36400 138400 36500
rect 138300 36500 138400 36600
rect 138300 36600 138400 36700
rect 138300 36700 138400 36800
rect 138300 36800 138400 36900
rect 138300 36900 138400 37000
rect 138300 37000 138400 37100
rect 138300 37100 138400 37200
rect 138300 37200 138400 37300
rect 138300 37300 138400 37400
rect 138300 37400 138400 37500
rect 138300 37500 138400 37600
rect 138300 37600 138400 37700
rect 138300 37700 138400 37800
rect 138400 21700 138500 21800
rect 138400 21800 138500 21900
rect 138400 21900 138500 22000
rect 138400 22000 138500 22100
rect 138400 22100 138500 22200
rect 138400 22200 138500 22300
rect 138400 22300 138500 22400
rect 138400 22400 138500 22500
rect 138400 22500 138500 22600
rect 138400 22600 138500 22700
rect 138400 22700 138500 22800
rect 138400 22800 138500 22900
rect 138400 22900 138500 23000
rect 138400 23000 138500 23100
rect 138400 23100 138500 23200
rect 138400 23200 138500 23300
rect 138400 23300 138500 23400
rect 138400 23400 138500 23500
rect 138400 23500 138500 23600
rect 138400 23600 138500 23700
rect 138400 23700 138500 23800
rect 138400 23800 138500 23900
rect 138400 23900 138500 24000
rect 138400 35500 138500 35600
rect 138400 35600 138500 35700
rect 138400 35700 138500 35800
rect 138400 35800 138500 35900
rect 138400 35900 138500 36000
rect 138400 36000 138500 36100
rect 138400 36100 138500 36200
rect 138400 36200 138500 36300
rect 138400 36300 138500 36400
rect 138400 36400 138500 36500
rect 138400 36500 138500 36600
rect 138400 36600 138500 36700
rect 138400 36700 138500 36800
rect 138400 36800 138500 36900
rect 138400 36900 138500 37000
rect 138400 37000 138500 37100
rect 138400 37100 138500 37200
rect 138400 37200 138500 37300
rect 138400 37300 138500 37400
rect 138400 37400 138500 37500
rect 138400 37500 138500 37600
rect 138400 37600 138500 37700
rect 138400 37700 138500 37800
rect 138400 37800 138500 37900
rect 138500 21700 138600 21800
rect 138500 21800 138600 21900
rect 138500 21900 138600 22000
rect 138500 22000 138600 22100
rect 138500 22100 138600 22200
rect 138500 22200 138600 22300
rect 138500 22300 138600 22400
rect 138500 22400 138600 22500
rect 138500 22500 138600 22600
rect 138500 22600 138600 22700
rect 138500 22700 138600 22800
rect 138500 22800 138600 22900
rect 138500 22900 138600 23000
rect 138500 23000 138600 23100
rect 138500 23100 138600 23200
rect 138500 23200 138600 23300
rect 138500 23300 138600 23400
rect 138500 23400 138600 23500
rect 138500 23500 138600 23600
rect 138500 23600 138600 23700
rect 138500 23700 138600 23800
rect 138500 23800 138600 23900
rect 138500 35500 138600 35600
rect 138500 35600 138600 35700
rect 138500 35700 138600 35800
rect 138500 35800 138600 35900
rect 138500 35900 138600 36000
rect 138500 36000 138600 36100
rect 138500 36100 138600 36200
rect 138500 36200 138600 36300
rect 138500 36300 138600 36400
rect 138500 36400 138600 36500
rect 138500 36500 138600 36600
rect 138500 36600 138600 36700
rect 138500 36700 138600 36800
rect 138500 36800 138600 36900
rect 138500 36900 138600 37000
rect 138500 37000 138600 37100
rect 138500 37100 138600 37200
rect 138500 37200 138600 37300
rect 138500 37300 138600 37400
rect 138500 37400 138600 37500
rect 138500 37500 138600 37600
rect 138500 37600 138600 37700
rect 138500 37700 138600 37800
rect 138500 37800 138600 37900
rect 138600 21700 138700 21800
rect 138600 21800 138700 21900
rect 138600 21900 138700 22000
rect 138600 22000 138700 22100
rect 138600 22100 138700 22200
rect 138600 22200 138700 22300
rect 138600 22300 138700 22400
rect 138600 22400 138700 22500
rect 138600 22500 138700 22600
rect 138600 22600 138700 22700
rect 138600 22700 138700 22800
rect 138600 22800 138700 22900
rect 138600 22900 138700 23000
rect 138600 23000 138700 23100
rect 138600 23100 138700 23200
rect 138600 23200 138700 23300
rect 138600 23300 138700 23400
rect 138600 23400 138700 23500
rect 138600 23500 138700 23600
rect 138600 23600 138700 23700
rect 138600 23700 138700 23800
rect 138600 23800 138700 23900
rect 138600 35600 138700 35700
rect 138600 35700 138700 35800
rect 138600 35800 138700 35900
rect 138600 35900 138700 36000
rect 138600 36000 138700 36100
rect 138600 36100 138700 36200
rect 138600 36200 138700 36300
rect 138600 36300 138700 36400
rect 138600 36400 138700 36500
rect 138600 36500 138700 36600
rect 138600 36600 138700 36700
rect 138600 36700 138700 36800
rect 138600 36800 138700 36900
rect 138600 36900 138700 37000
rect 138600 37000 138700 37100
rect 138600 37100 138700 37200
rect 138600 37200 138700 37300
rect 138600 37300 138700 37400
rect 138600 37400 138700 37500
rect 138600 37500 138700 37600
rect 138600 37600 138700 37700
rect 138600 37700 138700 37800
rect 138600 37800 138700 37900
rect 138700 21700 138800 21800
rect 138700 21800 138800 21900
rect 138700 21900 138800 22000
rect 138700 22000 138800 22100
rect 138700 22100 138800 22200
rect 138700 22200 138800 22300
rect 138700 22300 138800 22400
rect 138700 22400 138800 22500
rect 138700 22500 138800 22600
rect 138700 22600 138800 22700
rect 138700 22700 138800 22800
rect 138700 22800 138800 22900
rect 138700 22900 138800 23000
rect 138700 23000 138800 23100
rect 138700 23100 138800 23200
rect 138700 23200 138800 23300
rect 138700 23300 138800 23400
rect 138700 23400 138800 23500
rect 138700 23500 138800 23600
rect 138700 23600 138800 23700
rect 138700 23700 138800 23800
rect 138700 23800 138800 23900
rect 138700 35600 138800 35700
rect 138700 35700 138800 35800
rect 138700 35800 138800 35900
rect 138700 35900 138800 36000
rect 138700 36000 138800 36100
rect 138700 36100 138800 36200
rect 138700 36200 138800 36300
rect 138700 36300 138800 36400
rect 138700 36400 138800 36500
rect 138700 36500 138800 36600
rect 138700 36600 138800 36700
rect 138700 36700 138800 36800
rect 138700 36800 138800 36900
rect 138700 36900 138800 37000
rect 138700 37000 138800 37100
rect 138700 37100 138800 37200
rect 138700 37200 138800 37300
rect 138700 37300 138800 37400
rect 138700 37400 138800 37500
rect 138700 37500 138800 37600
rect 138700 37600 138800 37700
rect 138700 37700 138800 37800
rect 138700 37800 138800 37900
rect 138700 37900 138800 38000
rect 138800 21700 138900 21800
rect 138800 21800 138900 21900
rect 138800 21900 138900 22000
rect 138800 22000 138900 22100
rect 138800 22100 138900 22200
rect 138800 22200 138900 22300
rect 138800 22300 138900 22400
rect 138800 22400 138900 22500
rect 138800 22500 138900 22600
rect 138800 22600 138900 22700
rect 138800 22700 138900 22800
rect 138800 22800 138900 22900
rect 138800 22900 138900 23000
rect 138800 23000 138900 23100
rect 138800 23100 138900 23200
rect 138800 23200 138900 23300
rect 138800 23300 138900 23400
rect 138800 23400 138900 23500
rect 138800 23500 138900 23600
rect 138800 23600 138900 23700
rect 138800 23700 138900 23800
rect 138800 23800 138900 23900
rect 138800 35700 138900 35800
rect 138800 35800 138900 35900
rect 138800 35900 138900 36000
rect 138800 36000 138900 36100
rect 138800 36100 138900 36200
rect 138800 36200 138900 36300
rect 138800 36300 138900 36400
rect 138800 36400 138900 36500
rect 138800 36500 138900 36600
rect 138800 36600 138900 36700
rect 138800 36700 138900 36800
rect 138800 36800 138900 36900
rect 138800 36900 138900 37000
rect 138800 37000 138900 37100
rect 138800 37100 138900 37200
rect 138800 37200 138900 37300
rect 138800 37300 138900 37400
rect 138800 37400 138900 37500
rect 138800 37500 138900 37600
rect 138800 37600 138900 37700
rect 138800 37700 138900 37800
rect 138800 37800 138900 37900
rect 138800 37900 138900 38000
rect 138900 21600 139000 21700
rect 138900 21700 139000 21800
rect 138900 21800 139000 21900
rect 138900 21900 139000 22000
rect 138900 22000 139000 22100
rect 138900 22100 139000 22200
rect 138900 22200 139000 22300
rect 138900 22300 139000 22400
rect 138900 22400 139000 22500
rect 138900 22500 139000 22600
rect 138900 22600 139000 22700
rect 138900 22700 139000 22800
rect 138900 22800 139000 22900
rect 138900 22900 139000 23000
rect 138900 23000 139000 23100
rect 138900 23100 139000 23200
rect 138900 23200 139000 23300
rect 138900 23300 139000 23400
rect 138900 23400 139000 23500
rect 138900 23500 139000 23600
rect 138900 23600 139000 23700
rect 138900 23700 139000 23800
rect 138900 35700 139000 35800
rect 138900 35800 139000 35900
rect 138900 35900 139000 36000
rect 138900 36000 139000 36100
rect 138900 36100 139000 36200
rect 138900 36200 139000 36300
rect 138900 36300 139000 36400
rect 138900 36400 139000 36500
rect 138900 36500 139000 36600
rect 138900 36600 139000 36700
rect 138900 36700 139000 36800
rect 138900 36800 139000 36900
rect 138900 36900 139000 37000
rect 138900 37000 139000 37100
rect 138900 37100 139000 37200
rect 138900 37200 139000 37300
rect 138900 37300 139000 37400
rect 138900 37400 139000 37500
rect 138900 37500 139000 37600
rect 138900 37600 139000 37700
rect 138900 37700 139000 37800
rect 138900 37800 139000 37900
rect 138900 37900 139000 38000
rect 139000 21600 139100 21700
rect 139000 21700 139100 21800
rect 139000 21800 139100 21900
rect 139000 21900 139100 22000
rect 139000 22000 139100 22100
rect 139000 22100 139100 22200
rect 139000 22200 139100 22300
rect 139000 22300 139100 22400
rect 139000 22400 139100 22500
rect 139000 22500 139100 22600
rect 139000 22600 139100 22700
rect 139000 22700 139100 22800
rect 139000 22800 139100 22900
rect 139000 22900 139100 23000
rect 139000 23000 139100 23100
rect 139000 23100 139100 23200
rect 139000 23200 139100 23300
rect 139000 23300 139100 23400
rect 139000 23400 139100 23500
rect 139000 23500 139100 23600
rect 139000 23600 139100 23700
rect 139000 23700 139100 23800
rect 139000 35800 139100 35900
rect 139000 35900 139100 36000
rect 139000 36000 139100 36100
rect 139000 36100 139100 36200
rect 139000 36200 139100 36300
rect 139000 36300 139100 36400
rect 139000 36400 139100 36500
rect 139000 36500 139100 36600
rect 139000 36600 139100 36700
rect 139000 36700 139100 36800
rect 139000 36800 139100 36900
rect 139000 36900 139100 37000
rect 139000 37000 139100 37100
rect 139000 37100 139100 37200
rect 139000 37200 139100 37300
rect 139000 37300 139100 37400
rect 139000 37400 139100 37500
rect 139000 37500 139100 37600
rect 139000 37600 139100 37700
rect 139000 37700 139100 37800
rect 139000 37800 139100 37900
rect 139000 37900 139100 38000
rect 139000 38000 139100 38100
rect 139100 21600 139200 21700
rect 139100 21700 139200 21800
rect 139100 21800 139200 21900
rect 139100 21900 139200 22000
rect 139100 22000 139200 22100
rect 139100 22100 139200 22200
rect 139100 22200 139200 22300
rect 139100 22300 139200 22400
rect 139100 22400 139200 22500
rect 139100 22500 139200 22600
rect 139100 22600 139200 22700
rect 139100 22700 139200 22800
rect 139100 22800 139200 22900
rect 139100 22900 139200 23000
rect 139100 23000 139200 23100
rect 139100 23100 139200 23200
rect 139100 23200 139200 23300
rect 139100 23300 139200 23400
rect 139100 23400 139200 23500
rect 139100 23500 139200 23600
rect 139100 23600 139200 23700
rect 139100 23700 139200 23800
rect 139100 35800 139200 35900
rect 139100 35900 139200 36000
rect 139100 36000 139200 36100
rect 139100 36100 139200 36200
rect 139100 36200 139200 36300
rect 139100 36300 139200 36400
rect 139100 36400 139200 36500
rect 139100 36500 139200 36600
rect 139100 36600 139200 36700
rect 139100 36700 139200 36800
rect 139100 36800 139200 36900
rect 139100 36900 139200 37000
rect 139100 37000 139200 37100
rect 139100 37100 139200 37200
rect 139100 37200 139200 37300
rect 139100 37300 139200 37400
rect 139100 37400 139200 37500
rect 139100 37500 139200 37600
rect 139100 37600 139200 37700
rect 139100 37700 139200 37800
rect 139100 37800 139200 37900
rect 139100 37900 139200 38000
rect 139100 38000 139200 38100
rect 139200 21600 139300 21700
rect 139200 21700 139300 21800
rect 139200 21800 139300 21900
rect 139200 21900 139300 22000
rect 139200 22000 139300 22100
rect 139200 22100 139300 22200
rect 139200 22200 139300 22300
rect 139200 22300 139300 22400
rect 139200 22400 139300 22500
rect 139200 22500 139300 22600
rect 139200 22600 139300 22700
rect 139200 22700 139300 22800
rect 139200 22800 139300 22900
rect 139200 22900 139300 23000
rect 139200 23000 139300 23100
rect 139200 23100 139300 23200
rect 139200 23200 139300 23300
rect 139200 23300 139300 23400
rect 139200 23400 139300 23500
rect 139200 23500 139300 23600
rect 139200 23600 139300 23700
rect 139200 23700 139300 23800
rect 139200 35900 139300 36000
rect 139200 36000 139300 36100
rect 139200 36100 139300 36200
rect 139200 36200 139300 36300
rect 139200 36300 139300 36400
rect 139200 36400 139300 36500
rect 139200 36500 139300 36600
rect 139200 36600 139300 36700
rect 139200 36700 139300 36800
rect 139200 36800 139300 36900
rect 139200 36900 139300 37000
rect 139200 37000 139300 37100
rect 139200 37100 139300 37200
rect 139200 37200 139300 37300
rect 139200 37300 139300 37400
rect 139200 37400 139300 37500
rect 139200 37500 139300 37600
rect 139200 37600 139300 37700
rect 139200 37700 139300 37800
rect 139200 37800 139300 37900
rect 139200 37900 139300 38000
rect 139200 38000 139300 38100
rect 139300 21600 139400 21700
rect 139300 21700 139400 21800
rect 139300 21800 139400 21900
rect 139300 21900 139400 22000
rect 139300 22000 139400 22100
rect 139300 22100 139400 22200
rect 139300 22200 139400 22300
rect 139300 22300 139400 22400
rect 139300 22400 139400 22500
rect 139300 22500 139400 22600
rect 139300 22600 139400 22700
rect 139300 22700 139400 22800
rect 139300 22800 139400 22900
rect 139300 22900 139400 23000
rect 139300 23000 139400 23100
rect 139300 23100 139400 23200
rect 139300 23200 139400 23300
rect 139300 23300 139400 23400
rect 139300 23400 139400 23500
rect 139300 23500 139400 23600
rect 139300 23600 139400 23700
rect 139300 23700 139400 23800
rect 139300 35900 139400 36000
rect 139300 36000 139400 36100
rect 139300 36100 139400 36200
rect 139300 36200 139400 36300
rect 139300 36300 139400 36400
rect 139300 36400 139400 36500
rect 139300 36500 139400 36600
rect 139300 36600 139400 36700
rect 139300 36700 139400 36800
rect 139300 36800 139400 36900
rect 139300 36900 139400 37000
rect 139300 37000 139400 37100
rect 139300 37100 139400 37200
rect 139300 37200 139400 37300
rect 139300 37300 139400 37400
rect 139300 37400 139400 37500
rect 139300 37500 139400 37600
rect 139300 37600 139400 37700
rect 139300 37700 139400 37800
rect 139300 37800 139400 37900
rect 139300 37900 139400 38000
rect 139300 38000 139400 38100
rect 139400 21600 139500 21700
rect 139400 21700 139500 21800
rect 139400 21800 139500 21900
rect 139400 21900 139500 22000
rect 139400 22000 139500 22100
rect 139400 22100 139500 22200
rect 139400 22200 139500 22300
rect 139400 22300 139500 22400
rect 139400 22400 139500 22500
rect 139400 22500 139500 22600
rect 139400 22600 139500 22700
rect 139400 22700 139500 22800
rect 139400 22800 139500 22900
rect 139400 22900 139500 23000
rect 139400 23000 139500 23100
rect 139400 23100 139500 23200
rect 139400 23200 139500 23300
rect 139400 23300 139500 23400
rect 139400 23400 139500 23500
rect 139400 23500 139500 23600
rect 139400 23600 139500 23700
rect 139400 23700 139500 23800
rect 139400 35900 139500 36000
rect 139400 36000 139500 36100
rect 139400 36100 139500 36200
rect 139400 36200 139500 36300
rect 139400 36300 139500 36400
rect 139400 36400 139500 36500
rect 139400 36500 139500 36600
rect 139400 36600 139500 36700
rect 139400 36700 139500 36800
rect 139400 36800 139500 36900
rect 139400 36900 139500 37000
rect 139400 37000 139500 37100
rect 139400 37100 139500 37200
rect 139400 37200 139500 37300
rect 139400 37300 139500 37400
rect 139400 37400 139500 37500
rect 139400 37500 139500 37600
rect 139400 37600 139500 37700
rect 139400 37700 139500 37800
rect 139400 37800 139500 37900
rect 139400 37900 139500 38000
rect 139400 38000 139500 38100
rect 139400 38100 139500 38200
rect 139500 21600 139600 21700
rect 139500 21700 139600 21800
rect 139500 21800 139600 21900
rect 139500 21900 139600 22000
rect 139500 22000 139600 22100
rect 139500 22100 139600 22200
rect 139500 22200 139600 22300
rect 139500 22300 139600 22400
rect 139500 22400 139600 22500
rect 139500 22500 139600 22600
rect 139500 22600 139600 22700
rect 139500 22700 139600 22800
rect 139500 22800 139600 22900
rect 139500 22900 139600 23000
rect 139500 23000 139600 23100
rect 139500 23100 139600 23200
rect 139500 23200 139600 23300
rect 139500 23300 139600 23400
rect 139500 23400 139600 23500
rect 139500 23500 139600 23600
rect 139500 23600 139600 23700
rect 139500 23700 139600 23800
rect 139500 36000 139600 36100
rect 139500 36100 139600 36200
rect 139500 36200 139600 36300
rect 139500 36300 139600 36400
rect 139500 36400 139600 36500
rect 139500 36500 139600 36600
rect 139500 36600 139600 36700
rect 139500 36700 139600 36800
rect 139500 36800 139600 36900
rect 139500 36900 139600 37000
rect 139500 37000 139600 37100
rect 139500 37100 139600 37200
rect 139500 37200 139600 37300
rect 139500 37300 139600 37400
rect 139500 37400 139600 37500
rect 139500 37500 139600 37600
rect 139500 37600 139600 37700
rect 139500 37700 139600 37800
rect 139500 37800 139600 37900
rect 139500 37900 139600 38000
rect 139500 38000 139600 38100
rect 139500 38100 139600 38200
rect 139600 21600 139700 21700
rect 139600 21700 139700 21800
rect 139600 21800 139700 21900
rect 139600 21900 139700 22000
rect 139600 22000 139700 22100
rect 139600 22100 139700 22200
rect 139600 22200 139700 22300
rect 139600 22300 139700 22400
rect 139600 22400 139700 22500
rect 139600 22500 139700 22600
rect 139600 22600 139700 22700
rect 139600 22700 139700 22800
rect 139600 22800 139700 22900
rect 139600 22900 139700 23000
rect 139600 23000 139700 23100
rect 139600 23100 139700 23200
rect 139600 23200 139700 23300
rect 139600 23300 139700 23400
rect 139600 23400 139700 23500
rect 139600 23500 139700 23600
rect 139600 23600 139700 23700
rect 139600 23700 139700 23800
rect 139600 36000 139700 36100
rect 139600 36100 139700 36200
rect 139600 36200 139700 36300
rect 139600 36300 139700 36400
rect 139600 36400 139700 36500
rect 139600 36500 139700 36600
rect 139600 36600 139700 36700
rect 139600 36700 139700 36800
rect 139600 36800 139700 36900
rect 139600 36900 139700 37000
rect 139600 37000 139700 37100
rect 139600 37100 139700 37200
rect 139600 37200 139700 37300
rect 139600 37300 139700 37400
rect 139600 37400 139700 37500
rect 139600 37500 139700 37600
rect 139600 37600 139700 37700
rect 139600 37700 139700 37800
rect 139600 37800 139700 37900
rect 139600 37900 139700 38000
rect 139600 38000 139700 38100
rect 139600 38100 139700 38200
rect 139700 21600 139800 21700
rect 139700 21700 139800 21800
rect 139700 21800 139800 21900
rect 139700 21900 139800 22000
rect 139700 22000 139800 22100
rect 139700 22100 139800 22200
rect 139700 22200 139800 22300
rect 139700 22300 139800 22400
rect 139700 22400 139800 22500
rect 139700 22500 139800 22600
rect 139700 22600 139800 22700
rect 139700 22700 139800 22800
rect 139700 22800 139800 22900
rect 139700 22900 139800 23000
rect 139700 23000 139800 23100
rect 139700 23100 139800 23200
rect 139700 23200 139800 23300
rect 139700 23300 139800 23400
rect 139700 23400 139800 23500
rect 139700 23500 139800 23600
rect 139700 23600 139800 23700
rect 139700 23700 139800 23800
rect 139700 36000 139800 36100
rect 139700 36100 139800 36200
rect 139700 36200 139800 36300
rect 139700 36300 139800 36400
rect 139700 36400 139800 36500
rect 139700 36500 139800 36600
rect 139700 36600 139800 36700
rect 139700 36700 139800 36800
rect 139700 36800 139800 36900
rect 139700 36900 139800 37000
rect 139700 37000 139800 37100
rect 139700 37100 139800 37200
rect 139700 37200 139800 37300
rect 139700 37300 139800 37400
rect 139700 37400 139800 37500
rect 139700 37500 139800 37600
rect 139700 37600 139800 37700
rect 139700 37700 139800 37800
rect 139700 37800 139800 37900
rect 139700 37900 139800 38000
rect 139700 38000 139800 38100
rect 139700 38100 139800 38200
rect 139800 21600 139900 21700
rect 139800 21700 139900 21800
rect 139800 21800 139900 21900
rect 139800 21900 139900 22000
rect 139800 22000 139900 22100
rect 139800 22100 139900 22200
rect 139800 22200 139900 22300
rect 139800 22300 139900 22400
rect 139800 22400 139900 22500
rect 139800 22500 139900 22600
rect 139800 22600 139900 22700
rect 139800 22700 139900 22800
rect 139800 22800 139900 22900
rect 139800 22900 139900 23000
rect 139800 23000 139900 23100
rect 139800 23100 139900 23200
rect 139800 23200 139900 23300
rect 139800 23300 139900 23400
rect 139800 23400 139900 23500
rect 139800 23500 139900 23600
rect 139800 23600 139900 23700
rect 139800 23700 139900 23800
rect 139800 36000 139900 36100
rect 139800 36100 139900 36200
rect 139800 36200 139900 36300
rect 139800 36300 139900 36400
rect 139800 36400 139900 36500
rect 139800 36500 139900 36600
rect 139800 36600 139900 36700
rect 139800 36700 139900 36800
rect 139800 36800 139900 36900
rect 139800 36900 139900 37000
rect 139800 37000 139900 37100
rect 139800 37100 139900 37200
rect 139800 37200 139900 37300
rect 139800 37300 139900 37400
rect 139800 37400 139900 37500
rect 139800 37500 139900 37600
rect 139800 37600 139900 37700
rect 139800 37700 139900 37800
rect 139800 37800 139900 37900
rect 139800 37900 139900 38000
rect 139800 38000 139900 38100
rect 139800 38100 139900 38200
rect 139900 21600 140000 21700
rect 139900 21700 140000 21800
rect 139900 21800 140000 21900
rect 139900 21900 140000 22000
rect 139900 22000 140000 22100
rect 139900 22100 140000 22200
rect 139900 22200 140000 22300
rect 139900 22300 140000 22400
rect 139900 22400 140000 22500
rect 139900 22500 140000 22600
rect 139900 22600 140000 22700
rect 139900 22700 140000 22800
rect 139900 22800 140000 22900
rect 139900 22900 140000 23000
rect 139900 23000 140000 23100
rect 139900 23100 140000 23200
rect 139900 23200 140000 23300
rect 139900 23300 140000 23400
rect 139900 23400 140000 23500
rect 139900 23500 140000 23600
rect 139900 23600 140000 23700
rect 139900 23700 140000 23800
rect 139900 36000 140000 36100
rect 139900 36100 140000 36200
rect 139900 36200 140000 36300
rect 139900 36300 140000 36400
rect 139900 36400 140000 36500
rect 139900 36500 140000 36600
rect 139900 36600 140000 36700
rect 139900 36700 140000 36800
rect 139900 36800 140000 36900
rect 139900 36900 140000 37000
rect 139900 37000 140000 37100
rect 139900 37100 140000 37200
rect 139900 37200 140000 37300
rect 139900 37300 140000 37400
rect 139900 37400 140000 37500
rect 139900 37500 140000 37600
rect 139900 37600 140000 37700
rect 139900 37700 140000 37800
rect 139900 37800 140000 37900
rect 139900 37900 140000 38000
rect 139900 38000 140000 38100
rect 139900 38100 140000 38200
rect 140000 21600 140100 21700
rect 140000 21700 140100 21800
rect 140000 21800 140100 21900
rect 140000 21900 140100 22000
rect 140000 22000 140100 22100
rect 140000 22100 140100 22200
rect 140000 22200 140100 22300
rect 140000 22300 140100 22400
rect 140000 22400 140100 22500
rect 140000 22500 140100 22600
rect 140000 22600 140100 22700
rect 140000 22700 140100 22800
rect 140000 22800 140100 22900
rect 140000 22900 140100 23000
rect 140000 23000 140100 23100
rect 140000 23100 140100 23200
rect 140000 23200 140100 23300
rect 140000 23300 140100 23400
rect 140000 23400 140100 23500
rect 140000 23500 140100 23600
rect 140000 23600 140100 23700
rect 140000 23700 140100 23800
rect 140000 36100 140100 36200
rect 140000 36200 140100 36300
rect 140000 36300 140100 36400
rect 140000 36400 140100 36500
rect 140000 36500 140100 36600
rect 140000 36600 140100 36700
rect 140000 36700 140100 36800
rect 140000 36800 140100 36900
rect 140000 36900 140100 37000
rect 140000 37000 140100 37100
rect 140000 37100 140100 37200
rect 140000 37200 140100 37300
rect 140000 37300 140100 37400
rect 140000 37400 140100 37500
rect 140000 37500 140100 37600
rect 140000 37600 140100 37700
rect 140000 37700 140100 37800
rect 140000 37800 140100 37900
rect 140000 37900 140100 38000
rect 140000 38000 140100 38100
rect 140000 38100 140100 38200
rect 140100 21600 140200 21700
rect 140100 21700 140200 21800
rect 140100 21800 140200 21900
rect 140100 21900 140200 22000
rect 140100 22000 140200 22100
rect 140100 22100 140200 22200
rect 140100 22200 140200 22300
rect 140100 22300 140200 22400
rect 140100 22400 140200 22500
rect 140100 22500 140200 22600
rect 140100 22600 140200 22700
rect 140100 22700 140200 22800
rect 140100 22800 140200 22900
rect 140100 22900 140200 23000
rect 140100 23000 140200 23100
rect 140100 23100 140200 23200
rect 140100 23200 140200 23300
rect 140100 23300 140200 23400
rect 140100 23400 140200 23500
rect 140100 23500 140200 23600
rect 140100 23600 140200 23700
rect 140100 23700 140200 23800
rect 140100 36100 140200 36200
rect 140100 36200 140200 36300
rect 140100 36300 140200 36400
rect 140100 36400 140200 36500
rect 140100 36500 140200 36600
rect 140100 36600 140200 36700
rect 140100 36700 140200 36800
rect 140100 36800 140200 36900
rect 140100 36900 140200 37000
rect 140100 37000 140200 37100
rect 140100 37100 140200 37200
rect 140100 37200 140200 37300
rect 140100 37300 140200 37400
rect 140100 37400 140200 37500
rect 140100 37500 140200 37600
rect 140100 37600 140200 37700
rect 140100 37700 140200 37800
rect 140100 37800 140200 37900
rect 140100 37900 140200 38000
rect 140100 38000 140200 38100
rect 140100 38100 140200 38200
rect 140100 38200 140200 38300
rect 140200 21600 140300 21700
rect 140200 21700 140300 21800
rect 140200 21800 140300 21900
rect 140200 21900 140300 22000
rect 140200 22000 140300 22100
rect 140200 22100 140300 22200
rect 140200 22200 140300 22300
rect 140200 22300 140300 22400
rect 140200 22400 140300 22500
rect 140200 22500 140300 22600
rect 140200 22600 140300 22700
rect 140200 22700 140300 22800
rect 140200 22800 140300 22900
rect 140200 22900 140300 23000
rect 140200 23000 140300 23100
rect 140200 23100 140300 23200
rect 140200 23200 140300 23300
rect 140200 23300 140300 23400
rect 140200 23400 140300 23500
rect 140200 23500 140300 23600
rect 140200 23600 140300 23700
rect 140200 23700 140300 23800
rect 140200 36100 140300 36200
rect 140200 36200 140300 36300
rect 140200 36300 140300 36400
rect 140200 36400 140300 36500
rect 140200 36500 140300 36600
rect 140200 36600 140300 36700
rect 140200 36700 140300 36800
rect 140200 36800 140300 36900
rect 140200 36900 140300 37000
rect 140200 37000 140300 37100
rect 140200 37100 140300 37200
rect 140200 37200 140300 37300
rect 140200 37300 140300 37400
rect 140200 37400 140300 37500
rect 140200 37500 140300 37600
rect 140200 37600 140300 37700
rect 140200 37700 140300 37800
rect 140200 37800 140300 37900
rect 140200 37900 140300 38000
rect 140200 38000 140300 38100
rect 140200 38100 140300 38200
rect 140200 38200 140300 38300
rect 140300 21600 140400 21700
rect 140300 21700 140400 21800
rect 140300 21800 140400 21900
rect 140300 21900 140400 22000
rect 140300 22000 140400 22100
rect 140300 22100 140400 22200
rect 140300 22200 140400 22300
rect 140300 22300 140400 22400
rect 140300 22400 140400 22500
rect 140300 22500 140400 22600
rect 140300 22600 140400 22700
rect 140300 22700 140400 22800
rect 140300 22800 140400 22900
rect 140300 22900 140400 23000
rect 140300 23000 140400 23100
rect 140300 23100 140400 23200
rect 140300 23200 140400 23300
rect 140300 23300 140400 23400
rect 140300 23400 140400 23500
rect 140300 23500 140400 23600
rect 140300 23600 140400 23700
rect 140300 23700 140400 23800
rect 140300 36100 140400 36200
rect 140300 36200 140400 36300
rect 140300 36300 140400 36400
rect 140300 36400 140400 36500
rect 140300 36500 140400 36600
rect 140300 36600 140400 36700
rect 140300 36700 140400 36800
rect 140300 36800 140400 36900
rect 140300 36900 140400 37000
rect 140300 37000 140400 37100
rect 140300 37100 140400 37200
rect 140300 37200 140400 37300
rect 140300 37300 140400 37400
rect 140300 37400 140400 37500
rect 140300 37500 140400 37600
rect 140300 37600 140400 37700
rect 140300 37700 140400 37800
rect 140300 37800 140400 37900
rect 140300 37900 140400 38000
rect 140300 38000 140400 38100
rect 140300 38100 140400 38200
rect 140300 38200 140400 38300
rect 140400 21600 140500 21700
rect 140400 21700 140500 21800
rect 140400 21800 140500 21900
rect 140400 21900 140500 22000
rect 140400 22000 140500 22100
rect 140400 22100 140500 22200
rect 140400 22200 140500 22300
rect 140400 22300 140500 22400
rect 140400 22400 140500 22500
rect 140400 22500 140500 22600
rect 140400 22600 140500 22700
rect 140400 22700 140500 22800
rect 140400 22800 140500 22900
rect 140400 22900 140500 23000
rect 140400 23000 140500 23100
rect 140400 23100 140500 23200
rect 140400 23200 140500 23300
rect 140400 23300 140500 23400
rect 140400 23400 140500 23500
rect 140400 23500 140500 23600
rect 140400 23600 140500 23700
rect 140400 23700 140500 23800
rect 140400 36100 140500 36200
rect 140400 36200 140500 36300
rect 140400 36300 140500 36400
rect 140400 36400 140500 36500
rect 140400 36500 140500 36600
rect 140400 36600 140500 36700
rect 140400 36700 140500 36800
rect 140400 36800 140500 36900
rect 140400 36900 140500 37000
rect 140400 37000 140500 37100
rect 140400 37100 140500 37200
rect 140400 37200 140500 37300
rect 140400 37300 140500 37400
rect 140400 37400 140500 37500
rect 140400 37500 140500 37600
rect 140400 37600 140500 37700
rect 140400 37700 140500 37800
rect 140400 37800 140500 37900
rect 140400 37900 140500 38000
rect 140400 38000 140500 38100
rect 140400 38100 140500 38200
rect 140400 38200 140500 38300
rect 140500 21600 140600 21700
rect 140500 21700 140600 21800
rect 140500 21800 140600 21900
rect 140500 21900 140600 22000
rect 140500 22000 140600 22100
rect 140500 22100 140600 22200
rect 140500 22200 140600 22300
rect 140500 22300 140600 22400
rect 140500 22400 140600 22500
rect 140500 22500 140600 22600
rect 140500 22600 140600 22700
rect 140500 22700 140600 22800
rect 140500 22800 140600 22900
rect 140500 22900 140600 23000
rect 140500 23000 140600 23100
rect 140500 23100 140600 23200
rect 140500 23200 140600 23300
rect 140500 23300 140600 23400
rect 140500 23400 140600 23500
rect 140500 23500 140600 23600
rect 140500 23600 140600 23700
rect 140500 23700 140600 23800
rect 140500 36100 140600 36200
rect 140500 36200 140600 36300
rect 140500 36300 140600 36400
rect 140500 36400 140600 36500
rect 140500 36500 140600 36600
rect 140500 36600 140600 36700
rect 140500 36700 140600 36800
rect 140500 36800 140600 36900
rect 140500 36900 140600 37000
rect 140500 37000 140600 37100
rect 140500 37100 140600 37200
rect 140500 37200 140600 37300
rect 140500 37300 140600 37400
rect 140500 37400 140600 37500
rect 140500 37500 140600 37600
rect 140500 37600 140600 37700
rect 140500 37700 140600 37800
rect 140500 37800 140600 37900
rect 140500 37900 140600 38000
rect 140500 38000 140600 38100
rect 140500 38100 140600 38200
rect 140500 38200 140600 38300
rect 140600 21600 140700 21700
rect 140600 21700 140700 21800
rect 140600 21800 140700 21900
rect 140600 21900 140700 22000
rect 140600 22000 140700 22100
rect 140600 22100 140700 22200
rect 140600 22200 140700 22300
rect 140600 22300 140700 22400
rect 140600 22400 140700 22500
rect 140600 22500 140700 22600
rect 140600 22600 140700 22700
rect 140600 22700 140700 22800
rect 140600 22800 140700 22900
rect 140600 22900 140700 23000
rect 140600 23000 140700 23100
rect 140600 23100 140700 23200
rect 140600 23200 140700 23300
rect 140600 23300 140700 23400
rect 140600 23400 140700 23500
rect 140600 23500 140700 23600
rect 140600 23600 140700 23700
rect 140600 23700 140700 23800
rect 140600 36100 140700 36200
rect 140600 36200 140700 36300
rect 140600 36300 140700 36400
rect 140600 36400 140700 36500
rect 140600 36500 140700 36600
rect 140600 36600 140700 36700
rect 140600 36700 140700 36800
rect 140600 36800 140700 36900
rect 140600 36900 140700 37000
rect 140600 37000 140700 37100
rect 140600 37100 140700 37200
rect 140600 37200 140700 37300
rect 140600 37300 140700 37400
rect 140600 37400 140700 37500
rect 140600 37500 140700 37600
rect 140600 37600 140700 37700
rect 140600 37700 140700 37800
rect 140600 37800 140700 37900
rect 140600 37900 140700 38000
rect 140600 38000 140700 38100
rect 140600 38100 140700 38200
rect 140600 38200 140700 38300
rect 140700 21700 140800 21800
rect 140700 21800 140800 21900
rect 140700 21900 140800 22000
rect 140700 22000 140800 22100
rect 140700 22100 140800 22200
rect 140700 22200 140800 22300
rect 140700 22300 140800 22400
rect 140700 22400 140800 22500
rect 140700 22500 140800 22600
rect 140700 22600 140800 22700
rect 140700 22700 140800 22800
rect 140700 22800 140800 22900
rect 140700 22900 140800 23000
rect 140700 23000 140800 23100
rect 140700 23100 140800 23200
rect 140700 23200 140800 23300
rect 140700 23300 140800 23400
rect 140700 23400 140800 23500
rect 140700 23500 140800 23600
rect 140700 23600 140800 23700
rect 140700 23700 140800 23800
rect 140700 36100 140800 36200
rect 140700 36200 140800 36300
rect 140700 36300 140800 36400
rect 140700 36400 140800 36500
rect 140700 36500 140800 36600
rect 140700 36600 140800 36700
rect 140700 36700 140800 36800
rect 140700 36800 140800 36900
rect 140700 36900 140800 37000
rect 140700 37000 140800 37100
rect 140700 37100 140800 37200
rect 140700 37200 140800 37300
rect 140700 37300 140800 37400
rect 140700 37400 140800 37500
rect 140700 37500 140800 37600
rect 140700 37600 140800 37700
rect 140700 37700 140800 37800
rect 140700 37800 140800 37900
rect 140700 37900 140800 38000
rect 140700 38000 140800 38100
rect 140700 38100 140800 38200
rect 140700 38200 140800 38300
rect 140800 21700 140900 21800
rect 140800 21800 140900 21900
rect 140800 21900 140900 22000
rect 140800 22000 140900 22100
rect 140800 22100 140900 22200
rect 140800 22200 140900 22300
rect 140800 22300 140900 22400
rect 140800 22400 140900 22500
rect 140800 22500 140900 22600
rect 140800 22600 140900 22700
rect 140800 22700 140900 22800
rect 140800 22800 140900 22900
rect 140800 22900 140900 23000
rect 140800 23000 140900 23100
rect 140800 23100 140900 23200
rect 140800 23200 140900 23300
rect 140800 23300 140900 23400
rect 140800 23400 140900 23500
rect 140800 23500 140900 23600
rect 140800 23600 140900 23700
rect 140800 23700 140900 23800
rect 140800 23800 140900 23900
rect 140800 36100 140900 36200
rect 140800 36200 140900 36300
rect 140800 36300 140900 36400
rect 140800 36400 140900 36500
rect 140800 36500 140900 36600
rect 140800 36600 140900 36700
rect 140800 36700 140900 36800
rect 140800 36800 140900 36900
rect 140800 36900 140900 37000
rect 140800 37000 140900 37100
rect 140800 37100 140900 37200
rect 140800 37200 140900 37300
rect 140800 37300 140900 37400
rect 140800 37400 140900 37500
rect 140800 37500 140900 37600
rect 140800 37600 140900 37700
rect 140800 37700 140900 37800
rect 140800 37800 140900 37900
rect 140800 37900 140900 38000
rect 140800 38000 140900 38100
rect 140800 38100 140900 38200
rect 140800 38200 140900 38300
rect 140900 21700 141000 21800
rect 140900 21800 141000 21900
rect 140900 21900 141000 22000
rect 140900 22000 141000 22100
rect 140900 22100 141000 22200
rect 140900 22200 141000 22300
rect 140900 22300 141000 22400
rect 140900 22400 141000 22500
rect 140900 22500 141000 22600
rect 140900 22600 141000 22700
rect 140900 22700 141000 22800
rect 140900 22800 141000 22900
rect 140900 22900 141000 23000
rect 140900 23000 141000 23100
rect 140900 23100 141000 23200
rect 140900 23200 141000 23300
rect 140900 23300 141000 23400
rect 140900 23400 141000 23500
rect 140900 23500 141000 23600
rect 140900 23600 141000 23700
rect 140900 23700 141000 23800
rect 140900 23800 141000 23900
rect 140900 36100 141000 36200
rect 140900 36200 141000 36300
rect 140900 36300 141000 36400
rect 140900 36400 141000 36500
rect 140900 36500 141000 36600
rect 140900 36600 141000 36700
rect 140900 36700 141000 36800
rect 140900 36800 141000 36900
rect 140900 36900 141000 37000
rect 140900 37000 141000 37100
rect 140900 37100 141000 37200
rect 140900 37200 141000 37300
rect 140900 37300 141000 37400
rect 140900 37400 141000 37500
rect 140900 37500 141000 37600
rect 140900 37600 141000 37700
rect 140900 37700 141000 37800
rect 140900 37800 141000 37900
rect 140900 37900 141000 38000
rect 140900 38000 141000 38100
rect 140900 38100 141000 38200
rect 140900 38200 141000 38300
rect 141000 21700 141100 21800
rect 141000 21800 141100 21900
rect 141000 21900 141100 22000
rect 141000 22000 141100 22100
rect 141000 22100 141100 22200
rect 141000 22200 141100 22300
rect 141000 22300 141100 22400
rect 141000 22400 141100 22500
rect 141000 22500 141100 22600
rect 141000 22600 141100 22700
rect 141000 22700 141100 22800
rect 141000 22800 141100 22900
rect 141000 22900 141100 23000
rect 141000 23000 141100 23100
rect 141000 23100 141100 23200
rect 141000 23200 141100 23300
rect 141000 23300 141100 23400
rect 141000 23400 141100 23500
rect 141000 23500 141100 23600
rect 141000 23600 141100 23700
rect 141000 23700 141100 23800
rect 141000 23800 141100 23900
rect 141000 36200 141100 36300
rect 141000 36300 141100 36400
rect 141000 36400 141100 36500
rect 141000 36500 141100 36600
rect 141000 36600 141100 36700
rect 141000 36700 141100 36800
rect 141000 36800 141100 36900
rect 141000 36900 141100 37000
rect 141000 37000 141100 37100
rect 141000 37100 141100 37200
rect 141000 37200 141100 37300
rect 141000 37300 141100 37400
rect 141000 37400 141100 37500
rect 141000 37500 141100 37600
rect 141000 37600 141100 37700
rect 141000 37700 141100 37800
rect 141000 37800 141100 37900
rect 141000 37900 141100 38000
rect 141000 38000 141100 38100
rect 141000 38100 141100 38200
rect 141000 38200 141100 38300
rect 141100 21700 141200 21800
rect 141100 21800 141200 21900
rect 141100 21900 141200 22000
rect 141100 22000 141200 22100
rect 141100 22100 141200 22200
rect 141100 22200 141200 22300
rect 141100 22300 141200 22400
rect 141100 22400 141200 22500
rect 141100 22500 141200 22600
rect 141100 22600 141200 22700
rect 141100 22700 141200 22800
rect 141100 22800 141200 22900
rect 141100 22900 141200 23000
rect 141100 23000 141200 23100
rect 141100 23100 141200 23200
rect 141100 23200 141200 23300
rect 141100 23300 141200 23400
rect 141100 23400 141200 23500
rect 141100 23500 141200 23600
rect 141100 23600 141200 23700
rect 141100 23700 141200 23800
rect 141100 23800 141200 23900
rect 141100 36100 141200 36200
rect 141100 36200 141200 36300
rect 141100 36300 141200 36400
rect 141100 36400 141200 36500
rect 141100 36500 141200 36600
rect 141100 36600 141200 36700
rect 141100 36700 141200 36800
rect 141100 36800 141200 36900
rect 141100 36900 141200 37000
rect 141100 37000 141200 37100
rect 141100 37100 141200 37200
rect 141100 37200 141200 37300
rect 141100 37300 141200 37400
rect 141100 37400 141200 37500
rect 141100 37500 141200 37600
rect 141100 37600 141200 37700
rect 141100 37700 141200 37800
rect 141100 37800 141200 37900
rect 141100 37900 141200 38000
rect 141100 38000 141200 38100
rect 141100 38100 141200 38200
rect 141100 38200 141200 38300
rect 141200 21700 141300 21800
rect 141200 21800 141300 21900
rect 141200 21900 141300 22000
rect 141200 22000 141300 22100
rect 141200 22100 141300 22200
rect 141200 22200 141300 22300
rect 141200 22300 141300 22400
rect 141200 22400 141300 22500
rect 141200 22500 141300 22600
rect 141200 22600 141300 22700
rect 141200 22700 141300 22800
rect 141200 22800 141300 22900
rect 141200 22900 141300 23000
rect 141200 23000 141300 23100
rect 141200 23100 141300 23200
rect 141200 23200 141300 23300
rect 141200 23300 141300 23400
rect 141200 23400 141300 23500
rect 141200 23500 141300 23600
rect 141200 23600 141300 23700
rect 141200 23700 141300 23800
rect 141200 23800 141300 23900
rect 141200 23900 141300 24000
rect 141200 36200 141300 36300
rect 141200 36300 141300 36400
rect 141200 36400 141300 36500
rect 141200 36500 141300 36600
rect 141200 36600 141300 36700
rect 141200 36700 141300 36800
rect 141200 36800 141300 36900
rect 141200 36900 141300 37000
rect 141200 37000 141300 37100
rect 141200 37100 141300 37200
rect 141200 37200 141300 37300
rect 141200 37300 141300 37400
rect 141200 37400 141300 37500
rect 141200 37500 141300 37600
rect 141200 37600 141300 37700
rect 141200 37700 141300 37800
rect 141200 37800 141300 37900
rect 141200 37900 141300 38000
rect 141200 38000 141300 38100
rect 141200 38100 141300 38200
rect 141200 38200 141300 38300
rect 141300 21700 141400 21800
rect 141300 21800 141400 21900
rect 141300 21900 141400 22000
rect 141300 22000 141400 22100
rect 141300 22100 141400 22200
rect 141300 22200 141400 22300
rect 141300 22300 141400 22400
rect 141300 22400 141400 22500
rect 141300 22500 141400 22600
rect 141300 22600 141400 22700
rect 141300 22700 141400 22800
rect 141300 22800 141400 22900
rect 141300 22900 141400 23000
rect 141300 23000 141400 23100
rect 141300 23100 141400 23200
rect 141300 23200 141400 23300
rect 141300 23300 141400 23400
rect 141300 23400 141400 23500
rect 141300 23500 141400 23600
rect 141300 23600 141400 23700
rect 141300 23700 141400 23800
rect 141300 23800 141400 23900
rect 141300 23900 141400 24000
rect 141300 36100 141400 36200
rect 141300 36200 141400 36300
rect 141300 36300 141400 36400
rect 141300 36400 141400 36500
rect 141300 36500 141400 36600
rect 141300 36600 141400 36700
rect 141300 36700 141400 36800
rect 141300 36800 141400 36900
rect 141300 36900 141400 37000
rect 141300 37000 141400 37100
rect 141300 37100 141400 37200
rect 141300 37200 141400 37300
rect 141300 37300 141400 37400
rect 141300 37400 141400 37500
rect 141300 37500 141400 37600
rect 141300 37600 141400 37700
rect 141300 37700 141400 37800
rect 141300 37800 141400 37900
rect 141300 37900 141400 38000
rect 141300 38000 141400 38100
rect 141300 38100 141400 38200
rect 141300 38200 141400 38300
rect 141400 21800 141500 21900
rect 141400 21900 141500 22000
rect 141400 22000 141500 22100
rect 141400 22100 141500 22200
rect 141400 22200 141500 22300
rect 141400 22300 141500 22400
rect 141400 22400 141500 22500
rect 141400 22500 141500 22600
rect 141400 22600 141500 22700
rect 141400 22700 141500 22800
rect 141400 22800 141500 22900
rect 141400 22900 141500 23000
rect 141400 23000 141500 23100
rect 141400 23100 141500 23200
rect 141400 23200 141500 23300
rect 141400 23300 141500 23400
rect 141400 23400 141500 23500
rect 141400 23500 141500 23600
rect 141400 23600 141500 23700
rect 141400 23700 141500 23800
rect 141400 23800 141500 23900
rect 141400 23900 141500 24000
rect 141400 36100 141500 36200
rect 141400 36200 141500 36300
rect 141400 36300 141500 36400
rect 141400 36400 141500 36500
rect 141400 36500 141500 36600
rect 141400 36600 141500 36700
rect 141400 36700 141500 36800
rect 141400 36800 141500 36900
rect 141400 36900 141500 37000
rect 141400 37000 141500 37100
rect 141400 37100 141500 37200
rect 141400 37200 141500 37300
rect 141400 37300 141500 37400
rect 141400 37400 141500 37500
rect 141400 37500 141500 37600
rect 141400 37600 141500 37700
rect 141400 37700 141500 37800
rect 141400 37800 141500 37900
rect 141400 37900 141500 38000
rect 141400 38000 141500 38100
rect 141400 38100 141500 38200
rect 141400 38200 141500 38300
rect 141500 21800 141600 21900
rect 141500 21900 141600 22000
rect 141500 22000 141600 22100
rect 141500 22100 141600 22200
rect 141500 22200 141600 22300
rect 141500 22300 141600 22400
rect 141500 22400 141600 22500
rect 141500 22500 141600 22600
rect 141500 22600 141600 22700
rect 141500 22700 141600 22800
rect 141500 22800 141600 22900
rect 141500 22900 141600 23000
rect 141500 23000 141600 23100
rect 141500 23100 141600 23200
rect 141500 23200 141600 23300
rect 141500 23300 141600 23400
rect 141500 23400 141600 23500
rect 141500 23500 141600 23600
rect 141500 23600 141600 23700
rect 141500 23700 141600 23800
rect 141500 23800 141600 23900
rect 141500 23900 141600 24000
rect 141500 24000 141600 24100
rect 141500 36200 141600 36300
rect 141500 36300 141600 36400
rect 141500 36400 141600 36500
rect 141500 36500 141600 36600
rect 141500 36600 141600 36700
rect 141500 36700 141600 36800
rect 141500 36800 141600 36900
rect 141500 36900 141600 37000
rect 141500 37000 141600 37100
rect 141500 37100 141600 37200
rect 141500 37200 141600 37300
rect 141500 37300 141600 37400
rect 141500 37400 141600 37500
rect 141500 37500 141600 37600
rect 141500 37600 141600 37700
rect 141500 37700 141600 37800
rect 141500 37800 141600 37900
rect 141500 37900 141600 38000
rect 141500 38000 141600 38100
rect 141500 38100 141600 38200
rect 141500 38200 141600 38300
rect 141600 21800 141700 21900
rect 141600 21900 141700 22000
rect 141600 22000 141700 22100
rect 141600 22100 141700 22200
rect 141600 22200 141700 22300
rect 141600 22300 141700 22400
rect 141600 22400 141700 22500
rect 141600 22500 141700 22600
rect 141600 22600 141700 22700
rect 141600 22700 141700 22800
rect 141600 22800 141700 22900
rect 141600 22900 141700 23000
rect 141600 23000 141700 23100
rect 141600 23100 141700 23200
rect 141600 23200 141700 23300
rect 141600 23300 141700 23400
rect 141600 23400 141700 23500
rect 141600 23500 141700 23600
rect 141600 23600 141700 23700
rect 141600 23700 141700 23800
rect 141600 23800 141700 23900
rect 141600 23900 141700 24000
rect 141600 24000 141700 24100
rect 141600 36100 141700 36200
rect 141600 36200 141700 36300
rect 141600 36300 141700 36400
rect 141600 36400 141700 36500
rect 141600 36500 141700 36600
rect 141600 36600 141700 36700
rect 141600 36700 141700 36800
rect 141600 36800 141700 36900
rect 141600 36900 141700 37000
rect 141600 37000 141700 37100
rect 141600 37100 141700 37200
rect 141600 37200 141700 37300
rect 141600 37300 141700 37400
rect 141600 37400 141700 37500
rect 141600 37500 141700 37600
rect 141600 37600 141700 37700
rect 141600 37700 141700 37800
rect 141600 37800 141700 37900
rect 141600 37900 141700 38000
rect 141600 38000 141700 38100
rect 141600 38100 141700 38200
rect 141600 38200 141700 38300
rect 141700 21800 141800 21900
rect 141700 21900 141800 22000
rect 141700 22000 141800 22100
rect 141700 22100 141800 22200
rect 141700 22200 141800 22300
rect 141700 22300 141800 22400
rect 141700 22400 141800 22500
rect 141700 22500 141800 22600
rect 141700 22600 141800 22700
rect 141700 22700 141800 22800
rect 141700 22800 141800 22900
rect 141700 22900 141800 23000
rect 141700 23000 141800 23100
rect 141700 23100 141800 23200
rect 141700 23200 141800 23300
rect 141700 23300 141800 23400
rect 141700 23400 141800 23500
rect 141700 23500 141800 23600
rect 141700 23600 141800 23700
rect 141700 23700 141800 23800
rect 141700 23800 141800 23900
rect 141700 23900 141800 24000
rect 141700 24000 141800 24100
rect 141700 36100 141800 36200
rect 141700 36200 141800 36300
rect 141700 36300 141800 36400
rect 141700 36400 141800 36500
rect 141700 36500 141800 36600
rect 141700 36600 141800 36700
rect 141700 36700 141800 36800
rect 141700 36800 141800 36900
rect 141700 36900 141800 37000
rect 141700 37000 141800 37100
rect 141700 37100 141800 37200
rect 141700 37200 141800 37300
rect 141700 37300 141800 37400
rect 141700 37400 141800 37500
rect 141700 37500 141800 37600
rect 141700 37600 141800 37700
rect 141700 37700 141800 37800
rect 141700 37800 141800 37900
rect 141700 37900 141800 38000
rect 141700 38000 141800 38100
rect 141700 38100 141800 38200
rect 141700 38200 141800 38300
rect 141800 21900 141900 22000
rect 141800 22000 141900 22100
rect 141800 22100 141900 22200
rect 141800 22200 141900 22300
rect 141800 22300 141900 22400
rect 141800 22400 141900 22500
rect 141800 22500 141900 22600
rect 141800 22600 141900 22700
rect 141800 22700 141900 22800
rect 141800 22800 141900 22900
rect 141800 22900 141900 23000
rect 141800 23000 141900 23100
rect 141800 23100 141900 23200
rect 141800 23200 141900 23300
rect 141800 23300 141900 23400
rect 141800 23400 141900 23500
rect 141800 23500 141900 23600
rect 141800 23600 141900 23700
rect 141800 23700 141900 23800
rect 141800 23800 141900 23900
rect 141800 23900 141900 24000
rect 141800 24000 141900 24100
rect 141800 24100 141900 24200
rect 141800 36100 141900 36200
rect 141800 36200 141900 36300
rect 141800 36300 141900 36400
rect 141800 36400 141900 36500
rect 141800 36500 141900 36600
rect 141800 36600 141900 36700
rect 141800 36700 141900 36800
rect 141800 36800 141900 36900
rect 141800 36900 141900 37000
rect 141800 37000 141900 37100
rect 141800 37100 141900 37200
rect 141800 37200 141900 37300
rect 141800 37300 141900 37400
rect 141800 37400 141900 37500
rect 141800 37500 141900 37600
rect 141800 37600 141900 37700
rect 141800 37700 141900 37800
rect 141800 37800 141900 37900
rect 141800 37900 141900 38000
rect 141800 38000 141900 38100
rect 141800 38100 141900 38200
rect 141800 38200 141900 38300
rect 141900 21900 142000 22000
rect 141900 22000 142000 22100
rect 141900 22100 142000 22200
rect 141900 22200 142000 22300
rect 141900 22300 142000 22400
rect 141900 22400 142000 22500
rect 141900 22500 142000 22600
rect 141900 22600 142000 22700
rect 141900 22700 142000 22800
rect 141900 22800 142000 22900
rect 141900 22900 142000 23000
rect 141900 23000 142000 23100
rect 141900 23100 142000 23200
rect 141900 23200 142000 23300
rect 141900 23300 142000 23400
rect 141900 23400 142000 23500
rect 141900 23500 142000 23600
rect 141900 23600 142000 23700
rect 141900 23700 142000 23800
rect 141900 23800 142000 23900
rect 141900 23900 142000 24000
rect 141900 24000 142000 24100
rect 141900 24100 142000 24200
rect 141900 36100 142000 36200
rect 141900 36200 142000 36300
rect 141900 36300 142000 36400
rect 141900 36400 142000 36500
rect 141900 36500 142000 36600
rect 141900 36600 142000 36700
rect 141900 36700 142000 36800
rect 141900 36800 142000 36900
rect 141900 36900 142000 37000
rect 141900 37000 142000 37100
rect 141900 37100 142000 37200
rect 141900 37200 142000 37300
rect 141900 37300 142000 37400
rect 141900 37400 142000 37500
rect 141900 37500 142000 37600
rect 141900 37600 142000 37700
rect 141900 37700 142000 37800
rect 141900 37800 142000 37900
rect 141900 37900 142000 38000
rect 141900 38000 142000 38100
rect 141900 38100 142000 38200
rect 141900 38200 142000 38300
rect 142000 21900 142100 22000
rect 142000 22000 142100 22100
rect 142000 22100 142100 22200
rect 142000 22200 142100 22300
rect 142000 22300 142100 22400
rect 142000 22400 142100 22500
rect 142000 22500 142100 22600
rect 142000 22600 142100 22700
rect 142000 22700 142100 22800
rect 142000 22800 142100 22900
rect 142000 22900 142100 23000
rect 142000 23000 142100 23100
rect 142000 23100 142100 23200
rect 142000 23200 142100 23300
rect 142000 23300 142100 23400
rect 142000 23400 142100 23500
rect 142000 23500 142100 23600
rect 142000 23600 142100 23700
rect 142000 23700 142100 23800
rect 142000 23800 142100 23900
rect 142000 23900 142100 24000
rect 142000 24000 142100 24100
rect 142000 24100 142100 24200
rect 142000 24200 142100 24300
rect 142000 36100 142100 36200
rect 142000 36200 142100 36300
rect 142000 36300 142100 36400
rect 142000 36400 142100 36500
rect 142000 36500 142100 36600
rect 142000 36600 142100 36700
rect 142000 36700 142100 36800
rect 142000 36800 142100 36900
rect 142000 36900 142100 37000
rect 142000 37000 142100 37100
rect 142000 37100 142100 37200
rect 142000 37200 142100 37300
rect 142000 37300 142100 37400
rect 142000 37400 142100 37500
rect 142000 37500 142100 37600
rect 142000 37600 142100 37700
rect 142000 37700 142100 37800
rect 142000 37800 142100 37900
rect 142000 37900 142100 38000
rect 142000 38000 142100 38100
rect 142000 38100 142100 38200
rect 142000 38200 142100 38300
rect 142100 22000 142200 22100
rect 142100 22100 142200 22200
rect 142100 22200 142200 22300
rect 142100 22300 142200 22400
rect 142100 22400 142200 22500
rect 142100 22500 142200 22600
rect 142100 22600 142200 22700
rect 142100 22700 142200 22800
rect 142100 22800 142200 22900
rect 142100 22900 142200 23000
rect 142100 23000 142200 23100
rect 142100 23100 142200 23200
rect 142100 23200 142200 23300
rect 142100 23300 142200 23400
rect 142100 23400 142200 23500
rect 142100 23500 142200 23600
rect 142100 23600 142200 23700
rect 142100 23700 142200 23800
rect 142100 23800 142200 23900
rect 142100 23900 142200 24000
rect 142100 24000 142200 24100
rect 142100 24100 142200 24200
rect 142100 24200 142200 24300
rect 142100 24300 142200 24400
rect 142100 36100 142200 36200
rect 142100 36200 142200 36300
rect 142100 36300 142200 36400
rect 142100 36400 142200 36500
rect 142100 36500 142200 36600
rect 142100 36600 142200 36700
rect 142100 36700 142200 36800
rect 142100 36800 142200 36900
rect 142100 36900 142200 37000
rect 142100 37000 142200 37100
rect 142100 37100 142200 37200
rect 142100 37200 142200 37300
rect 142100 37300 142200 37400
rect 142100 37400 142200 37500
rect 142100 37500 142200 37600
rect 142100 37600 142200 37700
rect 142100 37700 142200 37800
rect 142100 37800 142200 37900
rect 142100 37900 142200 38000
rect 142100 38000 142200 38100
rect 142100 38100 142200 38200
rect 142100 38200 142200 38300
rect 142200 22000 142300 22100
rect 142200 22100 142300 22200
rect 142200 22200 142300 22300
rect 142200 22300 142300 22400
rect 142200 22400 142300 22500
rect 142200 22500 142300 22600
rect 142200 22600 142300 22700
rect 142200 22700 142300 22800
rect 142200 22800 142300 22900
rect 142200 22900 142300 23000
rect 142200 23000 142300 23100
rect 142200 23100 142300 23200
rect 142200 23200 142300 23300
rect 142200 23300 142300 23400
rect 142200 23400 142300 23500
rect 142200 23500 142300 23600
rect 142200 23600 142300 23700
rect 142200 23700 142300 23800
rect 142200 23800 142300 23900
rect 142200 23900 142300 24000
rect 142200 24000 142300 24100
rect 142200 24100 142300 24200
rect 142200 24200 142300 24300
rect 142200 24300 142300 24400
rect 142200 36100 142300 36200
rect 142200 36200 142300 36300
rect 142200 36300 142300 36400
rect 142200 36400 142300 36500
rect 142200 36500 142300 36600
rect 142200 36600 142300 36700
rect 142200 36700 142300 36800
rect 142200 36800 142300 36900
rect 142200 36900 142300 37000
rect 142200 37000 142300 37100
rect 142200 37100 142300 37200
rect 142200 37200 142300 37300
rect 142200 37300 142300 37400
rect 142200 37400 142300 37500
rect 142200 37500 142300 37600
rect 142200 37600 142300 37700
rect 142200 37700 142300 37800
rect 142200 37800 142300 37900
rect 142200 37900 142300 38000
rect 142200 38000 142300 38100
rect 142200 38100 142300 38200
rect 142200 38200 142300 38300
rect 142300 22000 142400 22100
rect 142300 22100 142400 22200
rect 142300 22200 142400 22300
rect 142300 22300 142400 22400
rect 142300 22400 142400 22500
rect 142300 22500 142400 22600
rect 142300 22600 142400 22700
rect 142300 22700 142400 22800
rect 142300 22800 142400 22900
rect 142300 22900 142400 23000
rect 142300 23000 142400 23100
rect 142300 23100 142400 23200
rect 142300 23200 142400 23300
rect 142300 23300 142400 23400
rect 142300 23400 142400 23500
rect 142300 23500 142400 23600
rect 142300 23600 142400 23700
rect 142300 23700 142400 23800
rect 142300 23800 142400 23900
rect 142300 23900 142400 24000
rect 142300 24000 142400 24100
rect 142300 24100 142400 24200
rect 142300 24200 142400 24300
rect 142300 24300 142400 24400
rect 142300 24400 142400 24500
rect 142300 36000 142400 36100
rect 142300 36100 142400 36200
rect 142300 36200 142400 36300
rect 142300 36300 142400 36400
rect 142300 36400 142400 36500
rect 142300 36500 142400 36600
rect 142300 36600 142400 36700
rect 142300 36700 142400 36800
rect 142300 36800 142400 36900
rect 142300 36900 142400 37000
rect 142300 37000 142400 37100
rect 142300 37100 142400 37200
rect 142300 37200 142400 37300
rect 142300 37300 142400 37400
rect 142300 37400 142400 37500
rect 142300 37500 142400 37600
rect 142300 37600 142400 37700
rect 142300 37700 142400 37800
rect 142300 37800 142400 37900
rect 142300 37900 142400 38000
rect 142300 38000 142400 38100
rect 142300 38100 142400 38200
rect 142300 38200 142400 38300
rect 142400 22100 142500 22200
rect 142400 22200 142500 22300
rect 142400 22300 142500 22400
rect 142400 22400 142500 22500
rect 142400 22500 142500 22600
rect 142400 22600 142500 22700
rect 142400 22700 142500 22800
rect 142400 22800 142500 22900
rect 142400 22900 142500 23000
rect 142400 23000 142500 23100
rect 142400 23100 142500 23200
rect 142400 23200 142500 23300
rect 142400 23300 142500 23400
rect 142400 23400 142500 23500
rect 142400 23500 142500 23600
rect 142400 23600 142500 23700
rect 142400 23700 142500 23800
rect 142400 23800 142500 23900
rect 142400 23900 142500 24000
rect 142400 24000 142500 24100
rect 142400 24100 142500 24200
rect 142400 24200 142500 24300
rect 142400 24300 142500 24400
rect 142400 24400 142500 24500
rect 142400 24500 142500 24600
rect 142400 36000 142500 36100
rect 142400 36100 142500 36200
rect 142400 36200 142500 36300
rect 142400 36300 142500 36400
rect 142400 36400 142500 36500
rect 142400 36500 142500 36600
rect 142400 36600 142500 36700
rect 142400 36700 142500 36800
rect 142400 36800 142500 36900
rect 142400 36900 142500 37000
rect 142400 37000 142500 37100
rect 142400 37100 142500 37200
rect 142400 37200 142500 37300
rect 142400 37300 142500 37400
rect 142400 37400 142500 37500
rect 142400 37500 142500 37600
rect 142400 37600 142500 37700
rect 142400 37700 142500 37800
rect 142400 37800 142500 37900
rect 142400 37900 142500 38000
rect 142400 38000 142500 38100
rect 142400 38100 142500 38200
rect 142500 22100 142600 22200
rect 142500 22200 142600 22300
rect 142500 22300 142600 22400
rect 142500 22400 142600 22500
rect 142500 22500 142600 22600
rect 142500 22600 142600 22700
rect 142500 22700 142600 22800
rect 142500 22800 142600 22900
rect 142500 22900 142600 23000
rect 142500 23000 142600 23100
rect 142500 23100 142600 23200
rect 142500 23200 142600 23300
rect 142500 23300 142600 23400
rect 142500 23400 142600 23500
rect 142500 23500 142600 23600
rect 142500 23600 142600 23700
rect 142500 23700 142600 23800
rect 142500 23800 142600 23900
rect 142500 23900 142600 24000
rect 142500 24000 142600 24100
rect 142500 24100 142600 24200
rect 142500 24200 142600 24300
rect 142500 24300 142600 24400
rect 142500 24400 142600 24500
rect 142500 24500 142600 24600
rect 142500 36000 142600 36100
rect 142500 36100 142600 36200
rect 142500 36200 142600 36300
rect 142500 36300 142600 36400
rect 142500 36400 142600 36500
rect 142500 36500 142600 36600
rect 142500 36600 142600 36700
rect 142500 36700 142600 36800
rect 142500 36800 142600 36900
rect 142500 36900 142600 37000
rect 142500 37000 142600 37100
rect 142500 37100 142600 37200
rect 142500 37200 142600 37300
rect 142500 37300 142600 37400
rect 142500 37400 142600 37500
rect 142500 37500 142600 37600
rect 142500 37600 142600 37700
rect 142500 37700 142600 37800
rect 142500 37800 142600 37900
rect 142500 37900 142600 38000
rect 142500 38000 142600 38100
rect 142500 38100 142600 38200
rect 142600 22200 142700 22300
rect 142600 22300 142700 22400
rect 142600 22400 142700 22500
rect 142600 22500 142700 22600
rect 142600 22600 142700 22700
rect 142600 22700 142700 22800
rect 142600 22800 142700 22900
rect 142600 22900 142700 23000
rect 142600 23000 142700 23100
rect 142600 23100 142700 23200
rect 142600 23200 142700 23300
rect 142600 23300 142700 23400
rect 142600 23400 142700 23500
rect 142600 23500 142700 23600
rect 142600 23600 142700 23700
rect 142600 23700 142700 23800
rect 142600 23800 142700 23900
rect 142600 23900 142700 24000
rect 142600 24000 142700 24100
rect 142600 24100 142700 24200
rect 142600 24200 142700 24300
rect 142600 24300 142700 24400
rect 142600 24400 142700 24500
rect 142600 24500 142700 24600
rect 142600 24600 142700 24700
rect 142600 36000 142700 36100
rect 142600 36100 142700 36200
rect 142600 36200 142700 36300
rect 142600 36300 142700 36400
rect 142600 36400 142700 36500
rect 142600 36500 142700 36600
rect 142600 36600 142700 36700
rect 142600 36700 142700 36800
rect 142600 36800 142700 36900
rect 142600 36900 142700 37000
rect 142600 37000 142700 37100
rect 142600 37100 142700 37200
rect 142600 37200 142700 37300
rect 142600 37300 142700 37400
rect 142600 37400 142700 37500
rect 142600 37500 142700 37600
rect 142600 37600 142700 37700
rect 142600 37700 142700 37800
rect 142600 37800 142700 37900
rect 142600 37900 142700 38000
rect 142600 38000 142700 38100
rect 142600 38100 142700 38200
rect 142700 22200 142800 22300
rect 142700 22300 142800 22400
rect 142700 22400 142800 22500
rect 142700 22500 142800 22600
rect 142700 22600 142800 22700
rect 142700 22700 142800 22800
rect 142700 22800 142800 22900
rect 142700 22900 142800 23000
rect 142700 23000 142800 23100
rect 142700 23100 142800 23200
rect 142700 23200 142800 23300
rect 142700 23300 142800 23400
rect 142700 23400 142800 23500
rect 142700 23500 142800 23600
rect 142700 23600 142800 23700
rect 142700 23700 142800 23800
rect 142700 23800 142800 23900
rect 142700 23900 142800 24000
rect 142700 24000 142800 24100
rect 142700 24100 142800 24200
rect 142700 24200 142800 24300
rect 142700 24300 142800 24400
rect 142700 24400 142800 24500
rect 142700 24500 142800 24600
rect 142700 24600 142800 24700
rect 142700 24700 142800 24800
rect 142700 35900 142800 36000
rect 142700 36000 142800 36100
rect 142700 36100 142800 36200
rect 142700 36200 142800 36300
rect 142700 36300 142800 36400
rect 142700 36400 142800 36500
rect 142700 36500 142800 36600
rect 142700 36600 142800 36700
rect 142700 36700 142800 36800
rect 142700 36800 142800 36900
rect 142700 36900 142800 37000
rect 142700 37000 142800 37100
rect 142700 37100 142800 37200
rect 142700 37200 142800 37300
rect 142700 37300 142800 37400
rect 142700 37400 142800 37500
rect 142700 37500 142800 37600
rect 142700 37600 142800 37700
rect 142700 37700 142800 37800
rect 142700 37800 142800 37900
rect 142700 37900 142800 38000
rect 142700 38000 142800 38100
rect 142700 38100 142800 38200
rect 142800 22300 142900 22400
rect 142800 22400 142900 22500
rect 142800 22500 142900 22600
rect 142800 22600 142900 22700
rect 142800 22700 142900 22800
rect 142800 22800 142900 22900
rect 142800 22900 142900 23000
rect 142800 23000 142900 23100
rect 142800 23100 142900 23200
rect 142800 23200 142900 23300
rect 142800 23300 142900 23400
rect 142800 23400 142900 23500
rect 142800 23500 142900 23600
rect 142800 23600 142900 23700
rect 142800 23700 142900 23800
rect 142800 23800 142900 23900
rect 142800 23900 142900 24000
rect 142800 24000 142900 24100
rect 142800 24100 142900 24200
rect 142800 24200 142900 24300
rect 142800 24300 142900 24400
rect 142800 24400 142900 24500
rect 142800 24500 142900 24600
rect 142800 24600 142900 24700
rect 142800 24700 142900 24800
rect 142800 24800 142900 24900
rect 142800 35900 142900 36000
rect 142800 36000 142900 36100
rect 142800 36100 142900 36200
rect 142800 36200 142900 36300
rect 142800 36300 142900 36400
rect 142800 36400 142900 36500
rect 142800 36500 142900 36600
rect 142800 36600 142900 36700
rect 142800 36700 142900 36800
rect 142800 36800 142900 36900
rect 142800 36900 142900 37000
rect 142800 37000 142900 37100
rect 142800 37100 142900 37200
rect 142800 37200 142900 37300
rect 142800 37300 142900 37400
rect 142800 37400 142900 37500
rect 142800 37500 142900 37600
rect 142800 37600 142900 37700
rect 142800 37700 142900 37800
rect 142800 37800 142900 37900
rect 142800 37900 142900 38000
rect 142800 38000 142900 38100
rect 142800 38100 142900 38200
rect 142900 22300 143000 22400
rect 142900 22400 143000 22500
rect 142900 22500 143000 22600
rect 142900 22600 143000 22700
rect 142900 22700 143000 22800
rect 142900 22800 143000 22900
rect 142900 22900 143000 23000
rect 142900 23000 143000 23100
rect 142900 23100 143000 23200
rect 142900 23200 143000 23300
rect 142900 23300 143000 23400
rect 142900 23400 143000 23500
rect 142900 23500 143000 23600
rect 142900 23600 143000 23700
rect 142900 23700 143000 23800
rect 142900 23800 143000 23900
rect 142900 23900 143000 24000
rect 142900 24000 143000 24100
rect 142900 24100 143000 24200
rect 142900 24200 143000 24300
rect 142900 24300 143000 24400
rect 142900 24400 143000 24500
rect 142900 24500 143000 24600
rect 142900 24600 143000 24700
rect 142900 24700 143000 24800
rect 142900 24800 143000 24900
rect 142900 24900 143000 25000
rect 142900 35900 143000 36000
rect 142900 36000 143000 36100
rect 142900 36100 143000 36200
rect 142900 36200 143000 36300
rect 142900 36300 143000 36400
rect 142900 36400 143000 36500
rect 142900 36500 143000 36600
rect 142900 36600 143000 36700
rect 142900 36700 143000 36800
rect 142900 36800 143000 36900
rect 142900 36900 143000 37000
rect 142900 37000 143000 37100
rect 142900 37100 143000 37200
rect 142900 37200 143000 37300
rect 142900 37300 143000 37400
rect 142900 37400 143000 37500
rect 142900 37500 143000 37600
rect 142900 37600 143000 37700
rect 142900 37700 143000 37800
rect 142900 37800 143000 37900
rect 142900 37900 143000 38000
rect 142900 38000 143000 38100
rect 142900 38100 143000 38200
rect 143000 22400 143100 22500
rect 143000 22500 143100 22600
rect 143000 22600 143100 22700
rect 143000 22700 143100 22800
rect 143000 22800 143100 22900
rect 143000 22900 143100 23000
rect 143000 23000 143100 23100
rect 143000 23100 143100 23200
rect 143000 23200 143100 23300
rect 143000 23300 143100 23400
rect 143000 23400 143100 23500
rect 143000 23500 143100 23600
rect 143000 23600 143100 23700
rect 143000 23700 143100 23800
rect 143000 23800 143100 23900
rect 143000 23900 143100 24000
rect 143000 24000 143100 24100
rect 143000 24100 143100 24200
rect 143000 24200 143100 24300
rect 143000 24300 143100 24400
rect 143000 24400 143100 24500
rect 143000 24500 143100 24600
rect 143000 24600 143100 24700
rect 143000 24700 143100 24800
rect 143000 24800 143100 24900
rect 143000 24900 143100 25000
rect 143000 25000 143100 25100
rect 143000 35800 143100 35900
rect 143000 35900 143100 36000
rect 143000 36000 143100 36100
rect 143000 36100 143100 36200
rect 143000 36200 143100 36300
rect 143000 36300 143100 36400
rect 143000 36400 143100 36500
rect 143000 36500 143100 36600
rect 143000 36600 143100 36700
rect 143000 36700 143100 36800
rect 143000 36800 143100 36900
rect 143000 36900 143100 37000
rect 143000 37000 143100 37100
rect 143000 37100 143100 37200
rect 143000 37200 143100 37300
rect 143000 37300 143100 37400
rect 143000 37400 143100 37500
rect 143000 37500 143100 37600
rect 143000 37600 143100 37700
rect 143000 37700 143100 37800
rect 143000 37800 143100 37900
rect 143000 37900 143100 38000
rect 143000 38000 143100 38100
rect 143100 22400 143200 22500
rect 143100 22500 143200 22600
rect 143100 22600 143200 22700
rect 143100 22700 143200 22800
rect 143100 22800 143200 22900
rect 143100 22900 143200 23000
rect 143100 23000 143200 23100
rect 143100 23100 143200 23200
rect 143100 23200 143200 23300
rect 143100 23300 143200 23400
rect 143100 23400 143200 23500
rect 143100 23500 143200 23600
rect 143100 23600 143200 23700
rect 143100 23700 143200 23800
rect 143100 23800 143200 23900
rect 143100 23900 143200 24000
rect 143100 24000 143200 24100
rect 143100 24100 143200 24200
rect 143100 24200 143200 24300
rect 143100 24300 143200 24400
rect 143100 24400 143200 24500
rect 143100 24500 143200 24600
rect 143100 24600 143200 24700
rect 143100 24700 143200 24800
rect 143100 24800 143200 24900
rect 143100 24900 143200 25000
rect 143100 25000 143200 25100
rect 143100 25100 143200 25200
rect 143100 35800 143200 35900
rect 143100 35900 143200 36000
rect 143100 36000 143200 36100
rect 143100 36100 143200 36200
rect 143100 36200 143200 36300
rect 143100 36300 143200 36400
rect 143100 36400 143200 36500
rect 143100 36500 143200 36600
rect 143100 36600 143200 36700
rect 143100 36700 143200 36800
rect 143100 36800 143200 36900
rect 143100 36900 143200 37000
rect 143100 37000 143200 37100
rect 143100 37100 143200 37200
rect 143100 37200 143200 37300
rect 143100 37300 143200 37400
rect 143100 37400 143200 37500
rect 143100 37500 143200 37600
rect 143100 37600 143200 37700
rect 143100 37700 143200 37800
rect 143100 37800 143200 37900
rect 143100 37900 143200 38000
rect 143100 38000 143200 38100
rect 143200 22500 143300 22600
rect 143200 22600 143300 22700
rect 143200 22700 143300 22800
rect 143200 22800 143300 22900
rect 143200 22900 143300 23000
rect 143200 23000 143300 23100
rect 143200 23100 143300 23200
rect 143200 23200 143300 23300
rect 143200 23300 143300 23400
rect 143200 23400 143300 23500
rect 143200 23500 143300 23600
rect 143200 23600 143300 23700
rect 143200 23700 143300 23800
rect 143200 23800 143300 23900
rect 143200 23900 143300 24000
rect 143200 24000 143300 24100
rect 143200 24100 143300 24200
rect 143200 24200 143300 24300
rect 143200 24300 143300 24400
rect 143200 24400 143300 24500
rect 143200 24500 143300 24600
rect 143200 24600 143300 24700
rect 143200 24700 143300 24800
rect 143200 24800 143300 24900
rect 143200 24900 143300 25000
rect 143200 25000 143300 25100
rect 143200 25100 143300 25200
rect 143200 25200 143300 25300
rect 143200 35700 143300 35800
rect 143200 35800 143300 35900
rect 143200 35900 143300 36000
rect 143200 36000 143300 36100
rect 143200 36100 143300 36200
rect 143200 36200 143300 36300
rect 143200 36300 143300 36400
rect 143200 36400 143300 36500
rect 143200 36500 143300 36600
rect 143200 36600 143300 36700
rect 143200 36700 143300 36800
rect 143200 36800 143300 36900
rect 143200 36900 143300 37000
rect 143200 37000 143300 37100
rect 143200 37100 143300 37200
rect 143200 37200 143300 37300
rect 143200 37300 143300 37400
rect 143200 37400 143300 37500
rect 143200 37500 143300 37600
rect 143200 37600 143300 37700
rect 143200 37700 143300 37800
rect 143200 37800 143300 37900
rect 143200 37900 143300 38000
rect 143200 38000 143300 38100
rect 143300 22600 143400 22700
rect 143300 22700 143400 22800
rect 143300 22800 143400 22900
rect 143300 22900 143400 23000
rect 143300 23000 143400 23100
rect 143300 23100 143400 23200
rect 143300 23200 143400 23300
rect 143300 23300 143400 23400
rect 143300 23400 143400 23500
rect 143300 23500 143400 23600
rect 143300 23600 143400 23700
rect 143300 23700 143400 23800
rect 143300 23800 143400 23900
rect 143300 23900 143400 24000
rect 143300 24000 143400 24100
rect 143300 24100 143400 24200
rect 143300 24200 143400 24300
rect 143300 24300 143400 24400
rect 143300 24400 143400 24500
rect 143300 24500 143400 24600
rect 143300 24600 143400 24700
rect 143300 24700 143400 24800
rect 143300 24800 143400 24900
rect 143300 24900 143400 25000
rect 143300 25000 143400 25100
rect 143300 25100 143400 25200
rect 143300 25200 143400 25300
rect 143300 25300 143400 25400
rect 143300 35600 143400 35700
rect 143300 35700 143400 35800
rect 143300 35800 143400 35900
rect 143300 35900 143400 36000
rect 143300 36000 143400 36100
rect 143300 36100 143400 36200
rect 143300 36200 143400 36300
rect 143300 36300 143400 36400
rect 143300 36400 143400 36500
rect 143300 36500 143400 36600
rect 143300 36600 143400 36700
rect 143300 36700 143400 36800
rect 143300 36800 143400 36900
rect 143300 36900 143400 37000
rect 143300 37000 143400 37100
rect 143300 37100 143400 37200
rect 143300 37200 143400 37300
rect 143300 37300 143400 37400
rect 143300 37400 143400 37500
rect 143300 37500 143400 37600
rect 143300 37600 143400 37700
rect 143300 37700 143400 37800
rect 143300 37800 143400 37900
rect 143300 37900 143400 38000
rect 143400 22600 143500 22700
rect 143400 22700 143500 22800
rect 143400 22800 143500 22900
rect 143400 22900 143500 23000
rect 143400 23000 143500 23100
rect 143400 23100 143500 23200
rect 143400 23200 143500 23300
rect 143400 23300 143500 23400
rect 143400 23400 143500 23500
rect 143400 23500 143500 23600
rect 143400 23600 143500 23700
rect 143400 23700 143500 23800
rect 143400 23800 143500 23900
rect 143400 23900 143500 24000
rect 143400 24000 143500 24100
rect 143400 24100 143500 24200
rect 143400 24200 143500 24300
rect 143400 24300 143500 24400
rect 143400 24400 143500 24500
rect 143400 24500 143500 24600
rect 143400 24600 143500 24700
rect 143400 24700 143500 24800
rect 143400 24800 143500 24900
rect 143400 24900 143500 25000
rect 143400 25000 143500 25100
rect 143400 25100 143500 25200
rect 143400 25200 143500 25300
rect 143400 25300 143500 25400
rect 143400 25400 143500 25500
rect 143400 25500 143500 25600
rect 143400 35600 143500 35700
rect 143400 35700 143500 35800
rect 143400 35800 143500 35900
rect 143400 35900 143500 36000
rect 143400 36000 143500 36100
rect 143400 36100 143500 36200
rect 143400 36200 143500 36300
rect 143400 36300 143500 36400
rect 143400 36400 143500 36500
rect 143400 36500 143500 36600
rect 143400 36600 143500 36700
rect 143400 36700 143500 36800
rect 143400 36800 143500 36900
rect 143400 36900 143500 37000
rect 143400 37000 143500 37100
rect 143400 37100 143500 37200
rect 143400 37200 143500 37300
rect 143400 37300 143500 37400
rect 143400 37400 143500 37500
rect 143400 37500 143500 37600
rect 143400 37600 143500 37700
rect 143400 37700 143500 37800
rect 143400 37800 143500 37900
rect 143400 37900 143500 38000
rect 143500 22700 143600 22800
rect 143500 22800 143600 22900
rect 143500 22900 143600 23000
rect 143500 23000 143600 23100
rect 143500 23100 143600 23200
rect 143500 23200 143600 23300
rect 143500 23300 143600 23400
rect 143500 23400 143600 23500
rect 143500 23500 143600 23600
rect 143500 23600 143600 23700
rect 143500 23700 143600 23800
rect 143500 23800 143600 23900
rect 143500 23900 143600 24000
rect 143500 24000 143600 24100
rect 143500 24100 143600 24200
rect 143500 24200 143600 24300
rect 143500 24300 143600 24400
rect 143500 24400 143600 24500
rect 143500 24500 143600 24600
rect 143500 24600 143600 24700
rect 143500 24700 143600 24800
rect 143500 24800 143600 24900
rect 143500 24900 143600 25000
rect 143500 25000 143600 25100
rect 143500 25100 143600 25200
rect 143500 25200 143600 25300
rect 143500 25300 143600 25400
rect 143500 25400 143600 25500
rect 143500 25500 143600 25600
rect 143500 25600 143600 25700
rect 143500 35500 143600 35600
rect 143500 35600 143600 35700
rect 143500 35700 143600 35800
rect 143500 35800 143600 35900
rect 143500 35900 143600 36000
rect 143500 36000 143600 36100
rect 143500 36100 143600 36200
rect 143500 36200 143600 36300
rect 143500 36300 143600 36400
rect 143500 36400 143600 36500
rect 143500 36500 143600 36600
rect 143500 36600 143600 36700
rect 143500 36700 143600 36800
rect 143500 36800 143600 36900
rect 143500 36900 143600 37000
rect 143500 37000 143600 37100
rect 143500 37100 143600 37200
rect 143500 37200 143600 37300
rect 143500 37300 143600 37400
rect 143500 37400 143600 37500
rect 143500 37500 143600 37600
rect 143500 37600 143600 37700
rect 143500 37700 143600 37800
rect 143500 37800 143600 37900
rect 143500 37900 143600 38000
rect 143600 22800 143700 22900
rect 143600 22900 143700 23000
rect 143600 23000 143700 23100
rect 143600 23100 143700 23200
rect 143600 23200 143700 23300
rect 143600 23300 143700 23400
rect 143600 23400 143700 23500
rect 143600 23500 143700 23600
rect 143600 23600 143700 23700
rect 143600 23700 143700 23800
rect 143600 23800 143700 23900
rect 143600 23900 143700 24000
rect 143600 24000 143700 24100
rect 143600 24100 143700 24200
rect 143600 24200 143700 24300
rect 143600 24300 143700 24400
rect 143600 24400 143700 24500
rect 143600 24500 143700 24600
rect 143600 24600 143700 24700
rect 143600 24700 143700 24800
rect 143600 24800 143700 24900
rect 143600 24900 143700 25000
rect 143600 25000 143700 25100
rect 143600 25100 143700 25200
rect 143600 25200 143700 25300
rect 143600 25300 143700 25400
rect 143600 25400 143700 25500
rect 143600 25500 143700 25600
rect 143600 25600 143700 25700
rect 143600 25700 143700 25800
rect 143600 25800 143700 25900
rect 143600 35400 143700 35500
rect 143600 35500 143700 35600
rect 143600 35600 143700 35700
rect 143600 35700 143700 35800
rect 143600 35800 143700 35900
rect 143600 35900 143700 36000
rect 143600 36000 143700 36100
rect 143600 36100 143700 36200
rect 143600 36200 143700 36300
rect 143600 36300 143700 36400
rect 143600 36400 143700 36500
rect 143600 36500 143700 36600
rect 143600 36600 143700 36700
rect 143600 36700 143700 36800
rect 143600 36800 143700 36900
rect 143600 36900 143700 37000
rect 143600 37000 143700 37100
rect 143600 37100 143700 37200
rect 143600 37200 143700 37300
rect 143600 37300 143700 37400
rect 143600 37400 143700 37500
rect 143600 37500 143700 37600
rect 143600 37600 143700 37700
rect 143600 37700 143700 37800
rect 143600 37800 143700 37900
rect 143700 22900 143800 23000
rect 143700 23000 143800 23100
rect 143700 23100 143800 23200
rect 143700 23200 143800 23300
rect 143700 23300 143800 23400
rect 143700 23400 143800 23500
rect 143700 23500 143800 23600
rect 143700 23600 143800 23700
rect 143700 23700 143800 23800
rect 143700 23800 143800 23900
rect 143700 23900 143800 24000
rect 143700 24000 143800 24100
rect 143700 24100 143800 24200
rect 143700 24200 143800 24300
rect 143700 24300 143800 24400
rect 143700 24400 143800 24500
rect 143700 24500 143800 24600
rect 143700 24600 143800 24700
rect 143700 24700 143800 24800
rect 143700 24800 143800 24900
rect 143700 24900 143800 25000
rect 143700 25000 143800 25100
rect 143700 25100 143800 25200
rect 143700 25200 143800 25300
rect 143700 25300 143800 25400
rect 143700 25400 143800 25500
rect 143700 25500 143800 25600
rect 143700 25600 143800 25700
rect 143700 25700 143800 25800
rect 143700 25800 143800 25900
rect 143700 25900 143800 26000
rect 143700 35300 143800 35400
rect 143700 35400 143800 35500
rect 143700 35500 143800 35600
rect 143700 35600 143800 35700
rect 143700 35700 143800 35800
rect 143700 35800 143800 35900
rect 143700 35900 143800 36000
rect 143700 36000 143800 36100
rect 143700 36100 143800 36200
rect 143700 36200 143800 36300
rect 143700 36300 143800 36400
rect 143700 36400 143800 36500
rect 143700 36500 143800 36600
rect 143700 36600 143800 36700
rect 143700 36700 143800 36800
rect 143700 36800 143800 36900
rect 143700 36900 143800 37000
rect 143700 37000 143800 37100
rect 143700 37100 143800 37200
rect 143700 37200 143800 37300
rect 143700 37300 143800 37400
rect 143700 37400 143800 37500
rect 143700 37500 143800 37600
rect 143700 37600 143800 37700
rect 143700 37700 143800 37800
rect 143700 37800 143800 37900
rect 143800 22900 143900 23000
rect 143800 23000 143900 23100
rect 143800 23100 143900 23200
rect 143800 23200 143900 23300
rect 143800 23300 143900 23400
rect 143800 23400 143900 23500
rect 143800 23500 143900 23600
rect 143800 23600 143900 23700
rect 143800 23700 143900 23800
rect 143800 23800 143900 23900
rect 143800 23900 143900 24000
rect 143800 24000 143900 24100
rect 143800 24100 143900 24200
rect 143800 24200 143900 24300
rect 143800 24300 143900 24400
rect 143800 24400 143900 24500
rect 143800 24500 143900 24600
rect 143800 24600 143900 24700
rect 143800 24700 143900 24800
rect 143800 24800 143900 24900
rect 143800 24900 143900 25000
rect 143800 25000 143900 25100
rect 143800 25100 143900 25200
rect 143800 25200 143900 25300
rect 143800 25300 143900 25400
rect 143800 25400 143900 25500
rect 143800 25500 143900 25600
rect 143800 25600 143900 25700
rect 143800 25700 143900 25800
rect 143800 25800 143900 25900
rect 143800 25900 143900 26000
rect 143800 26000 143900 26100
rect 143800 26100 143900 26200
rect 143800 35200 143900 35300
rect 143800 35300 143900 35400
rect 143800 35400 143900 35500
rect 143800 35500 143900 35600
rect 143800 35600 143900 35700
rect 143800 35700 143900 35800
rect 143800 35800 143900 35900
rect 143800 35900 143900 36000
rect 143800 36000 143900 36100
rect 143800 36100 143900 36200
rect 143800 36200 143900 36300
rect 143800 36300 143900 36400
rect 143800 36400 143900 36500
rect 143800 36500 143900 36600
rect 143800 36600 143900 36700
rect 143800 36700 143900 36800
rect 143800 36800 143900 36900
rect 143800 36900 143900 37000
rect 143800 37000 143900 37100
rect 143800 37100 143900 37200
rect 143800 37200 143900 37300
rect 143800 37300 143900 37400
rect 143800 37400 143900 37500
rect 143800 37500 143900 37600
rect 143800 37600 143900 37700
rect 143800 37700 143900 37800
rect 143900 23000 144000 23100
rect 143900 23100 144000 23200
rect 143900 23200 144000 23300
rect 143900 23300 144000 23400
rect 143900 23400 144000 23500
rect 143900 23500 144000 23600
rect 143900 23600 144000 23700
rect 143900 23700 144000 23800
rect 143900 23800 144000 23900
rect 143900 23900 144000 24000
rect 143900 24000 144000 24100
rect 143900 24100 144000 24200
rect 143900 24200 144000 24300
rect 143900 24300 144000 24400
rect 143900 24400 144000 24500
rect 143900 24500 144000 24600
rect 143900 24600 144000 24700
rect 143900 24700 144000 24800
rect 143900 24800 144000 24900
rect 143900 24900 144000 25000
rect 143900 25000 144000 25100
rect 143900 25100 144000 25200
rect 143900 25200 144000 25300
rect 143900 25300 144000 25400
rect 143900 25400 144000 25500
rect 143900 25500 144000 25600
rect 143900 25600 144000 25700
rect 143900 25700 144000 25800
rect 143900 25800 144000 25900
rect 143900 25900 144000 26000
rect 143900 26000 144000 26100
rect 143900 26100 144000 26200
rect 143900 26200 144000 26300
rect 143900 26300 144000 26400
rect 143900 35100 144000 35200
rect 143900 35200 144000 35300
rect 143900 35300 144000 35400
rect 143900 35400 144000 35500
rect 143900 35500 144000 35600
rect 143900 35600 144000 35700
rect 143900 35700 144000 35800
rect 143900 35800 144000 35900
rect 143900 35900 144000 36000
rect 143900 36000 144000 36100
rect 143900 36100 144000 36200
rect 143900 36200 144000 36300
rect 143900 36300 144000 36400
rect 143900 36400 144000 36500
rect 143900 36500 144000 36600
rect 143900 36600 144000 36700
rect 143900 36700 144000 36800
rect 143900 36800 144000 36900
rect 143900 36900 144000 37000
rect 143900 37000 144000 37100
rect 143900 37100 144000 37200
rect 143900 37200 144000 37300
rect 143900 37300 144000 37400
rect 143900 37400 144000 37500
rect 143900 37500 144000 37600
rect 143900 37600 144000 37700
rect 143900 37700 144000 37800
rect 144000 23100 144100 23200
rect 144000 23200 144100 23300
rect 144000 23300 144100 23400
rect 144000 23400 144100 23500
rect 144000 23500 144100 23600
rect 144000 23600 144100 23700
rect 144000 23700 144100 23800
rect 144000 23800 144100 23900
rect 144000 23900 144100 24000
rect 144000 24000 144100 24100
rect 144000 24100 144100 24200
rect 144000 24200 144100 24300
rect 144000 24300 144100 24400
rect 144000 24400 144100 24500
rect 144000 24500 144100 24600
rect 144000 24600 144100 24700
rect 144000 24700 144100 24800
rect 144000 24800 144100 24900
rect 144000 24900 144100 25000
rect 144000 25000 144100 25100
rect 144000 25100 144100 25200
rect 144000 25200 144100 25300
rect 144000 25300 144100 25400
rect 144000 25400 144100 25500
rect 144000 25500 144100 25600
rect 144000 25600 144100 25700
rect 144000 25700 144100 25800
rect 144000 25800 144100 25900
rect 144000 25900 144100 26000
rect 144000 26000 144100 26100
rect 144000 26100 144100 26200
rect 144000 26200 144100 26300
rect 144000 26300 144100 26400
rect 144000 26400 144100 26500
rect 144000 26500 144100 26600
rect 144000 34900 144100 35000
rect 144000 35000 144100 35100
rect 144000 35100 144100 35200
rect 144000 35200 144100 35300
rect 144000 35300 144100 35400
rect 144000 35400 144100 35500
rect 144000 35500 144100 35600
rect 144000 35600 144100 35700
rect 144000 35700 144100 35800
rect 144000 35800 144100 35900
rect 144000 35900 144100 36000
rect 144000 36000 144100 36100
rect 144000 36100 144100 36200
rect 144000 36200 144100 36300
rect 144000 36300 144100 36400
rect 144000 36400 144100 36500
rect 144000 36500 144100 36600
rect 144000 36600 144100 36700
rect 144000 36700 144100 36800
rect 144000 36800 144100 36900
rect 144000 36900 144100 37000
rect 144000 37000 144100 37100
rect 144000 37100 144100 37200
rect 144000 37200 144100 37300
rect 144000 37300 144100 37400
rect 144000 37400 144100 37500
rect 144000 37500 144100 37600
rect 144000 37600 144100 37700
rect 144100 23200 144200 23300
rect 144100 23300 144200 23400
rect 144100 23400 144200 23500
rect 144100 23500 144200 23600
rect 144100 23600 144200 23700
rect 144100 23700 144200 23800
rect 144100 23800 144200 23900
rect 144100 23900 144200 24000
rect 144100 24000 144200 24100
rect 144100 24100 144200 24200
rect 144100 24200 144200 24300
rect 144100 24300 144200 24400
rect 144100 24400 144200 24500
rect 144100 24500 144200 24600
rect 144100 24600 144200 24700
rect 144100 24700 144200 24800
rect 144100 24800 144200 24900
rect 144100 24900 144200 25000
rect 144100 25000 144200 25100
rect 144100 25100 144200 25200
rect 144100 25200 144200 25300
rect 144100 25300 144200 25400
rect 144100 25400 144200 25500
rect 144100 25500 144200 25600
rect 144100 25600 144200 25700
rect 144100 25700 144200 25800
rect 144100 25800 144200 25900
rect 144100 25900 144200 26000
rect 144100 26000 144200 26100
rect 144100 26100 144200 26200
rect 144100 26200 144200 26300
rect 144100 26300 144200 26400
rect 144100 26400 144200 26500
rect 144100 26500 144200 26600
rect 144100 26600 144200 26700
rect 144100 26700 144200 26800
rect 144100 34800 144200 34900
rect 144100 34900 144200 35000
rect 144100 35000 144200 35100
rect 144100 35100 144200 35200
rect 144100 35200 144200 35300
rect 144100 35300 144200 35400
rect 144100 35400 144200 35500
rect 144100 35500 144200 35600
rect 144100 35600 144200 35700
rect 144100 35700 144200 35800
rect 144100 35800 144200 35900
rect 144100 35900 144200 36000
rect 144100 36000 144200 36100
rect 144100 36100 144200 36200
rect 144100 36200 144200 36300
rect 144100 36300 144200 36400
rect 144100 36400 144200 36500
rect 144100 36500 144200 36600
rect 144100 36600 144200 36700
rect 144100 36700 144200 36800
rect 144100 36800 144200 36900
rect 144100 36900 144200 37000
rect 144100 37000 144200 37100
rect 144100 37100 144200 37200
rect 144100 37200 144200 37300
rect 144100 37300 144200 37400
rect 144100 37400 144200 37500
rect 144100 37500 144200 37600
rect 144100 37600 144200 37700
rect 144200 23300 144300 23400
rect 144200 23400 144300 23500
rect 144200 23500 144300 23600
rect 144200 23600 144300 23700
rect 144200 23700 144300 23800
rect 144200 23800 144300 23900
rect 144200 23900 144300 24000
rect 144200 24000 144300 24100
rect 144200 24100 144300 24200
rect 144200 24200 144300 24300
rect 144200 24300 144300 24400
rect 144200 24400 144300 24500
rect 144200 24500 144300 24600
rect 144200 24600 144300 24700
rect 144200 24700 144300 24800
rect 144200 24800 144300 24900
rect 144200 24900 144300 25000
rect 144200 25000 144300 25100
rect 144200 25100 144300 25200
rect 144200 25200 144300 25300
rect 144200 25300 144300 25400
rect 144200 25400 144300 25500
rect 144200 25500 144300 25600
rect 144200 25600 144300 25700
rect 144200 25700 144300 25800
rect 144200 25800 144300 25900
rect 144200 25900 144300 26000
rect 144200 26000 144300 26100
rect 144200 26100 144300 26200
rect 144200 26200 144300 26300
rect 144200 26300 144300 26400
rect 144200 26400 144300 26500
rect 144200 26500 144300 26600
rect 144200 26600 144300 26700
rect 144200 26700 144300 26800
rect 144200 26800 144300 26900
rect 144200 26900 144300 27000
rect 144200 34600 144300 34700
rect 144200 34700 144300 34800
rect 144200 34800 144300 34900
rect 144200 34900 144300 35000
rect 144200 35000 144300 35100
rect 144200 35100 144300 35200
rect 144200 35200 144300 35300
rect 144200 35300 144300 35400
rect 144200 35400 144300 35500
rect 144200 35500 144300 35600
rect 144200 35600 144300 35700
rect 144200 35700 144300 35800
rect 144200 35800 144300 35900
rect 144200 35900 144300 36000
rect 144200 36000 144300 36100
rect 144200 36100 144300 36200
rect 144200 36200 144300 36300
rect 144200 36300 144300 36400
rect 144200 36400 144300 36500
rect 144200 36500 144300 36600
rect 144200 36600 144300 36700
rect 144200 36700 144300 36800
rect 144200 36800 144300 36900
rect 144200 36900 144300 37000
rect 144200 37000 144300 37100
rect 144200 37100 144300 37200
rect 144200 37200 144300 37300
rect 144200 37300 144300 37400
rect 144200 37400 144300 37500
rect 144200 37500 144300 37600
rect 144300 23400 144400 23500
rect 144300 23500 144400 23600
rect 144300 23600 144400 23700
rect 144300 23700 144400 23800
rect 144300 23800 144400 23900
rect 144300 23900 144400 24000
rect 144300 24000 144400 24100
rect 144300 24100 144400 24200
rect 144300 24200 144400 24300
rect 144300 24300 144400 24400
rect 144300 24400 144400 24500
rect 144300 24500 144400 24600
rect 144300 24600 144400 24700
rect 144300 24700 144400 24800
rect 144300 24800 144400 24900
rect 144300 24900 144400 25000
rect 144300 25000 144400 25100
rect 144300 25100 144400 25200
rect 144300 25200 144400 25300
rect 144300 25300 144400 25400
rect 144300 25400 144400 25500
rect 144300 25500 144400 25600
rect 144300 25600 144400 25700
rect 144300 25700 144400 25800
rect 144300 25800 144400 25900
rect 144300 25900 144400 26000
rect 144300 26000 144400 26100
rect 144300 26100 144400 26200
rect 144300 26200 144400 26300
rect 144300 26300 144400 26400
rect 144300 26400 144400 26500
rect 144300 26500 144400 26600
rect 144300 26600 144400 26700
rect 144300 26700 144400 26800
rect 144300 26800 144400 26900
rect 144300 26900 144400 27000
rect 144300 27000 144400 27100
rect 144300 27100 144400 27200
rect 144300 27200 144400 27300
rect 144300 34400 144400 34500
rect 144300 34500 144400 34600
rect 144300 34600 144400 34700
rect 144300 34700 144400 34800
rect 144300 34800 144400 34900
rect 144300 34900 144400 35000
rect 144300 35000 144400 35100
rect 144300 35100 144400 35200
rect 144300 35200 144400 35300
rect 144300 35300 144400 35400
rect 144300 35400 144400 35500
rect 144300 35500 144400 35600
rect 144300 35600 144400 35700
rect 144300 35700 144400 35800
rect 144300 35800 144400 35900
rect 144300 35900 144400 36000
rect 144300 36000 144400 36100
rect 144300 36100 144400 36200
rect 144300 36200 144400 36300
rect 144300 36300 144400 36400
rect 144300 36400 144400 36500
rect 144300 36500 144400 36600
rect 144300 36600 144400 36700
rect 144300 36700 144400 36800
rect 144300 36800 144400 36900
rect 144300 36900 144400 37000
rect 144300 37000 144400 37100
rect 144300 37100 144400 37200
rect 144300 37200 144400 37300
rect 144300 37300 144400 37400
rect 144300 37400 144400 37500
rect 144300 37500 144400 37600
rect 144400 23500 144500 23600
rect 144400 23600 144500 23700
rect 144400 23700 144500 23800
rect 144400 23800 144500 23900
rect 144400 23900 144500 24000
rect 144400 24000 144500 24100
rect 144400 24100 144500 24200
rect 144400 24200 144500 24300
rect 144400 24300 144500 24400
rect 144400 24400 144500 24500
rect 144400 24500 144500 24600
rect 144400 24600 144500 24700
rect 144400 24700 144500 24800
rect 144400 24800 144500 24900
rect 144400 24900 144500 25000
rect 144400 25000 144500 25100
rect 144400 25100 144500 25200
rect 144400 25200 144500 25300
rect 144400 25300 144500 25400
rect 144400 25400 144500 25500
rect 144400 25500 144500 25600
rect 144400 25600 144500 25700
rect 144400 25700 144500 25800
rect 144400 25800 144500 25900
rect 144400 25900 144500 26000
rect 144400 26000 144500 26100
rect 144400 26100 144500 26200
rect 144400 26200 144500 26300
rect 144400 26300 144500 26400
rect 144400 26400 144500 26500
rect 144400 26500 144500 26600
rect 144400 26600 144500 26700
rect 144400 26700 144500 26800
rect 144400 26800 144500 26900
rect 144400 26900 144500 27000
rect 144400 27000 144500 27100
rect 144400 27100 144500 27200
rect 144400 27200 144500 27300
rect 144400 27300 144500 27400
rect 144400 27400 144500 27500
rect 144400 27500 144500 27600
rect 144400 34100 144500 34200
rect 144400 34200 144500 34300
rect 144400 34300 144500 34400
rect 144400 34400 144500 34500
rect 144400 34500 144500 34600
rect 144400 34600 144500 34700
rect 144400 34700 144500 34800
rect 144400 34800 144500 34900
rect 144400 34900 144500 35000
rect 144400 35000 144500 35100
rect 144400 35100 144500 35200
rect 144400 35200 144500 35300
rect 144400 35300 144500 35400
rect 144400 35400 144500 35500
rect 144400 35500 144500 35600
rect 144400 35600 144500 35700
rect 144400 35700 144500 35800
rect 144400 35800 144500 35900
rect 144400 35900 144500 36000
rect 144400 36000 144500 36100
rect 144400 36100 144500 36200
rect 144400 36200 144500 36300
rect 144400 36300 144500 36400
rect 144400 36400 144500 36500
rect 144400 36500 144500 36600
rect 144400 36600 144500 36700
rect 144400 36700 144500 36800
rect 144400 36800 144500 36900
rect 144400 36900 144500 37000
rect 144400 37000 144500 37100
rect 144400 37100 144500 37200
rect 144400 37200 144500 37300
rect 144400 37300 144500 37400
rect 144400 37400 144500 37500
rect 144500 23600 144600 23700
rect 144500 23700 144600 23800
rect 144500 23800 144600 23900
rect 144500 23900 144600 24000
rect 144500 24000 144600 24100
rect 144500 24100 144600 24200
rect 144500 24200 144600 24300
rect 144500 24300 144600 24400
rect 144500 24400 144600 24500
rect 144500 24500 144600 24600
rect 144500 24600 144600 24700
rect 144500 24700 144600 24800
rect 144500 24800 144600 24900
rect 144500 24900 144600 25000
rect 144500 25000 144600 25100
rect 144500 25100 144600 25200
rect 144500 25200 144600 25300
rect 144500 25300 144600 25400
rect 144500 25400 144600 25500
rect 144500 25500 144600 25600
rect 144500 25600 144600 25700
rect 144500 25700 144600 25800
rect 144500 25800 144600 25900
rect 144500 25900 144600 26000
rect 144500 26000 144600 26100
rect 144500 26100 144600 26200
rect 144500 26200 144600 26300
rect 144500 26300 144600 26400
rect 144500 26400 144600 26500
rect 144500 26500 144600 26600
rect 144500 26600 144600 26700
rect 144500 26700 144600 26800
rect 144500 26800 144600 26900
rect 144500 26900 144600 27000
rect 144500 27000 144600 27100
rect 144500 27100 144600 27200
rect 144500 27200 144600 27300
rect 144500 27300 144600 27400
rect 144500 27400 144600 27500
rect 144500 27500 144600 27600
rect 144500 27600 144600 27700
rect 144500 27700 144600 27800
rect 144500 27800 144600 27900
rect 144500 33900 144600 34000
rect 144500 34000 144600 34100
rect 144500 34100 144600 34200
rect 144500 34200 144600 34300
rect 144500 34300 144600 34400
rect 144500 34400 144600 34500
rect 144500 34500 144600 34600
rect 144500 34600 144600 34700
rect 144500 34700 144600 34800
rect 144500 34800 144600 34900
rect 144500 34900 144600 35000
rect 144500 35000 144600 35100
rect 144500 35100 144600 35200
rect 144500 35200 144600 35300
rect 144500 35300 144600 35400
rect 144500 35400 144600 35500
rect 144500 35500 144600 35600
rect 144500 35600 144600 35700
rect 144500 35700 144600 35800
rect 144500 35800 144600 35900
rect 144500 35900 144600 36000
rect 144500 36000 144600 36100
rect 144500 36100 144600 36200
rect 144500 36200 144600 36300
rect 144500 36300 144600 36400
rect 144500 36400 144600 36500
rect 144500 36500 144600 36600
rect 144500 36600 144600 36700
rect 144500 36700 144600 36800
rect 144500 36800 144600 36900
rect 144500 36900 144600 37000
rect 144500 37000 144600 37100
rect 144500 37100 144600 37200
rect 144500 37200 144600 37300
rect 144500 37300 144600 37400
rect 144600 23700 144700 23800
rect 144600 23800 144700 23900
rect 144600 23900 144700 24000
rect 144600 24000 144700 24100
rect 144600 24100 144700 24200
rect 144600 24200 144700 24300
rect 144600 24300 144700 24400
rect 144600 24400 144700 24500
rect 144600 24500 144700 24600
rect 144600 24600 144700 24700
rect 144600 24700 144700 24800
rect 144600 24800 144700 24900
rect 144600 24900 144700 25000
rect 144600 25000 144700 25100
rect 144600 25100 144700 25200
rect 144600 25200 144700 25300
rect 144600 25300 144700 25400
rect 144600 25400 144700 25500
rect 144600 25500 144700 25600
rect 144600 25600 144700 25700
rect 144600 25700 144700 25800
rect 144600 25800 144700 25900
rect 144600 25900 144700 26000
rect 144600 26000 144700 26100
rect 144600 26100 144700 26200
rect 144600 26200 144700 26300
rect 144600 26300 144700 26400
rect 144600 26400 144700 26500
rect 144600 26500 144700 26600
rect 144600 26600 144700 26700
rect 144600 26700 144700 26800
rect 144600 26800 144700 26900
rect 144600 26900 144700 27000
rect 144600 27000 144700 27100
rect 144600 27100 144700 27200
rect 144600 27200 144700 27300
rect 144600 27300 144700 27400
rect 144600 27400 144700 27500
rect 144600 27500 144700 27600
rect 144600 27600 144700 27700
rect 144600 27700 144700 27800
rect 144600 27800 144700 27900
rect 144600 27900 144700 28000
rect 144600 28000 144700 28100
rect 144600 28100 144700 28200
rect 144600 33500 144700 33600
rect 144600 33600 144700 33700
rect 144600 33700 144700 33800
rect 144600 33800 144700 33900
rect 144600 33900 144700 34000
rect 144600 34000 144700 34100
rect 144600 34100 144700 34200
rect 144600 34200 144700 34300
rect 144600 34300 144700 34400
rect 144600 34400 144700 34500
rect 144600 34500 144700 34600
rect 144600 34600 144700 34700
rect 144600 34700 144700 34800
rect 144600 34800 144700 34900
rect 144600 34900 144700 35000
rect 144600 35000 144700 35100
rect 144600 35100 144700 35200
rect 144600 35200 144700 35300
rect 144600 35300 144700 35400
rect 144600 35400 144700 35500
rect 144600 35500 144700 35600
rect 144600 35600 144700 35700
rect 144600 35700 144700 35800
rect 144600 35800 144700 35900
rect 144600 35900 144700 36000
rect 144600 36000 144700 36100
rect 144600 36100 144700 36200
rect 144600 36200 144700 36300
rect 144600 36300 144700 36400
rect 144600 36400 144700 36500
rect 144600 36500 144700 36600
rect 144600 36600 144700 36700
rect 144600 36700 144700 36800
rect 144600 36800 144700 36900
rect 144600 36900 144700 37000
rect 144600 37000 144700 37100
rect 144600 37100 144700 37200
rect 144600 37200 144700 37300
rect 144600 37300 144700 37400
rect 144700 23900 144800 24000
rect 144700 24000 144800 24100
rect 144700 24100 144800 24200
rect 144700 24200 144800 24300
rect 144700 24300 144800 24400
rect 144700 24400 144800 24500
rect 144700 24500 144800 24600
rect 144700 24600 144800 24700
rect 144700 24700 144800 24800
rect 144700 24800 144800 24900
rect 144700 24900 144800 25000
rect 144700 25000 144800 25100
rect 144700 25100 144800 25200
rect 144700 25200 144800 25300
rect 144700 25300 144800 25400
rect 144700 25400 144800 25500
rect 144700 25500 144800 25600
rect 144700 25600 144800 25700
rect 144700 25700 144800 25800
rect 144700 25800 144800 25900
rect 144700 25900 144800 26000
rect 144700 26000 144800 26100
rect 144700 26100 144800 26200
rect 144700 26200 144800 26300
rect 144700 26300 144800 26400
rect 144700 26400 144800 26500
rect 144700 26500 144800 26600
rect 144700 26600 144800 26700
rect 144700 26700 144800 26800
rect 144700 26800 144800 26900
rect 144700 26900 144800 27000
rect 144700 27000 144800 27100
rect 144700 27100 144800 27200
rect 144700 27200 144800 27300
rect 144700 27300 144800 27400
rect 144700 27400 144800 27500
rect 144700 27500 144800 27600
rect 144700 27600 144800 27700
rect 144700 27700 144800 27800
rect 144700 27800 144800 27900
rect 144700 27900 144800 28000
rect 144700 28000 144800 28100
rect 144700 28100 144800 28200
rect 144700 28200 144800 28300
rect 144700 28300 144800 28400
rect 144700 28400 144800 28500
rect 144700 28500 144800 28600
rect 144700 33100 144800 33200
rect 144700 33200 144800 33300
rect 144700 33300 144800 33400
rect 144700 33400 144800 33500
rect 144700 33500 144800 33600
rect 144700 33600 144800 33700
rect 144700 33700 144800 33800
rect 144700 33800 144800 33900
rect 144700 33900 144800 34000
rect 144700 34000 144800 34100
rect 144700 34100 144800 34200
rect 144700 34200 144800 34300
rect 144700 34300 144800 34400
rect 144700 34400 144800 34500
rect 144700 34500 144800 34600
rect 144700 34600 144800 34700
rect 144700 34700 144800 34800
rect 144700 34800 144800 34900
rect 144700 34900 144800 35000
rect 144700 35000 144800 35100
rect 144700 35100 144800 35200
rect 144700 35200 144800 35300
rect 144700 35300 144800 35400
rect 144700 35400 144800 35500
rect 144700 35500 144800 35600
rect 144700 35600 144800 35700
rect 144700 35700 144800 35800
rect 144700 35800 144800 35900
rect 144700 35900 144800 36000
rect 144700 36000 144800 36100
rect 144700 36100 144800 36200
rect 144700 36200 144800 36300
rect 144700 36300 144800 36400
rect 144700 36400 144800 36500
rect 144700 36500 144800 36600
rect 144700 36600 144800 36700
rect 144700 36700 144800 36800
rect 144700 36800 144800 36900
rect 144700 36900 144800 37000
rect 144700 37000 144800 37100
rect 144700 37100 144800 37200
rect 144700 37200 144800 37300
rect 144800 24000 144900 24100
rect 144800 24100 144900 24200
rect 144800 24200 144900 24300
rect 144800 24300 144900 24400
rect 144800 24400 144900 24500
rect 144800 24500 144900 24600
rect 144800 24600 144900 24700
rect 144800 24700 144900 24800
rect 144800 24800 144900 24900
rect 144800 24900 144900 25000
rect 144800 25000 144900 25100
rect 144800 25100 144900 25200
rect 144800 25200 144900 25300
rect 144800 25300 144900 25400
rect 144800 25400 144900 25500
rect 144800 25500 144900 25600
rect 144800 25600 144900 25700
rect 144800 25700 144900 25800
rect 144800 25800 144900 25900
rect 144800 25900 144900 26000
rect 144800 26000 144900 26100
rect 144800 26100 144900 26200
rect 144800 26200 144900 26300
rect 144800 26300 144900 26400
rect 144800 26400 144900 26500
rect 144800 26500 144900 26600
rect 144800 26600 144900 26700
rect 144800 26700 144900 26800
rect 144800 26800 144900 26900
rect 144800 26900 144900 27000
rect 144800 27000 144900 27100
rect 144800 27100 144900 27200
rect 144800 27200 144900 27300
rect 144800 27300 144900 27400
rect 144800 27400 144900 27500
rect 144800 27500 144900 27600
rect 144800 27600 144900 27700
rect 144800 27700 144900 27800
rect 144800 27800 144900 27900
rect 144800 27900 144900 28000
rect 144800 28000 144900 28100
rect 144800 28100 144900 28200
rect 144800 28200 144900 28300
rect 144800 28300 144900 28400
rect 144800 28400 144900 28500
rect 144800 28500 144900 28600
rect 144800 28600 144900 28700
rect 144800 28700 144900 28800
rect 144800 28800 144900 28900
rect 144800 28900 144900 29000
rect 144800 29000 144900 29100
rect 144800 32600 144900 32700
rect 144800 32700 144900 32800
rect 144800 32800 144900 32900
rect 144800 32900 144900 33000
rect 144800 33000 144900 33100
rect 144800 33100 144900 33200
rect 144800 33200 144900 33300
rect 144800 33300 144900 33400
rect 144800 33400 144900 33500
rect 144800 33500 144900 33600
rect 144800 33600 144900 33700
rect 144800 33700 144900 33800
rect 144800 33800 144900 33900
rect 144800 33900 144900 34000
rect 144800 34000 144900 34100
rect 144800 34100 144900 34200
rect 144800 34200 144900 34300
rect 144800 34300 144900 34400
rect 144800 34400 144900 34500
rect 144800 34500 144900 34600
rect 144800 34600 144900 34700
rect 144800 34700 144900 34800
rect 144800 34800 144900 34900
rect 144800 34900 144900 35000
rect 144800 35000 144900 35100
rect 144800 35100 144900 35200
rect 144800 35200 144900 35300
rect 144800 35300 144900 35400
rect 144800 35400 144900 35500
rect 144800 35500 144900 35600
rect 144800 35600 144900 35700
rect 144800 35700 144900 35800
rect 144800 35800 144900 35900
rect 144800 35900 144900 36000
rect 144800 36000 144900 36100
rect 144800 36100 144900 36200
rect 144800 36200 144900 36300
rect 144800 36300 144900 36400
rect 144800 36400 144900 36500
rect 144800 36500 144900 36600
rect 144800 36600 144900 36700
rect 144800 36700 144900 36800
rect 144800 36800 144900 36900
rect 144800 36900 144900 37000
rect 144800 37000 144900 37100
rect 144800 37100 144900 37200
rect 144900 24100 145000 24200
rect 144900 24200 145000 24300
rect 144900 24300 145000 24400
rect 144900 24400 145000 24500
rect 144900 24500 145000 24600
rect 144900 24600 145000 24700
rect 144900 24700 145000 24800
rect 144900 24800 145000 24900
rect 144900 24900 145000 25000
rect 144900 25000 145000 25100
rect 144900 25100 145000 25200
rect 144900 25200 145000 25300
rect 144900 25300 145000 25400
rect 144900 25400 145000 25500
rect 144900 25500 145000 25600
rect 144900 25600 145000 25700
rect 144900 25700 145000 25800
rect 144900 25800 145000 25900
rect 144900 25900 145000 26000
rect 144900 26000 145000 26100
rect 144900 26100 145000 26200
rect 144900 26200 145000 26300
rect 144900 26300 145000 26400
rect 144900 26400 145000 26500
rect 144900 26500 145000 26600
rect 144900 26600 145000 26700
rect 144900 26700 145000 26800
rect 144900 26800 145000 26900
rect 144900 26900 145000 27000
rect 144900 27000 145000 27100
rect 144900 27100 145000 27200
rect 144900 27200 145000 27300
rect 144900 27300 145000 27400
rect 144900 27400 145000 27500
rect 144900 27500 145000 27600
rect 144900 27600 145000 27700
rect 144900 27700 145000 27800
rect 144900 27800 145000 27900
rect 144900 27900 145000 28000
rect 144900 28000 145000 28100
rect 144900 28100 145000 28200
rect 144900 28200 145000 28300
rect 144900 28300 145000 28400
rect 144900 28400 145000 28500
rect 144900 28500 145000 28600
rect 144900 28600 145000 28700
rect 144900 28700 145000 28800
rect 144900 28800 145000 28900
rect 144900 28900 145000 29000
rect 144900 29000 145000 29100
rect 144900 29100 145000 29200
rect 144900 29200 145000 29300
rect 144900 29300 145000 29400
rect 144900 29400 145000 29500
rect 144900 29500 145000 29600
rect 144900 29600 145000 29700
rect 144900 29700 145000 29800
rect 144900 31800 145000 31900
rect 144900 31900 145000 32000
rect 144900 32000 145000 32100
rect 144900 32100 145000 32200
rect 144900 32200 145000 32300
rect 144900 32300 145000 32400
rect 144900 32400 145000 32500
rect 144900 32500 145000 32600
rect 144900 32600 145000 32700
rect 144900 32700 145000 32800
rect 144900 32800 145000 32900
rect 144900 32900 145000 33000
rect 144900 33000 145000 33100
rect 144900 33100 145000 33200
rect 144900 33200 145000 33300
rect 144900 33300 145000 33400
rect 144900 33400 145000 33500
rect 144900 33500 145000 33600
rect 144900 33600 145000 33700
rect 144900 33700 145000 33800
rect 144900 33800 145000 33900
rect 144900 33900 145000 34000
rect 144900 34000 145000 34100
rect 144900 34100 145000 34200
rect 144900 34200 145000 34300
rect 144900 34300 145000 34400
rect 144900 34400 145000 34500
rect 144900 34500 145000 34600
rect 144900 34600 145000 34700
rect 144900 34700 145000 34800
rect 144900 34800 145000 34900
rect 144900 34900 145000 35000
rect 144900 35000 145000 35100
rect 144900 35100 145000 35200
rect 144900 35200 145000 35300
rect 144900 35300 145000 35400
rect 144900 35400 145000 35500
rect 144900 35500 145000 35600
rect 144900 35600 145000 35700
rect 144900 35700 145000 35800
rect 144900 35800 145000 35900
rect 144900 35900 145000 36000
rect 144900 36000 145000 36100
rect 144900 36100 145000 36200
rect 144900 36200 145000 36300
rect 144900 36300 145000 36400
rect 144900 36400 145000 36500
rect 144900 36500 145000 36600
rect 144900 36600 145000 36700
rect 144900 36700 145000 36800
rect 144900 36800 145000 36900
rect 144900 36900 145000 37000
rect 144900 37000 145000 37100
rect 145000 24200 145100 24300
rect 145000 24300 145100 24400
rect 145000 24400 145100 24500
rect 145000 24500 145100 24600
rect 145000 24600 145100 24700
rect 145000 24700 145100 24800
rect 145000 24800 145100 24900
rect 145000 24900 145100 25000
rect 145000 25000 145100 25100
rect 145000 25100 145100 25200
rect 145000 25200 145100 25300
rect 145000 25300 145100 25400
rect 145000 25400 145100 25500
rect 145000 25500 145100 25600
rect 145000 25600 145100 25700
rect 145000 25700 145100 25800
rect 145000 25800 145100 25900
rect 145000 25900 145100 26000
rect 145000 26000 145100 26100
rect 145000 26100 145100 26200
rect 145000 26200 145100 26300
rect 145000 26300 145100 26400
rect 145000 26400 145100 26500
rect 145000 26500 145100 26600
rect 145000 26600 145100 26700
rect 145000 26700 145100 26800
rect 145000 26800 145100 26900
rect 145000 26900 145100 27000
rect 145000 27000 145100 27100
rect 145000 27100 145100 27200
rect 145000 27200 145100 27300
rect 145000 27300 145100 27400
rect 145000 27400 145100 27500
rect 145000 27500 145100 27600
rect 145000 27600 145100 27700
rect 145000 27700 145100 27800
rect 145000 27800 145100 27900
rect 145000 27900 145100 28000
rect 145000 28000 145100 28100
rect 145000 28100 145100 28200
rect 145000 28200 145100 28300
rect 145000 28300 145100 28400
rect 145000 28400 145100 28500
rect 145000 28500 145100 28600
rect 145000 28600 145100 28700
rect 145000 28700 145100 28800
rect 145000 28800 145100 28900
rect 145000 28900 145100 29000
rect 145000 29000 145100 29100
rect 145000 29100 145100 29200
rect 145000 29200 145100 29300
rect 145000 29300 145100 29400
rect 145000 29400 145100 29500
rect 145000 29500 145100 29600
rect 145000 29600 145100 29700
rect 145000 29700 145100 29800
rect 145000 29800 145100 29900
rect 145000 29900 145100 30000
rect 145000 30000 145100 30100
rect 145000 30100 145100 30200
rect 145000 30200 145100 30300
rect 145000 30300 145100 30400
rect 145000 30400 145100 30500
rect 145000 30500 145100 30600
rect 145000 30600 145100 30700
rect 145000 30700 145100 30800
rect 145000 30800 145100 30900
rect 145000 30900 145100 31000
rect 145000 31000 145100 31100
rect 145000 31100 145100 31200
rect 145000 31200 145100 31300
rect 145000 31300 145100 31400
rect 145000 31400 145100 31500
rect 145000 31500 145100 31600
rect 145000 31600 145100 31700
rect 145000 31700 145100 31800
rect 145000 31800 145100 31900
rect 145000 31900 145100 32000
rect 145000 32000 145100 32100
rect 145000 32100 145100 32200
rect 145000 32200 145100 32300
rect 145000 32300 145100 32400
rect 145000 32400 145100 32500
rect 145000 32500 145100 32600
rect 145000 32600 145100 32700
rect 145000 32700 145100 32800
rect 145000 32800 145100 32900
rect 145000 32900 145100 33000
rect 145000 33000 145100 33100
rect 145000 33100 145100 33200
rect 145000 33200 145100 33300
rect 145000 33300 145100 33400
rect 145000 33400 145100 33500
rect 145000 33500 145100 33600
rect 145000 33600 145100 33700
rect 145000 33700 145100 33800
rect 145000 33800 145100 33900
rect 145000 33900 145100 34000
rect 145000 34000 145100 34100
rect 145000 34100 145100 34200
rect 145000 34200 145100 34300
rect 145000 34300 145100 34400
rect 145000 34400 145100 34500
rect 145000 34500 145100 34600
rect 145000 34600 145100 34700
rect 145000 34700 145100 34800
rect 145000 34800 145100 34900
rect 145000 34900 145100 35000
rect 145000 35000 145100 35100
rect 145000 35100 145100 35200
rect 145000 35200 145100 35300
rect 145000 35300 145100 35400
rect 145000 35400 145100 35500
rect 145000 35500 145100 35600
rect 145000 35600 145100 35700
rect 145000 35700 145100 35800
rect 145000 35800 145100 35900
rect 145000 35900 145100 36000
rect 145000 36000 145100 36100
rect 145000 36100 145100 36200
rect 145000 36200 145100 36300
rect 145000 36300 145100 36400
rect 145000 36400 145100 36500
rect 145000 36500 145100 36600
rect 145000 36600 145100 36700
rect 145000 36700 145100 36800
rect 145000 36800 145100 36900
rect 145000 36900 145100 37000
rect 145100 24400 145200 24500
rect 145100 24500 145200 24600
rect 145100 24600 145200 24700
rect 145100 24700 145200 24800
rect 145100 24800 145200 24900
rect 145100 24900 145200 25000
rect 145100 25000 145200 25100
rect 145100 25100 145200 25200
rect 145100 25200 145200 25300
rect 145100 25300 145200 25400
rect 145100 25400 145200 25500
rect 145100 25500 145200 25600
rect 145100 25600 145200 25700
rect 145100 25700 145200 25800
rect 145100 25800 145200 25900
rect 145100 25900 145200 26000
rect 145100 26000 145200 26100
rect 145100 26100 145200 26200
rect 145100 26200 145200 26300
rect 145100 26300 145200 26400
rect 145100 26400 145200 26500
rect 145100 26500 145200 26600
rect 145100 26600 145200 26700
rect 145100 26700 145200 26800
rect 145100 26800 145200 26900
rect 145100 26900 145200 27000
rect 145100 27000 145200 27100
rect 145100 27100 145200 27200
rect 145100 27200 145200 27300
rect 145100 27300 145200 27400
rect 145100 27400 145200 27500
rect 145100 27500 145200 27600
rect 145100 27600 145200 27700
rect 145100 27700 145200 27800
rect 145100 27800 145200 27900
rect 145100 27900 145200 28000
rect 145100 28000 145200 28100
rect 145100 28100 145200 28200
rect 145100 28200 145200 28300
rect 145100 28300 145200 28400
rect 145100 28400 145200 28500
rect 145100 28500 145200 28600
rect 145100 28600 145200 28700
rect 145100 28700 145200 28800
rect 145100 28800 145200 28900
rect 145100 28900 145200 29000
rect 145100 29000 145200 29100
rect 145100 29100 145200 29200
rect 145100 29200 145200 29300
rect 145100 29300 145200 29400
rect 145100 29400 145200 29500
rect 145100 29500 145200 29600
rect 145100 29600 145200 29700
rect 145100 29700 145200 29800
rect 145100 29800 145200 29900
rect 145100 29900 145200 30000
rect 145100 30000 145200 30100
rect 145100 30100 145200 30200
rect 145100 30200 145200 30300
rect 145100 30300 145200 30400
rect 145100 30400 145200 30500
rect 145100 30500 145200 30600
rect 145100 30600 145200 30700
rect 145100 30700 145200 30800
rect 145100 30800 145200 30900
rect 145100 30900 145200 31000
rect 145100 31000 145200 31100
rect 145100 31100 145200 31200
rect 145100 31200 145200 31300
rect 145100 31300 145200 31400
rect 145100 31400 145200 31500
rect 145100 31500 145200 31600
rect 145100 31600 145200 31700
rect 145100 31700 145200 31800
rect 145100 31800 145200 31900
rect 145100 31900 145200 32000
rect 145100 32000 145200 32100
rect 145100 32100 145200 32200
rect 145100 32200 145200 32300
rect 145100 32300 145200 32400
rect 145100 32400 145200 32500
rect 145100 32500 145200 32600
rect 145100 32600 145200 32700
rect 145100 32700 145200 32800
rect 145100 32800 145200 32900
rect 145100 32900 145200 33000
rect 145100 33000 145200 33100
rect 145100 33100 145200 33200
rect 145100 33200 145200 33300
rect 145100 33300 145200 33400
rect 145100 33400 145200 33500
rect 145100 33500 145200 33600
rect 145100 33600 145200 33700
rect 145100 33700 145200 33800
rect 145100 33800 145200 33900
rect 145100 33900 145200 34000
rect 145100 34000 145200 34100
rect 145100 34100 145200 34200
rect 145100 34200 145200 34300
rect 145100 34300 145200 34400
rect 145100 34400 145200 34500
rect 145100 34500 145200 34600
rect 145100 34600 145200 34700
rect 145100 34700 145200 34800
rect 145100 34800 145200 34900
rect 145100 34900 145200 35000
rect 145100 35000 145200 35100
rect 145100 35100 145200 35200
rect 145100 35200 145200 35300
rect 145100 35300 145200 35400
rect 145100 35400 145200 35500
rect 145100 35500 145200 35600
rect 145100 35600 145200 35700
rect 145100 35700 145200 35800
rect 145100 35800 145200 35900
rect 145100 35900 145200 36000
rect 145100 36000 145200 36100
rect 145100 36100 145200 36200
rect 145100 36200 145200 36300
rect 145100 36300 145200 36400
rect 145100 36400 145200 36500
rect 145100 36500 145200 36600
rect 145100 36600 145200 36700
rect 145100 36700 145200 36800
rect 145100 36800 145200 36900
rect 145200 24500 145300 24600
rect 145200 24600 145300 24700
rect 145200 24700 145300 24800
rect 145200 24800 145300 24900
rect 145200 24900 145300 25000
rect 145200 25000 145300 25100
rect 145200 25100 145300 25200
rect 145200 25200 145300 25300
rect 145200 25300 145300 25400
rect 145200 25400 145300 25500
rect 145200 25500 145300 25600
rect 145200 25600 145300 25700
rect 145200 25700 145300 25800
rect 145200 25800 145300 25900
rect 145200 25900 145300 26000
rect 145200 26000 145300 26100
rect 145200 26100 145300 26200
rect 145200 26200 145300 26300
rect 145200 26300 145300 26400
rect 145200 26400 145300 26500
rect 145200 26500 145300 26600
rect 145200 26600 145300 26700
rect 145200 26700 145300 26800
rect 145200 26800 145300 26900
rect 145200 26900 145300 27000
rect 145200 27000 145300 27100
rect 145200 27100 145300 27200
rect 145200 27200 145300 27300
rect 145200 27300 145300 27400
rect 145200 27400 145300 27500
rect 145200 27500 145300 27600
rect 145200 27600 145300 27700
rect 145200 27700 145300 27800
rect 145200 27800 145300 27900
rect 145200 27900 145300 28000
rect 145200 28000 145300 28100
rect 145200 28100 145300 28200
rect 145200 28200 145300 28300
rect 145200 28300 145300 28400
rect 145200 28400 145300 28500
rect 145200 28500 145300 28600
rect 145200 28600 145300 28700
rect 145200 28700 145300 28800
rect 145200 28800 145300 28900
rect 145200 28900 145300 29000
rect 145200 29000 145300 29100
rect 145200 29100 145300 29200
rect 145200 29200 145300 29300
rect 145200 29300 145300 29400
rect 145200 29400 145300 29500
rect 145200 29500 145300 29600
rect 145200 29600 145300 29700
rect 145200 29700 145300 29800
rect 145200 29800 145300 29900
rect 145200 29900 145300 30000
rect 145200 30000 145300 30100
rect 145200 30100 145300 30200
rect 145200 30200 145300 30300
rect 145200 30300 145300 30400
rect 145200 30400 145300 30500
rect 145200 30500 145300 30600
rect 145200 30600 145300 30700
rect 145200 30700 145300 30800
rect 145200 30800 145300 30900
rect 145200 30900 145300 31000
rect 145200 31000 145300 31100
rect 145200 31100 145300 31200
rect 145200 31200 145300 31300
rect 145200 31300 145300 31400
rect 145200 31400 145300 31500
rect 145200 31500 145300 31600
rect 145200 31600 145300 31700
rect 145200 31700 145300 31800
rect 145200 31800 145300 31900
rect 145200 31900 145300 32000
rect 145200 32000 145300 32100
rect 145200 32100 145300 32200
rect 145200 32200 145300 32300
rect 145200 32300 145300 32400
rect 145200 32400 145300 32500
rect 145200 32500 145300 32600
rect 145200 32600 145300 32700
rect 145200 32700 145300 32800
rect 145200 32800 145300 32900
rect 145200 32900 145300 33000
rect 145200 33000 145300 33100
rect 145200 33100 145300 33200
rect 145200 33200 145300 33300
rect 145200 33300 145300 33400
rect 145200 33400 145300 33500
rect 145200 33500 145300 33600
rect 145200 33600 145300 33700
rect 145200 33700 145300 33800
rect 145200 33800 145300 33900
rect 145200 33900 145300 34000
rect 145200 34000 145300 34100
rect 145200 34100 145300 34200
rect 145200 34200 145300 34300
rect 145200 34300 145300 34400
rect 145200 34400 145300 34500
rect 145200 34500 145300 34600
rect 145200 34600 145300 34700
rect 145200 34700 145300 34800
rect 145200 34800 145300 34900
rect 145200 34900 145300 35000
rect 145200 35000 145300 35100
rect 145200 35100 145300 35200
rect 145200 35200 145300 35300
rect 145200 35300 145300 35400
rect 145200 35400 145300 35500
rect 145200 35500 145300 35600
rect 145200 35600 145300 35700
rect 145200 35700 145300 35800
rect 145200 35800 145300 35900
rect 145200 35900 145300 36000
rect 145200 36000 145300 36100
rect 145200 36100 145300 36200
rect 145200 36200 145300 36300
rect 145200 36300 145300 36400
rect 145200 36400 145300 36500
rect 145200 36500 145300 36600
rect 145200 36600 145300 36700
rect 145200 36700 145300 36800
rect 145300 24700 145400 24800
rect 145300 24800 145400 24900
rect 145300 24900 145400 25000
rect 145300 25000 145400 25100
rect 145300 25100 145400 25200
rect 145300 25200 145400 25300
rect 145300 25300 145400 25400
rect 145300 25400 145400 25500
rect 145300 25500 145400 25600
rect 145300 25600 145400 25700
rect 145300 25700 145400 25800
rect 145300 25800 145400 25900
rect 145300 25900 145400 26000
rect 145300 26000 145400 26100
rect 145300 26100 145400 26200
rect 145300 26200 145400 26300
rect 145300 26300 145400 26400
rect 145300 26400 145400 26500
rect 145300 26500 145400 26600
rect 145300 26600 145400 26700
rect 145300 26700 145400 26800
rect 145300 26800 145400 26900
rect 145300 26900 145400 27000
rect 145300 27000 145400 27100
rect 145300 27100 145400 27200
rect 145300 27200 145400 27300
rect 145300 27300 145400 27400
rect 145300 27400 145400 27500
rect 145300 27500 145400 27600
rect 145300 27600 145400 27700
rect 145300 27700 145400 27800
rect 145300 27800 145400 27900
rect 145300 27900 145400 28000
rect 145300 28000 145400 28100
rect 145300 28100 145400 28200
rect 145300 28200 145400 28300
rect 145300 28300 145400 28400
rect 145300 28400 145400 28500
rect 145300 28500 145400 28600
rect 145300 28600 145400 28700
rect 145300 28700 145400 28800
rect 145300 28800 145400 28900
rect 145300 28900 145400 29000
rect 145300 29000 145400 29100
rect 145300 29100 145400 29200
rect 145300 29200 145400 29300
rect 145300 29300 145400 29400
rect 145300 29400 145400 29500
rect 145300 29500 145400 29600
rect 145300 29600 145400 29700
rect 145300 29700 145400 29800
rect 145300 29800 145400 29900
rect 145300 29900 145400 30000
rect 145300 30000 145400 30100
rect 145300 30100 145400 30200
rect 145300 30200 145400 30300
rect 145300 30300 145400 30400
rect 145300 30400 145400 30500
rect 145300 30500 145400 30600
rect 145300 30600 145400 30700
rect 145300 30700 145400 30800
rect 145300 30800 145400 30900
rect 145300 30900 145400 31000
rect 145300 31000 145400 31100
rect 145300 31100 145400 31200
rect 145300 31200 145400 31300
rect 145300 31300 145400 31400
rect 145300 31400 145400 31500
rect 145300 31500 145400 31600
rect 145300 31600 145400 31700
rect 145300 31700 145400 31800
rect 145300 31800 145400 31900
rect 145300 31900 145400 32000
rect 145300 32000 145400 32100
rect 145300 32100 145400 32200
rect 145300 32200 145400 32300
rect 145300 32300 145400 32400
rect 145300 32400 145400 32500
rect 145300 32500 145400 32600
rect 145300 32600 145400 32700
rect 145300 32700 145400 32800
rect 145300 32800 145400 32900
rect 145300 32900 145400 33000
rect 145300 33000 145400 33100
rect 145300 33100 145400 33200
rect 145300 33200 145400 33300
rect 145300 33300 145400 33400
rect 145300 33400 145400 33500
rect 145300 33500 145400 33600
rect 145300 33600 145400 33700
rect 145300 33700 145400 33800
rect 145300 33800 145400 33900
rect 145300 33900 145400 34000
rect 145300 34000 145400 34100
rect 145300 34100 145400 34200
rect 145300 34200 145400 34300
rect 145300 34300 145400 34400
rect 145300 34400 145400 34500
rect 145300 34500 145400 34600
rect 145300 34600 145400 34700
rect 145300 34700 145400 34800
rect 145300 34800 145400 34900
rect 145300 34900 145400 35000
rect 145300 35000 145400 35100
rect 145300 35100 145400 35200
rect 145300 35200 145400 35300
rect 145300 35300 145400 35400
rect 145300 35400 145400 35500
rect 145300 35500 145400 35600
rect 145300 35600 145400 35700
rect 145300 35700 145400 35800
rect 145300 35800 145400 35900
rect 145300 35900 145400 36000
rect 145300 36000 145400 36100
rect 145300 36100 145400 36200
rect 145300 36200 145400 36300
rect 145300 36300 145400 36400
rect 145300 36400 145400 36500
rect 145300 36500 145400 36600
rect 145300 36600 145400 36700
rect 145400 24900 145500 25000
rect 145400 25000 145500 25100
rect 145400 25100 145500 25200
rect 145400 25200 145500 25300
rect 145400 25300 145500 25400
rect 145400 25400 145500 25500
rect 145400 25500 145500 25600
rect 145400 25600 145500 25700
rect 145400 25700 145500 25800
rect 145400 25800 145500 25900
rect 145400 25900 145500 26000
rect 145400 26000 145500 26100
rect 145400 26100 145500 26200
rect 145400 26200 145500 26300
rect 145400 26300 145500 26400
rect 145400 26400 145500 26500
rect 145400 26500 145500 26600
rect 145400 26600 145500 26700
rect 145400 26700 145500 26800
rect 145400 26800 145500 26900
rect 145400 26900 145500 27000
rect 145400 27000 145500 27100
rect 145400 27100 145500 27200
rect 145400 27200 145500 27300
rect 145400 27300 145500 27400
rect 145400 27400 145500 27500
rect 145400 27500 145500 27600
rect 145400 27600 145500 27700
rect 145400 27700 145500 27800
rect 145400 27800 145500 27900
rect 145400 27900 145500 28000
rect 145400 28000 145500 28100
rect 145400 28100 145500 28200
rect 145400 28200 145500 28300
rect 145400 28300 145500 28400
rect 145400 28400 145500 28500
rect 145400 28500 145500 28600
rect 145400 28600 145500 28700
rect 145400 28700 145500 28800
rect 145400 28800 145500 28900
rect 145400 28900 145500 29000
rect 145400 29000 145500 29100
rect 145400 29100 145500 29200
rect 145400 29200 145500 29300
rect 145400 29300 145500 29400
rect 145400 29400 145500 29500
rect 145400 29500 145500 29600
rect 145400 29600 145500 29700
rect 145400 29700 145500 29800
rect 145400 29800 145500 29900
rect 145400 29900 145500 30000
rect 145400 30000 145500 30100
rect 145400 30100 145500 30200
rect 145400 30200 145500 30300
rect 145400 30300 145500 30400
rect 145400 30400 145500 30500
rect 145400 30500 145500 30600
rect 145400 30600 145500 30700
rect 145400 30700 145500 30800
rect 145400 30800 145500 30900
rect 145400 30900 145500 31000
rect 145400 31000 145500 31100
rect 145400 31100 145500 31200
rect 145400 31200 145500 31300
rect 145400 31300 145500 31400
rect 145400 31400 145500 31500
rect 145400 31500 145500 31600
rect 145400 31600 145500 31700
rect 145400 31700 145500 31800
rect 145400 31800 145500 31900
rect 145400 31900 145500 32000
rect 145400 32000 145500 32100
rect 145400 32100 145500 32200
rect 145400 32200 145500 32300
rect 145400 32300 145500 32400
rect 145400 32400 145500 32500
rect 145400 32500 145500 32600
rect 145400 32600 145500 32700
rect 145400 32700 145500 32800
rect 145400 32800 145500 32900
rect 145400 32900 145500 33000
rect 145400 33000 145500 33100
rect 145400 33100 145500 33200
rect 145400 33200 145500 33300
rect 145400 33300 145500 33400
rect 145400 33400 145500 33500
rect 145400 33500 145500 33600
rect 145400 33600 145500 33700
rect 145400 33700 145500 33800
rect 145400 33800 145500 33900
rect 145400 33900 145500 34000
rect 145400 34000 145500 34100
rect 145400 34100 145500 34200
rect 145400 34200 145500 34300
rect 145400 34300 145500 34400
rect 145400 34400 145500 34500
rect 145400 34500 145500 34600
rect 145400 34600 145500 34700
rect 145400 34700 145500 34800
rect 145400 34800 145500 34900
rect 145400 34900 145500 35000
rect 145400 35000 145500 35100
rect 145400 35100 145500 35200
rect 145400 35200 145500 35300
rect 145400 35300 145500 35400
rect 145400 35400 145500 35500
rect 145400 35500 145500 35600
rect 145400 35600 145500 35700
rect 145400 35700 145500 35800
rect 145400 35800 145500 35900
rect 145400 35900 145500 36000
rect 145400 36000 145500 36100
rect 145400 36100 145500 36200
rect 145400 36200 145500 36300
rect 145400 36300 145500 36400
rect 145400 36400 145500 36500
rect 145400 36500 145500 36600
rect 145500 25000 145600 25100
rect 145500 25100 145600 25200
rect 145500 25200 145600 25300
rect 145500 25300 145600 25400
rect 145500 25400 145600 25500
rect 145500 25500 145600 25600
rect 145500 25600 145600 25700
rect 145500 25700 145600 25800
rect 145500 25800 145600 25900
rect 145500 25900 145600 26000
rect 145500 26000 145600 26100
rect 145500 26100 145600 26200
rect 145500 26200 145600 26300
rect 145500 26300 145600 26400
rect 145500 26400 145600 26500
rect 145500 26500 145600 26600
rect 145500 26600 145600 26700
rect 145500 26700 145600 26800
rect 145500 26800 145600 26900
rect 145500 26900 145600 27000
rect 145500 27000 145600 27100
rect 145500 27100 145600 27200
rect 145500 27200 145600 27300
rect 145500 27300 145600 27400
rect 145500 27400 145600 27500
rect 145500 27500 145600 27600
rect 145500 27600 145600 27700
rect 145500 27700 145600 27800
rect 145500 27800 145600 27900
rect 145500 27900 145600 28000
rect 145500 28000 145600 28100
rect 145500 28100 145600 28200
rect 145500 28200 145600 28300
rect 145500 28300 145600 28400
rect 145500 28400 145600 28500
rect 145500 28500 145600 28600
rect 145500 28600 145600 28700
rect 145500 28700 145600 28800
rect 145500 28800 145600 28900
rect 145500 28900 145600 29000
rect 145500 29000 145600 29100
rect 145500 29100 145600 29200
rect 145500 29200 145600 29300
rect 145500 29300 145600 29400
rect 145500 29400 145600 29500
rect 145500 29500 145600 29600
rect 145500 29600 145600 29700
rect 145500 29700 145600 29800
rect 145500 29800 145600 29900
rect 145500 29900 145600 30000
rect 145500 30000 145600 30100
rect 145500 30100 145600 30200
rect 145500 30200 145600 30300
rect 145500 30300 145600 30400
rect 145500 30400 145600 30500
rect 145500 30500 145600 30600
rect 145500 30600 145600 30700
rect 145500 30700 145600 30800
rect 145500 30800 145600 30900
rect 145500 30900 145600 31000
rect 145500 31000 145600 31100
rect 145500 31100 145600 31200
rect 145500 31200 145600 31300
rect 145500 31300 145600 31400
rect 145500 31400 145600 31500
rect 145500 31500 145600 31600
rect 145500 31600 145600 31700
rect 145500 31700 145600 31800
rect 145500 31800 145600 31900
rect 145500 31900 145600 32000
rect 145500 32000 145600 32100
rect 145500 32100 145600 32200
rect 145500 32200 145600 32300
rect 145500 32300 145600 32400
rect 145500 32400 145600 32500
rect 145500 32500 145600 32600
rect 145500 32600 145600 32700
rect 145500 32700 145600 32800
rect 145500 32800 145600 32900
rect 145500 32900 145600 33000
rect 145500 33000 145600 33100
rect 145500 33100 145600 33200
rect 145500 33200 145600 33300
rect 145500 33300 145600 33400
rect 145500 33400 145600 33500
rect 145500 33500 145600 33600
rect 145500 33600 145600 33700
rect 145500 33700 145600 33800
rect 145500 33800 145600 33900
rect 145500 33900 145600 34000
rect 145500 34000 145600 34100
rect 145500 34100 145600 34200
rect 145500 34200 145600 34300
rect 145500 34300 145600 34400
rect 145500 34400 145600 34500
rect 145500 34500 145600 34600
rect 145500 34600 145600 34700
rect 145500 34700 145600 34800
rect 145500 34800 145600 34900
rect 145500 34900 145600 35000
rect 145500 35000 145600 35100
rect 145500 35100 145600 35200
rect 145500 35200 145600 35300
rect 145500 35300 145600 35400
rect 145500 35400 145600 35500
rect 145500 35500 145600 35600
rect 145500 35600 145600 35700
rect 145500 35700 145600 35800
rect 145500 35800 145600 35900
rect 145500 35900 145600 36000
rect 145500 36000 145600 36100
rect 145500 36100 145600 36200
rect 145500 36200 145600 36300
rect 145500 36300 145600 36400
rect 145600 25200 145700 25300
rect 145600 25300 145700 25400
rect 145600 25400 145700 25500
rect 145600 25500 145700 25600
rect 145600 25600 145700 25700
rect 145600 25700 145700 25800
rect 145600 25800 145700 25900
rect 145600 25900 145700 26000
rect 145600 26000 145700 26100
rect 145600 26100 145700 26200
rect 145600 26200 145700 26300
rect 145600 26300 145700 26400
rect 145600 26400 145700 26500
rect 145600 26500 145700 26600
rect 145600 26600 145700 26700
rect 145600 26700 145700 26800
rect 145600 26800 145700 26900
rect 145600 26900 145700 27000
rect 145600 27000 145700 27100
rect 145600 27100 145700 27200
rect 145600 27200 145700 27300
rect 145600 27300 145700 27400
rect 145600 27400 145700 27500
rect 145600 27500 145700 27600
rect 145600 27600 145700 27700
rect 145600 27700 145700 27800
rect 145600 27800 145700 27900
rect 145600 27900 145700 28000
rect 145600 28000 145700 28100
rect 145600 28100 145700 28200
rect 145600 28200 145700 28300
rect 145600 28300 145700 28400
rect 145600 28400 145700 28500
rect 145600 28500 145700 28600
rect 145600 28600 145700 28700
rect 145600 28700 145700 28800
rect 145600 28800 145700 28900
rect 145600 28900 145700 29000
rect 145600 29000 145700 29100
rect 145600 29100 145700 29200
rect 145600 29200 145700 29300
rect 145600 29300 145700 29400
rect 145600 29400 145700 29500
rect 145600 29500 145700 29600
rect 145600 29600 145700 29700
rect 145600 29700 145700 29800
rect 145600 29800 145700 29900
rect 145600 29900 145700 30000
rect 145600 30000 145700 30100
rect 145600 30100 145700 30200
rect 145600 30200 145700 30300
rect 145600 30300 145700 30400
rect 145600 30400 145700 30500
rect 145600 30500 145700 30600
rect 145600 30600 145700 30700
rect 145600 30700 145700 30800
rect 145600 30800 145700 30900
rect 145600 30900 145700 31000
rect 145600 31000 145700 31100
rect 145600 31100 145700 31200
rect 145600 31200 145700 31300
rect 145600 31300 145700 31400
rect 145600 31400 145700 31500
rect 145600 31500 145700 31600
rect 145600 31600 145700 31700
rect 145600 31700 145700 31800
rect 145600 31800 145700 31900
rect 145600 31900 145700 32000
rect 145600 32000 145700 32100
rect 145600 32100 145700 32200
rect 145600 32200 145700 32300
rect 145600 32300 145700 32400
rect 145600 32400 145700 32500
rect 145600 32500 145700 32600
rect 145600 32600 145700 32700
rect 145600 32700 145700 32800
rect 145600 32800 145700 32900
rect 145600 32900 145700 33000
rect 145600 33000 145700 33100
rect 145600 33100 145700 33200
rect 145600 33200 145700 33300
rect 145600 33300 145700 33400
rect 145600 33400 145700 33500
rect 145600 33500 145700 33600
rect 145600 33600 145700 33700
rect 145600 33700 145700 33800
rect 145600 33800 145700 33900
rect 145600 33900 145700 34000
rect 145600 34000 145700 34100
rect 145600 34100 145700 34200
rect 145600 34200 145700 34300
rect 145600 34300 145700 34400
rect 145600 34400 145700 34500
rect 145600 34500 145700 34600
rect 145600 34600 145700 34700
rect 145600 34700 145700 34800
rect 145600 34800 145700 34900
rect 145600 34900 145700 35000
rect 145600 35000 145700 35100
rect 145600 35100 145700 35200
rect 145600 35200 145700 35300
rect 145600 35300 145700 35400
rect 145600 35400 145700 35500
rect 145600 35500 145700 35600
rect 145600 35600 145700 35700
rect 145600 35700 145700 35800
rect 145600 35800 145700 35900
rect 145600 35900 145700 36000
rect 145600 36000 145700 36100
rect 145600 36100 145700 36200
rect 145600 36200 145700 36300
rect 145700 25400 145800 25500
rect 145700 25500 145800 25600
rect 145700 25600 145800 25700
rect 145700 25700 145800 25800
rect 145700 25800 145800 25900
rect 145700 25900 145800 26000
rect 145700 26000 145800 26100
rect 145700 26100 145800 26200
rect 145700 26200 145800 26300
rect 145700 26300 145800 26400
rect 145700 26400 145800 26500
rect 145700 26500 145800 26600
rect 145700 26600 145800 26700
rect 145700 26700 145800 26800
rect 145700 26800 145800 26900
rect 145700 26900 145800 27000
rect 145700 27000 145800 27100
rect 145700 27100 145800 27200
rect 145700 27200 145800 27300
rect 145700 27300 145800 27400
rect 145700 27400 145800 27500
rect 145700 27500 145800 27600
rect 145700 27600 145800 27700
rect 145700 27700 145800 27800
rect 145700 27800 145800 27900
rect 145700 27900 145800 28000
rect 145700 28000 145800 28100
rect 145700 28100 145800 28200
rect 145700 28200 145800 28300
rect 145700 28300 145800 28400
rect 145700 28400 145800 28500
rect 145700 28500 145800 28600
rect 145700 28600 145800 28700
rect 145700 28700 145800 28800
rect 145700 28800 145800 28900
rect 145700 28900 145800 29000
rect 145700 29000 145800 29100
rect 145700 29100 145800 29200
rect 145700 29200 145800 29300
rect 145700 29300 145800 29400
rect 145700 29400 145800 29500
rect 145700 29500 145800 29600
rect 145700 29600 145800 29700
rect 145700 29700 145800 29800
rect 145700 29800 145800 29900
rect 145700 29900 145800 30000
rect 145700 30000 145800 30100
rect 145700 30100 145800 30200
rect 145700 30200 145800 30300
rect 145700 30300 145800 30400
rect 145700 30400 145800 30500
rect 145700 30500 145800 30600
rect 145700 30600 145800 30700
rect 145700 30700 145800 30800
rect 145700 30800 145800 30900
rect 145700 30900 145800 31000
rect 145700 31000 145800 31100
rect 145700 31100 145800 31200
rect 145700 31200 145800 31300
rect 145700 31300 145800 31400
rect 145700 31400 145800 31500
rect 145700 31500 145800 31600
rect 145700 31600 145800 31700
rect 145700 31700 145800 31800
rect 145700 31800 145800 31900
rect 145700 31900 145800 32000
rect 145700 32000 145800 32100
rect 145700 32100 145800 32200
rect 145700 32200 145800 32300
rect 145700 32300 145800 32400
rect 145700 32400 145800 32500
rect 145700 32500 145800 32600
rect 145700 32600 145800 32700
rect 145700 32700 145800 32800
rect 145700 32800 145800 32900
rect 145700 32900 145800 33000
rect 145700 33000 145800 33100
rect 145700 33100 145800 33200
rect 145700 33200 145800 33300
rect 145700 33300 145800 33400
rect 145700 33400 145800 33500
rect 145700 33500 145800 33600
rect 145700 33600 145800 33700
rect 145700 33700 145800 33800
rect 145700 33800 145800 33900
rect 145700 33900 145800 34000
rect 145700 34000 145800 34100
rect 145700 34100 145800 34200
rect 145700 34200 145800 34300
rect 145700 34300 145800 34400
rect 145700 34400 145800 34500
rect 145700 34500 145800 34600
rect 145700 34600 145800 34700
rect 145700 34700 145800 34800
rect 145700 34800 145800 34900
rect 145700 34900 145800 35000
rect 145700 35000 145800 35100
rect 145700 35100 145800 35200
rect 145700 35200 145800 35300
rect 145700 35300 145800 35400
rect 145700 35400 145800 35500
rect 145700 35500 145800 35600
rect 145700 35600 145800 35700
rect 145700 35700 145800 35800
rect 145700 35800 145800 35900
rect 145700 35900 145800 36000
rect 145700 36000 145800 36100
rect 145800 25600 145900 25700
rect 145800 25700 145900 25800
rect 145800 25800 145900 25900
rect 145800 25900 145900 26000
rect 145800 26000 145900 26100
rect 145800 26100 145900 26200
rect 145800 26200 145900 26300
rect 145800 26300 145900 26400
rect 145800 26400 145900 26500
rect 145800 26500 145900 26600
rect 145800 26600 145900 26700
rect 145800 26700 145900 26800
rect 145800 26800 145900 26900
rect 145800 26900 145900 27000
rect 145800 27000 145900 27100
rect 145800 27100 145900 27200
rect 145800 27200 145900 27300
rect 145800 27300 145900 27400
rect 145800 27400 145900 27500
rect 145800 27500 145900 27600
rect 145800 27600 145900 27700
rect 145800 27700 145900 27800
rect 145800 27800 145900 27900
rect 145800 27900 145900 28000
rect 145800 28000 145900 28100
rect 145800 28100 145900 28200
rect 145800 28200 145900 28300
rect 145800 28300 145900 28400
rect 145800 28400 145900 28500
rect 145800 28500 145900 28600
rect 145800 28600 145900 28700
rect 145800 28700 145900 28800
rect 145800 28800 145900 28900
rect 145800 28900 145900 29000
rect 145800 29000 145900 29100
rect 145800 29100 145900 29200
rect 145800 29200 145900 29300
rect 145800 29300 145900 29400
rect 145800 29400 145900 29500
rect 145800 29500 145900 29600
rect 145800 29600 145900 29700
rect 145800 29700 145900 29800
rect 145800 29800 145900 29900
rect 145800 29900 145900 30000
rect 145800 30000 145900 30100
rect 145800 30100 145900 30200
rect 145800 30200 145900 30300
rect 145800 30300 145900 30400
rect 145800 30400 145900 30500
rect 145800 30500 145900 30600
rect 145800 30600 145900 30700
rect 145800 30700 145900 30800
rect 145800 30800 145900 30900
rect 145800 30900 145900 31000
rect 145800 31000 145900 31100
rect 145800 31100 145900 31200
rect 145800 31200 145900 31300
rect 145800 31300 145900 31400
rect 145800 31400 145900 31500
rect 145800 31500 145900 31600
rect 145800 31600 145900 31700
rect 145800 31700 145900 31800
rect 145800 31800 145900 31900
rect 145800 31900 145900 32000
rect 145800 32000 145900 32100
rect 145800 32100 145900 32200
rect 145800 32200 145900 32300
rect 145800 32300 145900 32400
rect 145800 32400 145900 32500
rect 145800 32500 145900 32600
rect 145800 32600 145900 32700
rect 145800 32700 145900 32800
rect 145800 32800 145900 32900
rect 145800 32900 145900 33000
rect 145800 33000 145900 33100
rect 145800 33100 145900 33200
rect 145800 33200 145900 33300
rect 145800 33300 145900 33400
rect 145800 33400 145900 33500
rect 145800 33500 145900 33600
rect 145800 33600 145900 33700
rect 145800 33700 145900 33800
rect 145800 33800 145900 33900
rect 145800 33900 145900 34000
rect 145800 34000 145900 34100
rect 145800 34100 145900 34200
rect 145800 34200 145900 34300
rect 145800 34300 145900 34400
rect 145800 34400 145900 34500
rect 145800 34500 145900 34600
rect 145800 34600 145900 34700
rect 145800 34700 145900 34800
rect 145800 34800 145900 34900
rect 145800 34900 145900 35000
rect 145800 35000 145900 35100
rect 145800 35100 145900 35200
rect 145800 35200 145900 35300
rect 145800 35300 145900 35400
rect 145800 35400 145900 35500
rect 145800 35500 145900 35600
rect 145800 35600 145900 35700
rect 145800 35700 145900 35800
rect 145800 35800 145900 35900
rect 145800 35900 145900 36000
rect 145900 25800 146000 25900
rect 145900 25900 146000 26000
rect 145900 26000 146000 26100
rect 145900 26100 146000 26200
rect 145900 26200 146000 26300
rect 145900 26300 146000 26400
rect 145900 26400 146000 26500
rect 145900 26500 146000 26600
rect 145900 26600 146000 26700
rect 145900 26700 146000 26800
rect 145900 26800 146000 26900
rect 145900 26900 146000 27000
rect 145900 27000 146000 27100
rect 145900 27100 146000 27200
rect 145900 27200 146000 27300
rect 145900 27300 146000 27400
rect 145900 27400 146000 27500
rect 145900 27500 146000 27600
rect 145900 27600 146000 27700
rect 145900 27700 146000 27800
rect 145900 27800 146000 27900
rect 145900 27900 146000 28000
rect 145900 28000 146000 28100
rect 145900 28100 146000 28200
rect 145900 28200 146000 28300
rect 145900 28300 146000 28400
rect 145900 28400 146000 28500
rect 145900 28500 146000 28600
rect 145900 28600 146000 28700
rect 145900 28700 146000 28800
rect 145900 28800 146000 28900
rect 145900 28900 146000 29000
rect 145900 29000 146000 29100
rect 145900 29100 146000 29200
rect 145900 29200 146000 29300
rect 145900 29300 146000 29400
rect 145900 29400 146000 29500
rect 145900 29500 146000 29600
rect 145900 29600 146000 29700
rect 145900 29700 146000 29800
rect 145900 29800 146000 29900
rect 145900 29900 146000 30000
rect 145900 30000 146000 30100
rect 145900 30100 146000 30200
rect 145900 30200 146000 30300
rect 145900 30300 146000 30400
rect 145900 30400 146000 30500
rect 145900 30500 146000 30600
rect 145900 30600 146000 30700
rect 145900 30700 146000 30800
rect 145900 30800 146000 30900
rect 145900 30900 146000 31000
rect 145900 31000 146000 31100
rect 145900 31100 146000 31200
rect 145900 31200 146000 31300
rect 145900 31300 146000 31400
rect 145900 31400 146000 31500
rect 145900 31500 146000 31600
rect 145900 31600 146000 31700
rect 145900 31700 146000 31800
rect 145900 31800 146000 31900
rect 145900 31900 146000 32000
rect 145900 32000 146000 32100
rect 145900 32100 146000 32200
rect 145900 32200 146000 32300
rect 145900 32300 146000 32400
rect 145900 32400 146000 32500
rect 145900 32500 146000 32600
rect 145900 32600 146000 32700
rect 145900 32700 146000 32800
rect 145900 32800 146000 32900
rect 145900 32900 146000 33000
rect 145900 33000 146000 33100
rect 145900 33100 146000 33200
rect 145900 33200 146000 33300
rect 145900 33300 146000 33400
rect 145900 33400 146000 33500
rect 145900 33500 146000 33600
rect 145900 33600 146000 33700
rect 145900 33700 146000 33800
rect 145900 33800 146000 33900
rect 145900 33900 146000 34000
rect 145900 34000 146000 34100
rect 145900 34100 146000 34200
rect 145900 34200 146000 34300
rect 145900 34300 146000 34400
rect 145900 34400 146000 34500
rect 145900 34500 146000 34600
rect 145900 34600 146000 34700
rect 145900 34700 146000 34800
rect 145900 34800 146000 34900
rect 145900 34900 146000 35000
rect 145900 35000 146000 35100
rect 145900 35100 146000 35200
rect 145900 35200 146000 35300
rect 145900 35300 146000 35400
rect 145900 35400 146000 35500
rect 145900 35500 146000 35600
rect 145900 35600 146000 35700
rect 145900 35700 146000 35800
rect 146000 26100 146100 26200
rect 146000 26200 146100 26300
rect 146000 26300 146100 26400
rect 146000 26400 146100 26500
rect 146000 26500 146100 26600
rect 146000 26600 146100 26700
rect 146000 26700 146100 26800
rect 146000 26800 146100 26900
rect 146000 26900 146100 27000
rect 146000 27000 146100 27100
rect 146000 27100 146100 27200
rect 146000 27200 146100 27300
rect 146000 27300 146100 27400
rect 146000 27400 146100 27500
rect 146000 27500 146100 27600
rect 146000 27600 146100 27700
rect 146000 27700 146100 27800
rect 146000 27800 146100 27900
rect 146000 27900 146100 28000
rect 146000 28000 146100 28100
rect 146000 28100 146100 28200
rect 146000 28200 146100 28300
rect 146000 28300 146100 28400
rect 146000 28400 146100 28500
rect 146000 28500 146100 28600
rect 146000 28600 146100 28700
rect 146000 28700 146100 28800
rect 146000 28800 146100 28900
rect 146000 28900 146100 29000
rect 146000 29000 146100 29100
rect 146000 29100 146100 29200
rect 146000 29200 146100 29300
rect 146000 29300 146100 29400
rect 146000 29400 146100 29500
rect 146000 29500 146100 29600
rect 146000 29600 146100 29700
rect 146000 29700 146100 29800
rect 146000 29800 146100 29900
rect 146000 29900 146100 30000
rect 146000 30000 146100 30100
rect 146000 30100 146100 30200
rect 146000 30200 146100 30300
rect 146000 30300 146100 30400
rect 146000 30400 146100 30500
rect 146000 30500 146100 30600
rect 146000 30600 146100 30700
rect 146000 30700 146100 30800
rect 146000 30800 146100 30900
rect 146000 30900 146100 31000
rect 146000 31000 146100 31100
rect 146000 31100 146100 31200
rect 146000 31200 146100 31300
rect 146000 31300 146100 31400
rect 146000 31400 146100 31500
rect 146000 31500 146100 31600
rect 146000 31600 146100 31700
rect 146000 31700 146100 31800
rect 146000 31800 146100 31900
rect 146000 31900 146100 32000
rect 146000 32000 146100 32100
rect 146000 32100 146100 32200
rect 146000 32200 146100 32300
rect 146000 32300 146100 32400
rect 146000 32400 146100 32500
rect 146000 32500 146100 32600
rect 146000 32600 146100 32700
rect 146000 32700 146100 32800
rect 146000 32800 146100 32900
rect 146000 32900 146100 33000
rect 146000 33000 146100 33100
rect 146000 33100 146100 33200
rect 146000 33200 146100 33300
rect 146000 33300 146100 33400
rect 146000 33400 146100 33500
rect 146000 33500 146100 33600
rect 146000 33600 146100 33700
rect 146000 33700 146100 33800
rect 146000 33800 146100 33900
rect 146000 33900 146100 34000
rect 146000 34000 146100 34100
rect 146000 34100 146100 34200
rect 146000 34200 146100 34300
rect 146000 34300 146100 34400
rect 146000 34400 146100 34500
rect 146000 34500 146100 34600
rect 146000 34600 146100 34700
rect 146000 34700 146100 34800
rect 146000 34800 146100 34900
rect 146000 34900 146100 35000
rect 146000 35000 146100 35100
rect 146000 35100 146100 35200
rect 146000 35200 146100 35300
rect 146000 35300 146100 35400
rect 146000 35400 146100 35500
rect 146000 35500 146100 35600
rect 146100 26300 146200 26400
rect 146100 26400 146200 26500
rect 146100 26500 146200 26600
rect 146100 26600 146200 26700
rect 146100 26700 146200 26800
rect 146100 26800 146200 26900
rect 146100 26900 146200 27000
rect 146100 27000 146200 27100
rect 146100 27100 146200 27200
rect 146100 27200 146200 27300
rect 146100 27300 146200 27400
rect 146100 27400 146200 27500
rect 146100 27500 146200 27600
rect 146100 27600 146200 27700
rect 146100 27700 146200 27800
rect 146100 27800 146200 27900
rect 146100 27900 146200 28000
rect 146100 28000 146200 28100
rect 146100 28100 146200 28200
rect 146100 28200 146200 28300
rect 146100 28300 146200 28400
rect 146100 28400 146200 28500
rect 146100 28500 146200 28600
rect 146100 28600 146200 28700
rect 146100 28700 146200 28800
rect 146100 28800 146200 28900
rect 146100 28900 146200 29000
rect 146100 29000 146200 29100
rect 146100 29100 146200 29200
rect 146100 29200 146200 29300
rect 146100 29300 146200 29400
rect 146100 29400 146200 29500
rect 146100 29500 146200 29600
rect 146100 29600 146200 29700
rect 146100 29700 146200 29800
rect 146100 29800 146200 29900
rect 146100 29900 146200 30000
rect 146100 30000 146200 30100
rect 146100 30100 146200 30200
rect 146100 30200 146200 30300
rect 146100 30300 146200 30400
rect 146100 30400 146200 30500
rect 146100 30500 146200 30600
rect 146100 30600 146200 30700
rect 146100 30700 146200 30800
rect 146100 30800 146200 30900
rect 146100 30900 146200 31000
rect 146100 31000 146200 31100
rect 146100 31100 146200 31200
rect 146100 31200 146200 31300
rect 146100 31300 146200 31400
rect 146100 31400 146200 31500
rect 146100 31500 146200 31600
rect 146100 31600 146200 31700
rect 146100 31700 146200 31800
rect 146100 31800 146200 31900
rect 146100 31900 146200 32000
rect 146100 32000 146200 32100
rect 146100 32100 146200 32200
rect 146100 32200 146200 32300
rect 146100 32300 146200 32400
rect 146100 32400 146200 32500
rect 146100 32500 146200 32600
rect 146100 32600 146200 32700
rect 146100 32700 146200 32800
rect 146100 32800 146200 32900
rect 146100 32900 146200 33000
rect 146100 33000 146200 33100
rect 146100 33100 146200 33200
rect 146100 33200 146200 33300
rect 146100 33300 146200 33400
rect 146100 33400 146200 33500
rect 146100 33500 146200 33600
rect 146100 33600 146200 33700
rect 146100 33700 146200 33800
rect 146100 33800 146200 33900
rect 146100 33900 146200 34000
rect 146100 34000 146200 34100
rect 146100 34100 146200 34200
rect 146100 34200 146200 34300
rect 146100 34300 146200 34400
rect 146100 34400 146200 34500
rect 146100 34500 146200 34600
rect 146100 34600 146200 34700
rect 146100 34700 146200 34800
rect 146100 34800 146200 34900
rect 146100 34900 146200 35000
rect 146100 35000 146200 35100
rect 146100 35100 146200 35200
rect 146100 35200 146200 35300
rect 146100 35300 146200 35400
rect 146200 26600 146300 26700
rect 146200 26700 146300 26800
rect 146200 26800 146300 26900
rect 146200 26900 146300 27000
rect 146200 27000 146300 27100
rect 146200 27100 146300 27200
rect 146200 27200 146300 27300
rect 146200 27300 146300 27400
rect 146200 27400 146300 27500
rect 146200 27500 146300 27600
rect 146200 27600 146300 27700
rect 146200 27700 146300 27800
rect 146200 27800 146300 27900
rect 146200 27900 146300 28000
rect 146200 28000 146300 28100
rect 146200 28100 146300 28200
rect 146200 28200 146300 28300
rect 146200 28300 146300 28400
rect 146200 28400 146300 28500
rect 146200 28500 146300 28600
rect 146200 28600 146300 28700
rect 146200 28700 146300 28800
rect 146200 28800 146300 28900
rect 146200 28900 146300 29000
rect 146200 29000 146300 29100
rect 146200 29100 146300 29200
rect 146200 29200 146300 29300
rect 146200 29300 146300 29400
rect 146200 29400 146300 29500
rect 146200 29500 146300 29600
rect 146200 29600 146300 29700
rect 146200 29700 146300 29800
rect 146200 29800 146300 29900
rect 146200 29900 146300 30000
rect 146200 30000 146300 30100
rect 146200 30100 146300 30200
rect 146200 30200 146300 30300
rect 146200 30300 146300 30400
rect 146200 30400 146300 30500
rect 146200 30500 146300 30600
rect 146200 30600 146300 30700
rect 146200 30700 146300 30800
rect 146200 30800 146300 30900
rect 146200 30900 146300 31000
rect 146200 31000 146300 31100
rect 146200 31100 146300 31200
rect 146200 31200 146300 31300
rect 146200 31300 146300 31400
rect 146200 31400 146300 31500
rect 146200 31500 146300 31600
rect 146200 31600 146300 31700
rect 146200 31700 146300 31800
rect 146200 31800 146300 31900
rect 146200 31900 146300 32000
rect 146200 32000 146300 32100
rect 146200 32100 146300 32200
rect 146200 32200 146300 32300
rect 146200 32300 146300 32400
rect 146200 32400 146300 32500
rect 146200 32500 146300 32600
rect 146200 32600 146300 32700
rect 146200 32700 146300 32800
rect 146200 32800 146300 32900
rect 146200 32900 146300 33000
rect 146200 33000 146300 33100
rect 146200 33100 146300 33200
rect 146200 33200 146300 33300
rect 146200 33300 146300 33400
rect 146200 33400 146300 33500
rect 146200 33500 146300 33600
rect 146200 33600 146300 33700
rect 146200 33700 146300 33800
rect 146200 33800 146300 33900
rect 146200 33900 146300 34000
rect 146200 34000 146300 34100
rect 146200 34100 146300 34200
rect 146200 34200 146300 34300
rect 146200 34300 146300 34400
rect 146200 34400 146300 34500
rect 146200 34500 146300 34600
rect 146200 34600 146300 34700
rect 146200 34700 146300 34800
rect 146200 34800 146300 34900
rect 146200 34900 146300 35000
rect 146200 35000 146300 35100
rect 146200 35100 146300 35200
rect 146300 26800 146400 26900
rect 146300 26900 146400 27000
rect 146300 27000 146400 27100
rect 146300 27100 146400 27200
rect 146300 27200 146400 27300
rect 146300 27300 146400 27400
rect 146300 27400 146400 27500
rect 146300 27500 146400 27600
rect 146300 27600 146400 27700
rect 146300 27700 146400 27800
rect 146300 27800 146400 27900
rect 146300 27900 146400 28000
rect 146300 28000 146400 28100
rect 146300 28100 146400 28200
rect 146300 28200 146400 28300
rect 146300 28300 146400 28400
rect 146300 28400 146400 28500
rect 146300 28500 146400 28600
rect 146300 28600 146400 28700
rect 146300 28700 146400 28800
rect 146300 28800 146400 28900
rect 146300 28900 146400 29000
rect 146300 29000 146400 29100
rect 146300 29100 146400 29200
rect 146300 29200 146400 29300
rect 146300 29300 146400 29400
rect 146300 29400 146400 29500
rect 146300 29500 146400 29600
rect 146300 29600 146400 29700
rect 146300 29700 146400 29800
rect 146300 29800 146400 29900
rect 146300 29900 146400 30000
rect 146300 30000 146400 30100
rect 146300 30100 146400 30200
rect 146300 30200 146400 30300
rect 146300 30300 146400 30400
rect 146300 30400 146400 30500
rect 146300 30500 146400 30600
rect 146300 30600 146400 30700
rect 146300 30700 146400 30800
rect 146300 30800 146400 30900
rect 146300 30900 146400 31000
rect 146300 31000 146400 31100
rect 146300 31100 146400 31200
rect 146300 31200 146400 31300
rect 146300 31300 146400 31400
rect 146300 31400 146400 31500
rect 146300 31500 146400 31600
rect 146300 31600 146400 31700
rect 146300 31700 146400 31800
rect 146300 31800 146400 31900
rect 146300 31900 146400 32000
rect 146300 32000 146400 32100
rect 146300 32100 146400 32200
rect 146300 32200 146400 32300
rect 146300 32300 146400 32400
rect 146300 32400 146400 32500
rect 146300 32500 146400 32600
rect 146300 32600 146400 32700
rect 146300 32700 146400 32800
rect 146300 32800 146400 32900
rect 146300 32900 146400 33000
rect 146300 33000 146400 33100
rect 146300 33100 146400 33200
rect 146300 33200 146400 33300
rect 146300 33300 146400 33400
rect 146300 33400 146400 33500
rect 146300 33500 146400 33600
rect 146300 33600 146400 33700
rect 146300 33700 146400 33800
rect 146300 33800 146400 33900
rect 146300 33900 146400 34000
rect 146300 34000 146400 34100
rect 146300 34100 146400 34200
rect 146300 34200 146400 34300
rect 146300 34300 146400 34400
rect 146300 34400 146400 34500
rect 146300 34500 146400 34600
rect 146300 34600 146400 34700
rect 146300 34700 146400 34800
rect 146300 34800 146400 34900
rect 146400 27100 146500 27200
rect 146400 27200 146500 27300
rect 146400 27300 146500 27400
rect 146400 27400 146500 27500
rect 146400 27500 146500 27600
rect 146400 27600 146500 27700
rect 146400 27700 146500 27800
rect 146400 27800 146500 27900
rect 146400 27900 146500 28000
rect 146400 28000 146500 28100
rect 146400 28100 146500 28200
rect 146400 28200 146500 28300
rect 146400 28300 146500 28400
rect 146400 28400 146500 28500
rect 146400 28500 146500 28600
rect 146400 28600 146500 28700
rect 146400 28700 146500 28800
rect 146400 28800 146500 28900
rect 146400 28900 146500 29000
rect 146400 29000 146500 29100
rect 146400 29100 146500 29200
rect 146400 29200 146500 29300
rect 146400 29300 146500 29400
rect 146400 29400 146500 29500
rect 146400 29500 146500 29600
rect 146400 29600 146500 29700
rect 146400 29700 146500 29800
rect 146400 29800 146500 29900
rect 146400 29900 146500 30000
rect 146400 30000 146500 30100
rect 146400 30100 146500 30200
rect 146400 30200 146500 30300
rect 146400 30300 146500 30400
rect 146400 30400 146500 30500
rect 146400 30500 146500 30600
rect 146400 30600 146500 30700
rect 146400 30700 146500 30800
rect 146400 30800 146500 30900
rect 146400 30900 146500 31000
rect 146400 31000 146500 31100
rect 146400 31100 146500 31200
rect 146400 31200 146500 31300
rect 146400 31300 146500 31400
rect 146400 31400 146500 31500
rect 146400 31500 146500 31600
rect 146400 31600 146500 31700
rect 146400 31700 146500 31800
rect 146400 31800 146500 31900
rect 146400 31900 146500 32000
rect 146400 32000 146500 32100
rect 146400 32100 146500 32200
rect 146400 32200 146500 32300
rect 146400 32300 146500 32400
rect 146400 32400 146500 32500
rect 146400 32500 146500 32600
rect 146400 32600 146500 32700
rect 146400 32700 146500 32800
rect 146400 32800 146500 32900
rect 146400 32900 146500 33000
rect 146400 33000 146500 33100
rect 146400 33100 146500 33200
rect 146400 33200 146500 33300
rect 146400 33300 146500 33400
rect 146400 33400 146500 33500
rect 146400 33500 146500 33600
rect 146400 33600 146500 33700
rect 146400 33700 146500 33800
rect 146400 33800 146500 33900
rect 146400 33900 146500 34000
rect 146400 34000 146500 34100
rect 146400 34100 146500 34200
rect 146400 34200 146500 34300
rect 146400 34300 146500 34400
rect 146400 34400 146500 34500
rect 146400 34500 146500 34600
rect 146500 27500 146600 27600
rect 146500 27600 146600 27700
rect 146500 27700 146600 27800
rect 146500 27800 146600 27900
rect 146500 27900 146600 28000
rect 146500 28000 146600 28100
rect 146500 28100 146600 28200
rect 146500 28200 146600 28300
rect 146500 28300 146600 28400
rect 146500 28400 146600 28500
rect 146500 28500 146600 28600
rect 146500 28600 146600 28700
rect 146500 28700 146600 28800
rect 146500 28800 146600 28900
rect 146500 28900 146600 29000
rect 146500 29000 146600 29100
rect 146500 29100 146600 29200
rect 146500 29200 146600 29300
rect 146500 29300 146600 29400
rect 146500 29400 146600 29500
rect 146500 29500 146600 29600
rect 146500 29600 146600 29700
rect 146500 29700 146600 29800
rect 146500 29800 146600 29900
rect 146500 29900 146600 30000
rect 146500 30000 146600 30100
rect 146500 30100 146600 30200
rect 146500 30200 146600 30300
rect 146500 30300 146600 30400
rect 146500 30400 146600 30500
rect 146500 30500 146600 30600
rect 146500 30600 146600 30700
rect 146500 30700 146600 30800
rect 146500 30800 146600 30900
rect 146500 30900 146600 31000
rect 146500 31000 146600 31100
rect 146500 31100 146600 31200
rect 146500 31200 146600 31300
rect 146500 31300 146600 31400
rect 146500 31400 146600 31500
rect 146500 31500 146600 31600
rect 146500 31600 146600 31700
rect 146500 31700 146600 31800
rect 146500 31800 146600 31900
rect 146500 31900 146600 32000
rect 146500 32000 146600 32100
rect 146500 32100 146600 32200
rect 146500 32200 146600 32300
rect 146500 32300 146600 32400
rect 146500 32400 146600 32500
rect 146500 32500 146600 32600
rect 146500 32600 146600 32700
rect 146500 32700 146600 32800
rect 146500 32800 146600 32900
rect 146500 32900 146600 33000
rect 146500 33000 146600 33100
rect 146500 33100 146600 33200
rect 146500 33200 146600 33300
rect 146500 33300 146600 33400
rect 146500 33400 146600 33500
rect 146500 33500 146600 33600
rect 146500 33600 146600 33700
rect 146500 33700 146600 33800
rect 146500 33800 146600 33900
rect 146500 33900 146600 34000
rect 146500 34000 146600 34100
rect 146500 34100 146600 34200
rect 146500 34200 146600 34300
rect 146600 27800 146700 27900
rect 146600 27900 146700 28000
rect 146600 28000 146700 28100
rect 146600 28100 146700 28200
rect 146600 28200 146700 28300
rect 146600 28300 146700 28400
rect 146600 28400 146700 28500
rect 146600 28500 146700 28600
rect 146600 28600 146700 28700
rect 146600 28700 146700 28800
rect 146600 28800 146700 28900
rect 146600 28900 146700 29000
rect 146600 29000 146700 29100
rect 146600 29100 146700 29200
rect 146600 29200 146700 29300
rect 146600 29300 146700 29400
rect 146600 29400 146700 29500
rect 146600 29500 146700 29600
rect 146600 29600 146700 29700
rect 146600 29700 146700 29800
rect 146600 29800 146700 29900
rect 146600 29900 146700 30000
rect 146600 30000 146700 30100
rect 146600 30100 146700 30200
rect 146600 30200 146700 30300
rect 146600 30300 146700 30400
rect 146600 30400 146700 30500
rect 146600 30500 146700 30600
rect 146600 30600 146700 30700
rect 146600 30700 146700 30800
rect 146600 30800 146700 30900
rect 146600 30900 146700 31000
rect 146600 31000 146700 31100
rect 146600 31100 146700 31200
rect 146600 31200 146700 31300
rect 146600 31300 146700 31400
rect 146600 31400 146700 31500
rect 146600 31500 146700 31600
rect 146600 31600 146700 31700
rect 146600 31700 146700 31800
rect 146600 31800 146700 31900
rect 146600 31900 146700 32000
rect 146600 32000 146700 32100
rect 146600 32100 146700 32200
rect 146600 32200 146700 32300
rect 146600 32300 146700 32400
rect 146600 32400 146700 32500
rect 146600 32500 146700 32600
rect 146600 32600 146700 32700
rect 146600 32700 146700 32800
rect 146600 32800 146700 32900
rect 146600 32900 146700 33000
rect 146600 33000 146700 33100
rect 146600 33100 146700 33200
rect 146600 33200 146700 33300
rect 146600 33300 146700 33400
rect 146600 33400 146700 33500
rect 146600 33500 146700 33600
rect 146600 33600 146700 33700
rect 146600 33700 146700 33800
rect 146600 33800 146700 33900
rect 146700 28300 146800 28400
rect 146700 28400 146800 28500
rect 146700 28500 146800 28600
rect 146700 28600 146800 28700
rect 146700 28700 146800 28800
rect 146700 28800 146800 28900
rect 146700 28900 146800 29000
rect 146700 29000 146800 29100
rect 146700 29100 146800 29200
rect 146700 29200 146800 29300
rect 146700 29300 146800 29400
rect 146700 29400 146800 29500
rect 146700 29500 146800 29600
rect 146700 29600 146800 29700
rect 146700 29700 146800 29800
rect 146700 29800 146800 29900
rect 146700 29900 146800 30000
rect 146700 30000 146800 30100
rect 146700 30100 146800 30200
rect 146700 30200 146800 30300
rect 146700 30300 146800 30400
rect 146700 30400 146800 30500
rect 146700 30500 146800 30600
rect 146700 30600 146800 30700
rect 146700 30700 146800 30800
rect 146700 30800 146800 30900
rect 146700 30900 146800 31000
rect 146700 31000 146800 31100
rect 146700 31100 146800 31200
rect 146700 31200 146800 31300
rect 146700 31300 146800 31400
rect 146700 31400 146800 31500
rect 146700 31500 146800 31600
rect 146700 31600 146800 31700
rect 146700 31700 146800 31800
rect 146700 31800 146800 31900
rect 146700 31900 146800 32000
rect 146700 32000 146800 32100
rect 146700 32100 146800 32200
rect 146700 32200 146800 32300
rect 146700 32300 146800 32400
rect 146700 32400 146800 32500
rect 146700 32500 146800 32600
rect 146700 32600 146800 32700
rect 146700 32700 146800 32800
rect 146700 32800 146800 32900
rect 146700 32900 146800 33000
rect 146700 33000 146800 33100
rect 146700 33100 146800 33200
rect 146700 33200 146800 33300
rect 146700 33300 146800 33400
rect 146700 33400 146800 33500
rect 146800 28800 146900 28900
rect 146800 28900 146900 29000
rect 146800 29000 146900 29100
rect 146800 29100 146900 29200
rect 146800 29200 146900 29300
rect 146800 29300 146900 29400
rect 146800 29400 146900 29500
rect 146800 29500 146900 29600
rect 146800 29600 146900 29700
rect 146800 29700 146900 29800
rect 146800 29800 146900 29900
rect 146800 29900 146900 30000
rect 146800 30000 146900 30100
rect 146800 30100 146900 30200
rect 146800 30200 146900 30300
rect 146800 30300 146900 30400
rect 146800 30400 146900 30500
rect 146800 30500 146900 30600
rect 146800 30600 146900 30700
rect 146800 30700 146900 30800
rect 146800 30800 146900 30900
rect 146800 30900 146900 31000
rect 146800 31000 146900 31100
rect 146800 31100 146900 31200
rect 146800 31200 146900 31300
rect 146800 31300 146900 31400
rect 146800 31400 146900 31500
rect 146800 31500 146900 31600
rect 146800 31600 146900 31700
rect 146800 31700 146900 31800
rect 146800 31800 146900 31900
rect 146800 31900 146900 32000
rect 146800 32000 146900 32100
rect 146800 32100 146900 32200
rect 146800 32200 146900 32300
rect 146800 32300 146900 32400
rect 146800 32400 146900 32500
rect 146800 32500 146900 32600
rect 146800 32600 146900 32700
rect 146800 32700 146900 32800
rect 146800 32800 146900 32900
rect 146900 29500 147000 29600
rect 146900 29600 147000 29700
rect 146900 29700 147000 29800
rect 146900 29800 147000 29900
rect 146900 29900 147000 30000
rect 146900 30000 147000 30100
rect 146900 30100 147000 30200
rect 146900 30200 147000 30300
rect 146900 30300 147000 30400
rect 146900 30400 147000 30500
rect 146900 30500 147000 30600
rect 146900 30600 147000 30700
rect 146900 30700 147000 30800
rect 146900 30800 147000 30900
rect 146900 30900 147000 31000
rect 146900 31000 147000 31100
rect 146900 31100 147000 31200
rect 146900 31200 147000 31300
rect 146900 31300 147000 31400
rect 146900 31400 147000 31500
rect 146900 31500 147000 31600
rect 146900 31600 147000 31700
rect 146900 31700 147000 31800
rect 146900 31800 147000 31900
rect 146900 31900 147000 32000
rect 146900 32000 147000 32100
rect 149900 29100 150000 29200
rect 149900 29200 150000 29300
rect 149900 29300 150000 29400
rect 149900 29400 150000 29500
rect 149900 29500 150000 29600
rect 149900 29600 150000 29700
rect 149900 29700 150000 29800
rect 149900 29800 150000 29900
rect 149900 29900 150000 30000
rect 149900 30000 150000 30100
rect 150000 28800 150100 28900
rect 150000 28900 150100 29000
rect 150000 29000 150100 29100
rect 150000 29100 150100 29200
rect 150000 29200 150100 29300
rect 150000 29300 150100 29400
rect 150000 29400 150100 29500
rect 150000 29500 150100 29600
rect 150000 29600 150100 29700
rect 150000 29700 150100 29800
rect 150000 29800 150100 29900
rect 150000 29900 150100 30000
rect 150000 30000 150100 30100
rect 150000 30100 150100 30200
rect 150000 30200 150100 30300
rect 150000 30300 150100 30400
rect 150100 28700 150200 28800
rect 150100 28800 150200 28900
rect 150100 28900 150200 29000
rect 150100 29000 150200 29100
rect 150100 29100 150200 29200
rect 150100 29200 150200 29300
rect 150100 29300 150200 29400
rect 150100 29400 150200 29500
rect 150100 29500 150200 29600
rect 150100 29600 150200 29700
rect 150100 29700 150200 29800
rect 150100 29800 150200 29900
rect 150100 29900 150200 30000
rect 150100 30000 150200 30100
rect 150100 30100 150200 30200
rect 150100 30200 150200 30300
rect 150100 30300 150200 30400
rect 150100 30400 150200 30500
rect 150100 30500 150200 30600
rect 150100 30600 150200 30700
rect 150200 22200 150300 22300
rect 150200 22300 150300 22400
rect 150200 22400 150300 22500
rect 150200 22500 150300 22600
rect 150200 22600 150300 22700
rect 150200 22700 150300 22800
rect 150200 22800 150300 22900
rect 150200 22900 150300 23000
rect 150200 23000 150300 23100
rect 150200 23100 150300 23200
rect 150200 23200 150300 23300
rect 150200 23300 150300 23400
rect 150200 23400 150300 23500
rect 150200 23500 150300 23600
rect 150200 23600 150300 23700
rect 150200 23700 150300 23800
rect 150200 23800 150300 23900
rect 150200 23900 150300 24000
rect 150200 24000 150300 24100
rect 150200 24100 150300 24200
rect 150200 24200 150300 24300
rect 150200 24300 150300 24400
rect 150200 24400 150300 24500
rect 150200 24500 150300 24600
rect 150200 24600 150300 24700
rect 150200 24700 150300 24800
rect 150200 24800 150300 24900
rect 150200 24900 150300 25000
rect 150200 25000 150300 25100
rect 150200 25100 150300 25200
rect 150200 25200 150300 25300
rect 150200 25300 150300 25400
rect 150200 25400 150300 25500
rect 150200 25500 150300 25600
rect 150200 25600 150300 25700
rect 150200 25800 150300 25900
rect 150200 26000 150300 26100
rect 150200 28500 150300 28600
rect 150200 28600 150300 28700
rect 150200 28700 150300 28800
rect 150200 28800 150300 28900
rect 150200 28900 150300 29000
rect 150200 29000 150300 29100
rect 150200 29100 150300 29200
rect 150200 29200 150300 29300
rect 150200 29300 150300 29400
rect 150200 29400 150300 29500
rect 150200 29500 150300 29600
rect 150200 29600 150300 29700
rect 150200 29700 150300 29800
rect 150200 29800 150300 29900
rect 150200 29900 150300 30000
rect 150200 30000 150300 30100
rect 150200 30100 150300 30200
rect 150200 30200 150300 30300
rect 150200 30300 150300 30400
rect 150200 30400 150300 30500
rect 150200 30500 150300 30600
rect 150200 30600 150300 30700
rect 150200 30700 150300 30800
rect 150200 30800 150300 30900
rect 150300 21900 150400 22000
rect 150300 22000 150400 22100
rect 150300 22100 150400 22200
rect 150300 22200 150400 22300
rect 150300 22300 150400 22400
rect 150300 22400 150400 22500
rect 150300 22500 150400 22600
rect 150300 22600 150400 22700
rect 150300 22700 150400 22800
rect 150300 22800 150400 22900
rect 150300 22900 150400 23000
rect 150300 23000 150400 23100
rect 150300 23100 150400 23200
rect 150300 23200 150400 23300
rect 150300 23300 150400 23400
rect 150300 23400 150400 23500
rect 150300 23500 150400 23600
rect 150300 23600 150400 23700
rect 150300 23700 150400 23800
rect 150300 23800 150400 23900
rect 150300 23900 150400 24000
rect 150300 24000 150400 24100
rect 150300 24100 150400 24200
rect 150300 24200 150400 24300
rect 150300 24300 150400 24400
rect 150300 24400 150400 24500
rect 150300 24500 150400 24600
rect 150300 24600 150400 24700
rect 150300 24700 150400 24800
rect 150300 24800 150400 24900
rect 150300 24900 150400 25000
rect 150300 25000 150400 25100
rect 150300 25100 150400 25200
rect 150300 25200 150400 25300
rect 150300 25300 150400 25400
rect 150300 25400 150400 25500
rect 150300 25500 150400 25600
rect 150300 25600 150400 25700
rect 150300 25700 150400 25800
rect 150300 25800 150400 25900
rect 150300 25900 150400 26000
rect 150300 26000 150400 26100
rect 150300 26100 150400 26200
rect 150300 26200 150400 26300
rect 150300 26300 150400 26400
rect 150300 26400 150400 26500
rect 150300 26500 150400 26600
rect 150300 26600 150400 26700
rect 150300 26700 150400 26800
rect 150300 26800 150400 26900
rect 150300 26900 150400 27000
rect 150300 27000 150400 27100
rect 150300 27100 150400 27200
rect 150300 27200 150400 27300
rect 150300 27300 150400 27400
rect 150300 27400 150400 27500
rect 150300 27500 150400 27600
rect 150300 27600 150400 27700
rect 150300 27700 150400 27800
rect 150300 27800 150400 27900
rect 150300 27900 150400 28000
rect 150300 28000 150400 28100
rect 150300 28100 150400 28200
rect 150300 28200 150400 28300
rect 150300 28300 150400 28400
rect 150300 28400 150400 28500
rect 150300 28500 150400 28600
rect 150300 28600 150400 28700
rect 150300 28700 150400 28800
rect 150300 28800 150400 28900
rect 150300 28900 150400 29000
rect 150300 29000 150400 29100
rect 150300 29100 150400 29200
rect 150300 29200 150400 29300
rect 150300 29300 150400 29400
rect 150300 29400 150400 29500
rect 150300 29500 150400 29600
rect 150300 29600 150400 29700
rect 150300 29700 150400 29800
rect 150300 29800 150400 29900
rect 150300 29900 150400 30000
rect 150300 30000 150400 30100
rect 150300 30100 150400 30200
rect 150300 30200 150400 30300
rect 150300 30300 150400 30400
rect 150300 30400 150400 30500
rect 150300 30500 150400 30600
rect 150300 30600 150400 30700
rect 150300 30700 150400 30800
rect 150300 30800 150400 30900
rect 150300 30900 150400 31000
rect 150300 31000 150400 31100
rect 150400 21700 150500 21800
rect 150400 21800 150500 21900
rect 150400 21900 150500 22000
rect 150400 22000 150500 22100
rect 150400 22100 150500 22200
rect 150400 22200 150500 22300
rect 150400 22300 150500 22400
rect 150400 22400 150500 22500
rect 150400 22500 150500 22600
rect 150400 22600 150500 22700
rect 150400 22700 150500 22800
rect 150400 22800 150500 22900
rect 150400 22900 150500 23000
rect 150400 23000 150500 23100
rect 150400 23100 150500 23200
rect 150400 23200 150500 23300
rect 150400 23300 150500 23400
rect 150400 23400 150500 23500
rect 150400 23500 150500 23600
rect 150400 23600 150500 23700
rect 150400 23700 150500 23800
rect 150400 23800 150500 23900
rect 150400 23900 150500 24000
rect 150400 24000 150500 24100
rect 150400 24100 150500 24200
rect 150400 24200 150500 24300
rect 150400 24300 150500 24400
rect 150400 24400 150500 24500
rect 150400 24500 150500 24600
rect 150400 24600 150500 24700
rect 150400 24700 150500 24800
rect 150400 24800 150500 24900
rect 150400 24900 150500 25000
rect 150400 25000 150500 25100
rect 150400 25100 150500 25200
rect 150400 25200 150500 25300
rect 150400 25300 150500 25400
rect 150400 25400 150500 25500
rect 150400 25500 150500 25600
rect 150400 25600 150500 25700
rect 150400 25700 150500 25800
rect 150400 25800 150500 25900
rect 150400 25900 150500 26000
rect 150400 26000 150500 26100
rect 150400 26100 150500 26200
rect 150400 26200 150500 26300
rect 150400 26300 150500 26400
rect 150400 26400 150500 26500
rect 150400 26500 150500 26600
rect 150400 26600 150500 26700
rect 150400 26700 150500 26800
rect 150400 26800 150500 26900
rect 150400 26900 150500 27000
rect 150400 27000 150500 27100
rect 150400 27100 150500 27200
rect 150400 27200 150500 27300
rect 150400 27300 150500 27400
rect 150400 27400 150500 27500
rect 150400 27500 150500 27600
rect 150400 27600 150500 27700
rect 150400 27700 150500 27800
rect 150400 27800 150500 27900
rect 150400 27900 150500 28000
rect 150400 28000 150500 28100
rect 150400 28100 150500 28200
rect 150400 28200 150500 28300
rect 150400 28300 150500 28400
rect 150400 28400 150500 28500
rect 150400 28500 150500 28600
rect 150400 28600 150500 28700
rect 150400 28700 150500 28800
rect 150400 28800 150500 28900
rect 150400 28900 150500 29000
rect 150400 29000 150500 29100
rect 150400 29100 150500 29200
rect 150400 29200 150500 29300
rect 150400 29300 150500 29400
rect 150400 29400 150500 29500
rect 150400 29500 150500 29600
rect 150400 29600 150500 29700
rect 150400 29700 150500 29800
rect 150400 29800 150500 29900
rect 150400 29900 150500 30000
rect 150400 30000 150500 30100
rect 150400 30100 150500 30200
rect 150400 30200 150500 30300
rect 150400 30300 150500 30400
rect 150400 30400 150500 30500
rect 150400 30500 150500 30600
rect 150400 30600 150500 30700
rect 150400 30700 150500 30800
rect 150400 30800 150500 30900
rect 150400 30900 150500 31000
rect 150400 31000 150500 31100
rect 150400 31100 150500 31200
rect 150400 31200 150500 31300
rect 150400 31300 150500 31400
rect 150400 31400 150500 31500
rect 150400 31500 150500 31600
rect 150400 31600 150500 31700
rect 150400 31700 150500 31800
rect 150400 31800 150500 31900
rect 150400 31900 150500 32000
rect 150400 32000 150500 32100
rect 150400 32100 150500 32200
rect 150400 32200 150500 32300
rect 150400 32300 150500 32400
rect 150400 32400 150500 32500
rect 150400 32500 150500 32600
rect 150400 32600 150500 32700
rect 150400 32700 150500 32800
rect 150400 32800 150500 32900
rect 150400 32900 150500 33000
rect 150400 33000 150500 33100
rect 150400 33100 150500 33200
rect 150400 33200 150500 33300
rect 150400 33300 150500 33400
rect 150400 33400 150500 33500
rect 150400 33500 150500 33600
rect 150400 33600 150500 33700
rect 150400 33700 150500 33800
rect 150400 33800 150500 33900
rect 150400 34000 150500 34100
rect 150400 34200 150500 34300
rect 150500 21600 150600 21700
rect 150500 21700 150600 21800
rect 150500 21800 150600 21900
rect 150500 21900 150600 22000
rect 150500 22000 150600 22100
rect 150500 22100 150600 22200
rect 150500 22200 150600 22300
rect 150500 22300 150600 22400
rect 150500 22400 150600 22500
rect 150500 22500 150600 22600
rect 150500 22600 150600 22700
rect 150500 22700 150600 22800
rect 150500 22800 150600 22900
rect 150500 22900 150600 23000
rect 150500 23000 150600 23100
rect 150500 23100 150600 23200
rect 150500 23200 150600 23300
rect 150500 23300 150600 23400
rect 150500 23400 150600 23500
rect 150500 23500 150600 23600
rect 150500 23600 150600 23700
rect 150500 23700 150600 23800
rect 150500 23800 150600 23900
rect 150500 23900 150600 24000
rect 150500 24000 150600 24100
rect 150500 24100 150600 24200
rect 150500 24200 150600 24300
rect 150500 24300 150600 24400
rect 150500 24400 150600 24500
rect 150500 24500 150600 24600
rect 150500 24600 150600 24700
rect 150500 24700 150600 24800
rect 150500 24800 150600 24900
rect 150500 24900 150600 25000
rect 150500 25000 150600 25100
rect 150500 25100 150600 25200
rect 150500 25200 150600 25300
rect 150500 25300 150600 25400
rect 150500 25400 150600 25500
rect 150500 25500 150600 25600
rect 150500 25600 150600 25700
rect 150500 25700 150600 25800
rect 150500 25800 150600 25900
rect 150500 25900 150600 26000
rect 150500 26000 150600 26100
rect 150500 26100 150600 26200
rect 150500 26200 150600 26300
rect 150500 26300 150600 26400
rect 150500 26400 150600 26500
rect 150500 26500 150600 26600
rect 150500 26600 150600 26700
rect 150500 26700 150600 26800
rect 150500 26800 150600 26900
rect 150500 26900 150600 27000
rect 150500 27000 150600 27100
rect 150500 27100 150600 27200
rect 150500 27200 150600 27300
rect 150500 27300 150600 27400
rect 150500 27400 150600 27500
rect 150500 27500 150600 27600
rect 150500 27600 150600 27700
rect 150500 27700 150600 27800
rect 150500 27800 150600 27900
rect 150500 27900 150600 28000
rect 150500 28000 150600 28100
rect 150500 28100 150600 28200
rect 150500 28200 150600 28300
rect 150500 28300 150600 28400
rect 150500 28400 150600 28500
rect 150500 28500 150600 28600
rect 150500 28600 150600 28700
rect 150500 28700 150600 28800
rect 150500 28800 150600 28900
rect 150500 28900 150600 29000
rect 150500 29000 150600 29100
rect 150500 29100 150600 29200
rect 150500 29200 150600 29300
rect 150500 29300 150600 29400
rect 150500 29400 150600 29500
rect 150500 29500 150600 29600
rect 150500 29600 150600 29700
rect 150500 29700 150600 29800
rect 150500 29800 150600 29900
rect 150500 29900 150600 30000
rect 150500 30000 150600 30100
rect 150500 30100 150600 30200
rect 150500 30200 150600 30300
rect 150500 30300 150600 30400
rect 150500 30400 150600 30500
rect 150500 30500 150600 30600
rect 150500 30600 150600 30700
rect 150500 30700 150600 30800
rect 150500 30800 150600 30900
rect 150500 30900 150600 31000
rect 150500 31000 150600 31100
rect 150500 31100 150600 31200
rect 150500 31200 150600 31300
rect 150500 31300 150600 31400
rect 150500 31400 150600 31500
rect 150500 31500 150600 31600
rect 150500 31600 150600 31700
rect 150500 31700 150600 31800
rect 150500 31800 150600 31900
rect 150500 31900 150600 32000
rect 150500 32000 150600 32100
rect 150500 32100 150600 32200
rect 150500 32200 150600 32300
rect 150500 32300 150600 32400
rect 150500 32400 150600 32500
rect 150500 32500 150600 32600
rect 150500 32600 150600 32700
rect 150500 32700 150600 32800
rect 150500 32800 150600 32900
rect 150500 32900 150600 33000
rect 150500 33000 150600 33100
rect 150500 33100 150600 33200
rect 150500 33200 150600 33300
rect 150500 33300 150600 33400
rect 150500 33400 150600 33500
rect 150500 33500 150600 33600
rect 150500 33600 150600 33700
rect 150500 33700 150600 33800
rect 150500 33800 150600 33900
rect 150500 33900 150600 34000
rect 150500 34000 150600 34100
rect 150500 34100 150600 34200
rect 150500 34200 150600 34300
rect 150500 34300 150600 34400
rect 150500 34400 150600 34500
rect 150500 34500 150600 34600
rect 150500 34600 150600 34700
rect 150500 34700 150600 34800
rect 150500 34800 150600 34900
rect 150500 34900 150600 35000
rect 150500 35000 150600 35100
rect 150500 35100 150600 35200
rect 150500 35200 150600 35300
rect 150500 35300 150600 35400
rect 150500 35400 150600 35500
rect 150500 35500 150600 35600
rect 150500 35600 150600 35700
rect 150500 35700 150600 35800
rect 150500 35800 150600 35900
rect 150500 35900 150600 36000
rect 150500 36000 150600 36100
rect 150500 36100 150600 36200
rect 150500 36200 150600 36300
rect 150500 36300 150600 36400
rect 150500 36400 150600 36500
rect 150500 36500 150600 36600
rect 150500 36600 150600 36700
rect 150500 36700 150600 36800
rect 150500 36800 150600 36900
rect 150500 36900 150600 37000
rect 150500 37000 150600 37100
rect 150500 37100 150600 37200
rect 150500 37200 150600 37300
rect 150500 37300 150600 37400
rect 150500 37400 150600 37500
rect 150500 37500 150600 37600
rect 150600 21500 150700 21600
rect 150600 21600 150700 21700
rect 150600 21700 150700 21800
rect 150600 21800 150700 21900
rect 150600 21900 150700 22000
rect 150600 22000 150700 22100
rect 150600 22100 150700 22200
rect 150600 22200 150700 22300
rect 150600 22300 150700 22400
rect 150600 22400 150700 22500
rect 150600 22500 150700 22600
rect 150600 22600 150700 22700
rect 150600 22700 150700 22800
rect 150600 22800 150700 22900
rect 150600 22900 150700 23000
rect 150600 23000 150700 23100
rect 150600 23100 150700 23200
rect 150600 23200 150700 23300
rect 150600 23300 150700 23400
rect 150600 23400 150700 23500
rect 150600 23500 150700 23600
rect 150600 23600 150700 23700
rect 150600 23700 150700 23800
rect 150600 23800 150700 23900
rect 150600 23900 150700 24000
rect 150600 24000 150700 24100
rect 150600 24100 150700 24200
rect 150600 24200 150700 24300
rect 150600 24300 150700 24400
rect 150600 24400 150700 24500
rect 150600 24500 150700 24600
rect 150600 24600 150700 24700
rect 150600 24700 150700 24800
rect 150600 24800 150700 24900
rect 150600 24900 150700 25000
rect 150600 25000 150700 25100
rect 150600 25100 150700 25200
rect 150600 25200 150700 25300
rect 150600 25300 150700 25400
rect 150600 25400 150700 25500
rect 150600 25500 150700 25600
rect 150600 25600 150700 25700
rect 150600 25700 150700 25800
rect 150600 25800 150700 25900
rect 150600 25900 150700 26000
rect 150600 26000 150700 26100
rect 150600 26100 150700 26200
rect 150600 26200 150700 26300
rect 150600 26300 150700 26400
rect 150600 26400 150700 26500
rect 150600 26500 150700 26600
rect 150600 26600 150700 26700
rect 150600 26700 150700 26800
rect 150600 26800 150700 26900
rect 150600 26900 150700 27000
rect 150600 27000 150700 27100
rect 150600 27100 150700 27200
rect 150600 27200 150700 27300
rect 150600 27300 150700 27400
rect 150600 27400 150700 27500
rect 150600 27500 150700 27600
rect 150600 27600 150700 27700
rect 150600 27700 150700 27800
rect 150600 27800 150700 27900
rect 150600 27900 150700 28000
rect 150600 28000 150700 28100
rect 150600 28100 150700 28200
rect 150600 28200 150700 28300
rect 150600 28300 150700 28400
rect 150600 28400 150700 28500
rect 150600 28500 150700 28600
rect 150600 28600 150700 28700
rect 150600 28700 150700 28800
rect 150600 28800 150700 28900
rect 150600 28900 150700 29000
rect 150600 29000 150700 29100
rect 150600 29100 150700 29200
rect 150600 29200 150700 29300
rect 150600 29300 150700 29400
rect 150600 29400 150700 29500
rect 150600 29500 150700 29600
rect 150600 29600 150700 29700
rect 150600 29700 150700 29800
rect 150600 29800 150700 29900
rect 150600 29900 150700 30000
rect 150600 30000 150700 30100
rect 150600 30100 150700 30200
rect 150600 30200 150700 30300
rect 150600 30300 150700 30400
rect 150600 30400 150700 30500
rect 150600 30500 150700 30600
rect 150600 30600 150700 30700
rect 150600 30700 150700 30800
rect 150600 30800 150700 30900
rect 150600 30900 150700 31000
rect 150600 31000 150700 31100
rect 150600 31100 150700 31200
rect 150600 31200 150700 31300
rect 150600 31300 150700 31400
rect 150600 31400 150700 31500
rect 150600 31500 150700 31600
rect 150600 31600 150700 31700
rect 150600 31700 150700 31800
rect 150600 31800 150700 31900
rect 150600 31900 150700 32000
rect 150600 32000 150700 32100
rect 150600 32100 150700 32200
rect 150600 32200 150700 32300
rect 150600 32300 150700 32400
rect 150600 32400 150700 32500
rect 150600 32500 150700 32600
rect 150600 32600 150700 32700
rect 150600 32700 150700 32800
rect 150600 32800 150700 32900
rect 150600 32900 150700 33000
rect 150600 33000 150700 33100
rect 150600 33100 150700 33200
rect 150600 33200 150700 33300
rect 150600 33300 150700 33400
rect 150600 33400 150700 33500
rect 150600 33500 150700 33600
rect 150600 33600 150700 33700
rect 150600 33700 150700 33800
rect 150600 33800 150700 33900
rect 150600 33900 150700 34000
rect 150600 34000 150700 34100
rect 150600 34100 150700 34200
rect 150600 34200 150700 34300
rect 150600 34300 150700 34400
rect 150600 34400 150700 34500
rect 150600 34500 150700 34600
rect 150600 34600 150700 34700
rect 150600 34700 150700 34800
rect 150600 34800 150700 34900
rect 150600 34900 150700 35000
rect 150600 35000 150700 35100
rect 150600 35100 150700 35200
rect 150600 35200 150700 35300
rect 150600 35300 150700 35400
rect 150600 35400 150700 35500
rect 150600 35500 150700 35600
rect 150600 35600 150700 35700
rect 150600 35700 150700 35800
rect 150600 35800 150700 35900
rect 150600 35900 150700 36000
rect 150600 36000 150700 36100
rect 150600 36100 150700 36200
rect 150600 36200 150700 36300
rect 150600 36300 150700 36400
rect 150600 36400 150700 36500
rect 150600 36500 150700 36600
rect 150600 36600 150700 36700
rect 150600 36700 150700 36800
rect 150600 36800 150700 36900
rect 150600 36900 150700 37000
rect 150600 37000 150700 37100
rect 150600 37100 150700 37200
rect 150600 37200 150700 37300
rect 150600 37300 150700 37400
rect 150600 37400 150700 37500
rect 150600 37500 150700 37600
rect 150600 37600 150700 37700
rect 150600 37700 150700 37800
rect 150600 37800 150700 37900
rect 150700 21400 150800 21500
rect 150700 21500 150800 21600
rect 150700 21600 150800 21700
rect 150700 21700 150800 21800
rect 150700 21800 150800 21900
rect 150700 21900 150800 22000
rect 150700 22000 150800 22100
rect 150700 22100 150800 22200
rect 150700 22200 150800 22300
rect 150700 22300 150800 22400
rect 150700 22400 150800 22500
rect 150700 22500 150800 22600
rect 150700 22600 150800 22700
rect 150700 22700 150800 22800
rect 150700 22800 150800 22900
rect 150700 22900 150800 23000
rect 150700 23000 150800 23100
rect 150700 23100 150800 23200
rect 150700 23200 150800 23300
rect 150700 23300 150800 23400
rect 150700 23400 150800 23500
rect 150700 23500 150800 23600
rect 150700 23600 150800 23700
rect 150700 23700 150800 23800
rect 150700 23800 150800 23900
rect 150700 23900 150800 24000
rect 150700 24000 150800 24100
rect 150700 24100 150800 24200
rect 150700 24200 150800 24300
rect 150700 24300 150800 24400
rect 150700 24400 150800 24500
rect 150700 24500 150800 24600
rect 150700 24600 150800 24700
rect 150700 24700 150800 24800
rect 150700 24800 150800 24900
rect 150700 24900 150800 25000
rect 150700 25000 150800 25100
rect 150700 25100 150800 25200
rect 150700 25200 150800 25300
rect 150700 25300 150800 25400
rect 150700 25400 150800 25500
rect 150700 25500 150800 25600
rect 150700 25600 150800 25700
rect 150700 25700 150800 25800
rect 150700 25800 150800 25900
rect 150700 25900 150800 26000
rect 150700 26000 150800 26100
rect 150700 26100 150800 26200
rect 150700 26200 150800 26300
rect 150700 26300 150800 26400
rect 150700 26400 150800 26500
rect 150700 26500 150800 26600
rect 150700 26600 150800 26700
rect 150700 26700 150800 26800
rect 150700 26800 150800 26900
rect 150700 26900 150800 27000
rect 150700 27000 150800 27100
rect 150700 27100 150800 27200
rect 150700 27200 150800 27300
rect 150700 27300 150800 27400
rect 150700 27400 150800 27500
rect 150700 27500 150800 27600
rect 150700 27600 150800 27700
rect 150700 27700 150800 27800
rect 150700 27800 150800 27900
rect 150700 27900 150800 28000
rect 150700 28000 150800 28100
rect 150700 28100 150800 28200
rect 150700 28200 150800 28300
rect 150700 28300 150800 28400
rect 150700 28400 150800 28500
rect 150700 28500 150800 28600
rect 150700 28600 150800 28700
rect 150700 28700 150800 28800
rect 150700 28800 150800 28900
rect 150700 28900 150800 29000
rect 150700 29000 150800 29100
rect 150700 29100 150800 29200
rect 150700 29200 150800 29300
rect 150700 29300 150800 29400
rect 150700 29400 150800 29500
rect 150700 29500 150800 29600
rect 150700 29600 150800 29700
rect 150700 29700 150800 29800
rect 150700 29800 150800 29900
rect 150700 29900 150800 30000
rect 150700 30000 150800 30100
rect 150700 30100 150800 30200
rect 150700 30200 150800 30300
rect 150700 30300 150800 30400
rect 150700 30400 150800 30500
rect 150700 30500 150800 30600
rect 150700 30600 150800 30700
rect 150700 30700 150800 30800
rect 150700 30800 150800 30900
rect 150700 30900 150800 31000
rect 150700 31000 150800 31100
rect 150700 31100 150800 31200
rect 150700 31200 150800 31300
rect 150700 31300 150800 31400
rect 150700 31400 150800 31500
rect 150700 31500 150800 31600
rect 150700 31600 150800 31700
rect 150700 31700 150800 31800
rect 150700 31800 150800 31900
rect 150700 31900 150800 32000
rect 150700 32000 150800 32100
rect 150700 32100 150800 32200
rect 150700 32200 150800 32300
rect 150700 32300 150800 32400
rect 150700 32400 150800 32500
rect 150700 32500 150800 32600
rect 150700 32600 150800 32700
rect 150700 32700 150800 32800
rect 150700 32800 150800 32900
rect 150700 32900 150800 33000
rect 150700 33000 150800 33100
rect 150700 33100 150800 33200
rect 150700 33200 150800 33300
rect 150700 33300 150800 33400
rect 150700 33400 150800 33500
rect 150700 33500 150800 33600
rect 150700 33600 150800 33700
rect 150700 33700 150800 33800
rect 150700 33800 150800 33900
rect 150700 33900 150800 34000
rect 150700 34000 150800 34100
rect 150700 34100 150800 34200
rect 150700 34200 150800 34300
rect 150700 34300 150800 34400
rect 150700 34400 150800 34500
rect 150700 34500 150800 34600
rect 150700 34600 150800 34700
rect 150700 34700 150800 34800
rect 150700 34800 150800 34900
rect 150700 34900 150800 35000
rect 150700 35000 150800 35100
rect 150700 35100 150800 35200
rect 150700 35200 150800 35300
rect 150700 35300 150800 35400
rect 150700 35400 150800 35500
rect 150700 35500 150800 35600
rect 150700 35600 150800 35700
rect 150700 35700 150800 35800
rect 150700 35800 150800 35900
rect 150700 35900 150800 36000
rect 150700 36000 150800 36100
rect 150700 36100 150800 36200
rect 150700 36200 150800 36300
rect 150700 36300 150800 36400
rect 150700 36400 150800 36500
rect 150700 36500 150800 36600
rect 150700 36600 150800 36700
rect 150700 36700 150800 36800
rect 150700 36800 150800 36900
rect 150700 36900 150800 37000
rect 150700 37000 150800 37100
rect 150700 37100 150800 37200
rect 150700 37200 150800 37300
rect 150700 37300 150800 37400
rect 150700 37400 150800 37500
rect 150700 37500 150800 37600
rect 150700 37600 150800 37700
rect 150700 37700 150800 37800
rect 150700 37800 150800 37900
rect 150700 37900 150800 38000
rect 150800 21300 150900 21400
rect 150800 21400 150900 21500
rect 150800 21500 150900 21600
rect 150800 21600 150900 21700
rect 150800 21700 150900 21800
rect 150800 21800 150900 21900
rect 150800 21900 150900 22000
rect 150800 22000 150900 22100
rect 150800 22100 150900 22200
rect 150800 22200 150900 22300
rect 150800 22300 150900 22400
rect 150800 22400 150900 22500
rect 150800 22500 150900 22600
rect 150800 22600 150900 22700
rect 150800 22700 150900 22800
rect 150800 22800 150900 22900
rect 150800 22900 150900 23000
rect 150800 23000 150900 23100
rect 150800 23100 150900 23200
rect 150800 23200 150900 23300
rect 150800 23300 150900 23400
rect 150800 23400 150900 23500
rect 150800 23500 150900 23600
rect 150800 23600 150900 23700
rect 150800 23700 150900 23800
rect 150800 23800 150900 23900
rect 150800 23900 150900 24000
rect 150800 24000 150900 24100
rect 150800 24100 150900 24200
rect 150800 24200 150900 24300
rect 150800 24300 150900 24400
rect 150800 24400 150900 24500
rect 150800 24500 150900 24600
rect 150800 24600 150900 24700
rect 150800 24700 150900 24800
rect 150800 24800 150900 24900
rect 150800 24900 150900 25000
rect 150800 25000 150900 25100
rect 150800 25100 150900 25200
rect 150800 25200 150900 25300
rect 150800 25300 150900 25400
rect 150800 25400 150900 25500
rect 150800 25500 150900 25600
rect 150800 25600 150900 25700
rect 150800 25700 150900 25800
rect 150800 25800 150900 25900
rect 150800 25900 150900 26000
rect 150800 26000 150900 26100
rect 150800 26100 150900 26200
rect 150800 26200 150900 26300
rect 150800 26300 150900 26400
rect 150800 26400 150900 26500
rect 150800 26500 150900 26600
rect 150800 26600 150900 26700
rect 150800 26700 150900 26800
rect 150800 26800 150900 26900
rect 150800 26900 150900 27000
rect 150800 27000 150900 27100
rect 150800 27100 150900 27200
rect 150800 27200 150900 27300
rect 150800 27300 150900 27400
rect 150800 27400 150900 27500
rect 150800 27500 150900 27600
rect 150800 27600 150900 27700
rect 150800 27700 150900 27800
rect 150800 27800 150900 27900
rect 150800 27900 150900 28000
rect 150800 28000 150900 28100
rect 150800 28100 150900 28200
rect 150800 28200 150900 28300
rect 150800 28300 150900 28400
rect 150800 28400 150900 28500
rect 150800 28500 150900 28600
rect 150800 28600 150900 28700
rect 150800 28700 150900 28800
rect 150800 28800 150900 28900
rect 150800 28900 150900 29000
rect 150800 29000 150900 29100
rect 150800 29100 150900 29200
rect 150800 29200 150900 29300
rect 150800 29300 150900 29400
rect 150800 29400 150900 29500
rect 150800 29500 150900 29600
rect 150800 29600 150900 29700
rect 150800 29700 150900 29800
rect 150800 29800 150900 29900
rect 150800 29900 150900 30000
rect 150800 30000 150900 30100
rect 150800 30100 150900 30200
rect 150800 30200 150900 30300
rect 150800 30300 150900 30400
rect 150800 30400 150900 30500
rect 150800 30500 150900 30600
rect 150800 30600 150900 30700
rect 150800 30700 150900 30800
rect 150800 30800 150900 30900
rect 150800 30900 150900 31000
rect 150800 31000 150900 31100
rect 150800 31100 150900 31200
rect 150800 31200 150900 31300
rect 150800 31300 150900 31400
rect 150800 31400 150900 31500
rect 150800 31500 150900 31600
rect 150800 31600 150900 31700
rect 150800 31700 150900 31800
rect 150800 31800 150900 31900
rect 150800 31900 150900 32000
rect 150800 32000 150900 32100
rect 150800 32100 150900 32200
rect 150800 32200 150900 32300
rect 150800 32300 150900 32400
rect 150800 32400 150900 32500
rect 150800 32500 150900 32600
rect 150800 32600 150900 32700
rect 150800 32700 150900 32800
rect 150800 32800 150900 32900
rect 150800 32900 150900 33000
rect 150800 33000 150900 33100
rect 150800 33100 150900 33200
rect 150800 33200 150900 33300
rect 150800 33300 150900 33400
rect 150800 33400 150900 33500
rect 150800 33500 150900 33600
rect 150800 33600 150900 33700
rect 150800 33700 150900 33800
rect 150800 33800 150900 33900
rect 150800 33900 150900 34000
rect 150800 34000 150900 34100
rect 150800 34100 150900 34200
rect 150800 34200 150900 34300
rect 150800 34300 150900 34400
rect 150800 34400 150900 34500
rect 150800 34500 150900 34600
rect 150800 34600 150900 34700
rect 150800 34700 150900 34800
rect 150800 34800 150900 34900
rect 150800 34900 150900 35000
rect 150800 35000 150900 35100
rect 150800 35100 150900 35200
rect 150800 35200 150900 35300
rect 150800 35300 150900 35400
rect 150800 35400 150900 35500
rect 150800 35500 150900 35600
rect 150800 35600 150900 35700
rect 150800 35700 150900 35800
rect 150800 35800 150900 35900
rect 150800 35900 150900 36000
rect 150800 36000 150900 36100
rect 150800 36100 150900 36200
rect 150800 36200 150900 36300
rect 150800 36300 150900 36400
rect 150800 36400 150900 36500
rect 150800 36500 150900 36600
rect 150800 36600 150900 36700
rect 150800 36700 150900 36800
rect 150800 36800 150900 36900
rect 150800 36900 150900 37000
rect 150800 37000 150900 37100
rect 150800 37100 150900 37200
rect 150800 37200 150900 37300
rect 150800 37300 150900 37400
rect 150800 37400 150900 37500
rect 150800 37500 150900 37600
rect 150800 37600 150900 37700
rect 150800 37700 150900 37800
rect 150800 37800 150900 37900
rect 150800 37900 150900 38000
rect 150800 38000 150900 38100
rect 150900 21200 151000 21300
rect 150900 21300 151000 21400
rect 150900 21400 151000 21500
rect 150900 21500 151000 21600
rect 150900 21600 151000 21700
rect 150900 21700 151000 21800
rect 150900 21800 151000 21900
rect 150900 21900 151000 22000
rect 150900 22000 151000 22100
rect 150900 22100 151000 22200
rect 150900 22200 151000 22300
rect 150900 22300 151000 22400
rect 150900 22400 151000 22500
rect 150900 22500 151000 22600
rect 150900 22600 151000 22700
rect 150900 22700 151000 22800
rect 150900 22800 151000 22900
rect 150900 22900 151000 23000
rect 150900 23000 151000 23100
rect 150900 23100 151000 23200
rect 150900 23200 151000 23300
rect 150900 23300 151000 23400
rect 150900 23400 151000 23500
rect 150900 23500 151000 23600
rect 150900 23600 151000 23700
rect 150900 23700 151000 23800
rect 150900 23800 151000 23900
rect 150900 23900 151000 24000
rect 150900 24000 151000 24100
rect 150900 24100 151000 24200
rect 150900 24200 151000 24300
rect 150900 24300 151000 24400
rect 150900 24400 151000 24500
rect 150900 24500 151000 24600
rect 150900 24600 151000 24700
rect 150900 24700 151000 24800
rect 150900 24800 151000 24900
rect 150900 24900 151000 25000
rect 150900 25000 151000 25100
rect 150900 25100 151000 25200
rect 150900 25200 151000 25300
rect 150900 25300 151000 25400
rect 150900 25400 151000 25500
rect 150900 25500 151000 25600
rect 150900 25600 151000 25700
rect 150900 25700 151000 25800
rect 150900 25800 151000 25900
rect 150900 25900 151000 26000
rect 150900 26000 151000 26100
rect 150900 26100 151000 26200
rect 150900 26200 151000 26300
rect 150900 26300 151000 26400
rect 150900 26400 151000 26500
rect 150900 26500 151000 26600
rect 150900 26600 151000 26700
rect 150900 26700 151000 26800
rect 150900 26800 151000 26900
rect 150900 26900 151000 27000
rect 150900 27000 151000 27100
rect 150900 27100 151000 27200
rect 150900 27200 151000 27300
rect 150900 27300 151000 27400
rect 150900 27400 151000 27500
rect 150900 27500 151000 27600
rect 150900 27600 151000 27700
rect 150900 27700 151000 27800
rect 150900 27800 151000 27900
rect 150900 27900 151000 28000
rect 150900 28000 151000 28100
rect 150900 28100 151000 28200
rect 150900 28200 151000 28300
rect 150900 28300 151000 28400
rect 150900 28400 151000 28500
rect 150900 28500 151000 28600
rect 150900 28600 151000 28700
rect 150900 28700 151000 28800
rect 150900 28800 151000 28900
rect 150900 28900 151000 29000
rect 150900 29000 151000 29100
rect 150900 29100 151000 29200
rect 150900 29200 151000 29300
rect 150900 29300 151000 29400
rect 150900 29400 151000 29500
rect 150900 29500 151000 29600
rect 150900 29600 151000 29700
rect 150900 29700 151000 29800
rect 150900 29800 151000 29900
rect 150900 29900 151000 30000
rect 150900 30000 151000 30100
rect 150900 30100 151000 30200
rect 150900 30200 151000 30300
rect 150900 30300 151000 30400
rect 150900 30400 151000 30500
rect 150900 30500 151000 30600
rect 150900 30600 151000 30700
rect 150900 30700 151000 30800
rect 150900 30800 151000 30900
rect 150900 30900 151000 31000
rect 150900 31000 151000 31100
rect 150900 31100 151000 31200
rect 150900 31200 151000 31300
rect 150900 31300 151000 31400
rect 150900 31400 151000 31500
rect 150900 31500 151000 31600
rect 150900 31600 151000 31700
rect 150900 31700 151000 31800
rect 150900 31800 151000 31900
rect 150900 31900 151000 32000
rect 150900 32000 151000 32100
rect 150900 32100 151000 32200
rect 150900 32200 151000 32300
rect 150900 32300 151000 32400
rect 150900 32400 151000 32500
rect 150900 32500 151000 32600
rect 150900 32600 151000 32700
rect 150900 32700 151000 32800
rect 150900 32800 151000 32900
rect 150900 32900 151000 33000
rect 150900 33000 151000 33100
rect 150900 33100 151000 33200
rect 150900 33200 151000 33300
rect 150900 33300 151000 33400
rect 150900 33400 151000 33500
rect 150900 33500 151000 33600
rect 150900 33600 151000 33700
rect 150900 33700 151000 33800
rect 150900 33800 151000 33900
rect 150900 33900 151000 34000
rect 150900 34000 151000 34100
rect 150900 34100 151000 34200
rect 150900 34200 151000 34300
rect 150900 34300 151000 34400
rect 150900 34400 151000 34500
rect 150900 34500 151000 34600
rect 150900 34600 151000 34700
rect 150900 34700 151000 34800
rect 150900 34800 151000 34900
rect 150900 34900 151000 35000
rect 150900 35000 151000 35100
rect 150900 35100 151000 35200
rect 150900 35200 151000 35300
rect 150900 35300 151000 35400
rect 150900 35400 151000 35500
rect 150900 35500 151000 35600
rect 150900 35600 151000 35700
rect 150900 35700 151000 35800
rect 150900 35800 151000 35900
rect 150900 35900 151000 36000
rect 150900 36000 151000 36100
rect 150900 36100 151000 36200
rect 150900 36200 151000 36300
rect 150900 36300 151000 36400
rect 150900 36400 151000 36500
rect 150900 36500 151000 36600
rect 150900 36600 151000 36700
rect 150900 36700 151000 36800
rect 150900 36800 151000 36900
rect 150900 36900 151000 37000
rect 150900 37000 151000 37100
rect 150900 37100 151000 37200
rect 150900 37200 151000 37300
rect 150900 37300 151000 37400
rect 150900 37400 151000 37500
rect 150900 37500 151000 37600
rect 150900 37600 151000 37700
rect 150900 37700 151000 37800
rect 150900 37800 151000 37900
rect 150900 37900 151000 38000
rect 150900 38000 151000 38100
rect 150900 38100 151000 38200
rect 151000 21200 151100 21300
rect 151000 21300 151100 21400
rect 151000 21400 151100 21500
rect 151000 21500 151100 21600
rect 151000 21600 151100 21700
rect 151000 21700 151100 21800
rect 151000 21800 151100 21900
rect 151000 21900 151100 22000
rect 151000 22000 151100 22100
rect 151000 22100 151100 22200
rect 151000 22200 151100 22300
rect 151000 22300 151100 22400
rect 151000 22400 151100 22500
rect 151000 22500 151100 22600
rect 151000 22600 151100 22700
rect 151000 22700 151100 22800
rect 151000 22800 151100 22900
rect 151000 22900 151100 23000
rect 151000 23000 151100 23100
rect 151000 23100 151100 23200
rect 151000 23200 151100 23300
rect 151000 23300 151100 23400
rect 151000 23400 151100 23500
rect 151000 23500 151100 23600
rect 151000 23600 151100 23700
rect 151000 23700 151100 23800
rect 151000 23800 151100 23900
rect 151000 23900 151100 24000
rect 151000 24000 151100 24100
rect 151000 24100 151100 24200
rect 151000 24200 151100 24300
rect 151000 24300 151100 24400
rect 151000 24400 151100 24500
rect 151000 24500 151100 24600
rect 151000 24600 151100 24700
rect 151000 24700 151100 24800
rect 151000 24800 151100 24900
rect 151000 24900 151100 25000
rect 151000 25000 151100 25100
rect 151000 25100 151100 25200
rect 151000 25200 151100 25300
rect 151000 25300 151100 25400
rect 151000 25400 151100 25500
rect 151000 25500 151100 25600
rect 151000 25600 151100 25700
rect 151000 25700 151100 25800
rect 151000 25800 151100 25900
rect 151000 25900 151100 26000
rect 151000 26000 151100 26100
rect 151000 26100 151100 26200
rect 151000 26200 151100 26300
rect 151000 26300 151100 26400
rect 151000 26400 151100 26500
rect 151000 26500 151100 26600
rect 151000 26600 151100 26700
rect 151000 26700 151100 26800
rect 151000 26800 151100 26900
rect 151000 26900 151100 27000
rect 151000 27000 151100 27100
rect 151000 27100 151100 27200
rect 151000 27200 151100 27300
rect 151000 27300 151100 27400
rect 151000 27400 151100 27500
rect 151000 27500 151100 27600
rect 151000 27600 151100 27700
rect 151000 27700 151100 27800
rect 151000 27800 151100 27900
rect 151000 27900 151100 28000
rect 151000 28000 151100 28100
rect 151000 28100 151100 28200
rect 151000 28200 151100 28300
rect 151000 28300 151100 28400
rect 151000 28400 151100 28500
rect 151000 28500 151100 28600
rect 151000 28600 151100 28700
rect 151000 28700 151100 28800
rect 151000 28800 151100 28900
rect 151000 28900 151100 29000
rect 151000 29000 151100 29100
rect 151000 29100 151100 29200
rect 151000 29200 151100 29300
rect 151000 29300 151100 29400
rect 151000 29400 151100 29500
rect 151000 29500 151100 29600
rect 151000 29600 151100 29700
rect 151000 29700 151100 29800
rect 151000 29800 151100 29900
rect 151000 29900 151100 30000
rect 151000 30000 151100 30100
rect 151000 30100 151100 30200
rect 151000 30200 151100 30300
rect 151000 30300 151100 30400
rect 151000 30400 151100 30500
rect 151000 30500 151100 30600
rect 151000 30600 151100 30700
rect 151000 30700 151100 30800
rect 151000 30800 151100 30900
rect 151000 30900 151100 31000
rect 151000 31000 151100 31100
rect 151000 31100 151100 31200
rect 151000 31200 151100 31300
rect 151000 31300 151100 31400
rect 151000 31400 151100 31500
rect 151000 31500 151100 31600
rect 151000 31600 151100 31700
rect 151000 31700 151100 31800
rect 151000 31800 151100 31900
rect 151000 31900 151100 32000
rect 151000 32000 151100 32100
rect 151000 32100 151100 32200
rect 151000 32200 151100 32300
rect 151000 32300 151100 32400
rect 151000 32400 151100 32500
rect 151000 32500 151100 32600
rect 151000 32600 151100 32700
rect 151000 32700 151100 32800
rect 151000 32800 151100 32900
rect 151000 32900 151100 33000
rect 151000 33000 151100 33100
rect 151000 33100 151100 33200
rect 151000 33200 151100 33300
rect 151000 33300 151100 33400
rect 151000 33400 151100 33500
rect 151000 33500 151100 33600
rect 151000 33600 151100 33700
rect 151000 33700 151100 33800
rect 151000 33800 151100 33900
rect 151000 33900 151100 34000
rect 151000 34000 151100 34100
rect 151000 34100 151100 34200
rect 151000 34200 151100 34300
rect 151000 34300 151100 34400
rect 151000 34400 151100 34500
rect 151000 34500 151100 34600
rect 151000 34600 151100 34700
rect 151000 34700 151100 34800
rect 151000 34800 151100 34900
rect 151000 34900 151100 35000
rect 151000 35000 151100 35100
rect 151000 35100 151100 35200
rect 151000 35200 151100 35300
rect 151000 35300 151100 35400
rect 151000 35400 151100 35500
rect 151000 35500 151100 35600
rect 151000 35600 151100 35700
rect 151000 35700 151100 35800
rect 151000 35800 151100 35900
rect 151000 35900 151100 36000
rect 151000 36000 151100 36100
rect 151000 36100 151100 36200
rect 151000 36200 151100 36300
rect 151000 36300 151100 36400
rect 151000 36400 151100 36500
rect 151000 36500 151100 36600
rect 151000 36600 151100 36700
rect 151000 36700 151100 36800
rect 151000 36800 151100 36900
rect 151000 36900 151100 37000
rect 151000 37000 151100 37100
rect 151000 37100 151100 37200
rect 151000 37200 151100 37300
rect 151000 37300 151100 37400
rect 151000 37400 151100 37500
rect 151000 37500 151100 37600
rect 151000 37600 151100 37700
rect 151000 37700 151100 37800
rect 151000 37800 151100 37900
rect 151000 37900 151100 38000
rect 151000 38000 151100 38100
rect 151000 38100 151100 38200
rect 151100 21200 151200 21300
rect 151100 21300 151200 21400
rect 151100 21400 151200 21500
rect 151100 21500 151200 21600
rect 151100 21600 151200 21700
rect 151100 21700 151200 21800
rect 151100 21800 151200 21900
rect 151100 21900 151200 22000
rect 151100 22000 151200 22100
rect 151100 22100 151200 22200
rect 151100 22200 151200 22300
rect 151100 22300 151200 22400
rect 151100 22400 151200 22500
rect 151100 22500 151200 22600
rect 151100 22600 151200 22700
rect 151100 22700 151200 22800
rect 151100 22800 151200 22900
rect 151100 22900 151200 23000
rect 151100 23000 151200 23100
rect 151100 23100 151200 23200
rect 151100 23200 151200 23300
rect 151100 23300 151200 23400
rect 151100 23400 151200 23500
rect 151100 23500 151200 23600
rect 151100 23600 151200 23700
rect 151100 23700 151200 23800
rect 151100 23800 151200 23900
rect 151100 23900 151200 24000
rect 151100 24000 151200 24100
rect 151100 24100 151200 24200
rect 151100 24200 151200 24300
rect 151100 24300 151200 24400
rect 151100 24400 151200 24500
rect 151100 24500 151200 24600
rect 151100 24600 151200 24700
rect 151100 24700 151200 24800
rect 151100 24800 151200 24900
rect 151100 24900 151200 25000
rect 151100 25000 151200 25100
rect 151100 25100 151200 25200
rect 151100 25200 151200 25300
rect 151100 25300 151200 25400
rect 151100 25400 151200 25500
rect 151100 25500 151200 25600
rect 151100 25600 151200 25700
rect 151100 25700 151200 25800
rect 151100 25800 151200 25900
rect 151100 25900 151200 26000
rect 151100 26000 151200 26100
rect 151100 26100 151200 26200
rect 151100 26200 151200 26300
rect 151100 26300 151200 26400
rect 151100 26400 151200 26500
rect 151100 26500 151200 26600
rect 151100 26600 151200 26700
rect 151100 26700 151200 26800
rect 151100 26800 151200 26900
rect 151100 26900 151200 27000
rect 151100 27000 151200 27100
rect 151100 27100 151200 27200
rect 151100 27200 151200 27300
rect 151100 27300 151200 27400
rect 151100 27400 151200 27500
rect 151100 27500 151200 27600
rect 151100 27600 151200 27700
rect 151100 27700 151200 27800
rect 151100 27800 151200 27900
rect 151100 27900 151200 28000
rect 151100 28000 151200 28100
rect 151100 28100 151200 28200
rect 151100 28200 151200 28300
rect 151100 28300 151200 28400
rect 151100 28400 151200 28500
rect 151100 28500 151200 28600
rect 151100 28600 151200 28700
rect 151100 28700 151200 28800
rect 151100 28800 151200 28900
rect 151100 28900 151200 29000
rect 151100 29000 151200 29100
rect 151100 29100 151200 29200
rect 151100 29200 151200 29300
rect 151100 29300 151200 29400
rect 151100 29400 151200 29500
rect 151100 29500 151200 29600
rect 151100 29600 151200 29700
rect 151100 29700 151200 29800
rect 151100 29800 151200 29900
rect 151100 29900 151200 30000
rect 151100 30000 151200 30100
rect 151100 30100 151200 30200
rect 151100 30200 151200 30300
rect 151100 30300 151200 30400
rect 151100 30400 151200 30500
rect 151100 30500 151200 30600
rect 151100 30600 151200 30700
rect 151100 30700 151200 30800
rect 151100 30800 151200 30900
rect 151100 30900 151200 31000
rect 151100 31000 151200 31100
rect 151100 31100 151200 31200
rect 151100 31200 151200 31300
rect 151100 31300 151200 31400
rect 151100 31400 151200 31500
rect 151100 31500 151200 31600
rect 151100 31600 151200 31700
rect 151100 31700 151200 31800
rect 151100 31800 151200 31900
rect 151100 31900 151200 32000
rect 151100 32000 151200 32100
rect 151100 32100 151200 32200
rect 151100 32200 151200 32300
rect 151100 32300 151200 32400
rect 151100 32400 151200 32500
rect 151100 32500 151200 32600
rect 151100 32600 151200 32700
rect 151100 32700 151200 32800
rect 151100 32800 151200 32900
rect 151100 32900 151200 33000
rect 151100 33000 151200 33100
rect 151100 33100 151200 33200
rect 151100 33200 151200 33300
rect 151100 33300 151200 33400
rect 151100 33400 151200 33500
rect 151100 33500 151200 33600
rect 151100 33600 151200 33700
rect 151100 33700 151200 33800
rect 151100 33800 151200 33900
rect 151100 33900 151200 34000
rect 151100 34000 151200 34100
rect 151100 34100 151200 34200
rect 151100 34200 151200 34300
rect 151100 34300 151200 34400
rect 151100 34400 151200 34500
rect 151100 34500 151200 34600
rect 151100 34600 151200 34700
rect 151100 34700 151200 34800
rect 151100 34800 151200 34900
rect 151100 34900 151200 35000
rect 151100 35000 151200 35100
rect 151100 35100 151200 35200
rect 151100 35200 151200 35300
rect 151100 35300 151200 35400
rect 151100 35400 151200 35500
rect 151100 35500 151200 35600
rect 151100 35600 151200 35700
rect 151100 35700 151200 35800
rect 151100 35800 151200 35900
rect 151100 35900 151200 36000
rect 151100 36000 151200 36100
rect 151100 36100 151200 36200
rect 151100 36200 151200 36300
rect 151100 36300 151200 36400
rect 151100 36400 151200 36500
rect 151100 36500 151200 36600
rect 151100 36600 151200 36700
rect 151100 36700 151200 36800
rect 151100 36800 151200 36900
rect 151100 36900 151200 37000
rect 151100 37000 151200 37100
rect 151100 37100 151200 37200
rect 151100 37200 151200 37300
rect 151100 37300 151200 37400
rect 151100 37400 151200 37500
rect 151100 37500 151200 37600
rect 151100 37600 151200 37700
rect 151100 37700 151200 37800
rect 151100 37800 151200 37900
rect 151100 37900 151200 38000
rect 151100 38000 151200 38100
rect 151100 38100 151200 38200
rect 151100 38200 151200 38300
rect 151200 21200 151300 21300
rect 151200 21300 151300 21400
rect 151200 21400 151300 21500
rect 151200 21500 151300 21600
rect 151200 21600 151300 21700
rect 151200 21700 151300 21800
rect 151200 21800 151300 21900
rect 151200 21900 151300 22000
rect 151200 22000 151300 22100
rect 151200 22100 151300 22200
rect 151200 22200 151300 22300
rect 151200 22300 151300 22400
rect 151200 22400 151300 22500
rect 151200 22500 151300 22600
rect 151200 22600 151300 22700
rect 151200 22700 151300 22800
rect 151200 22800 151300 22900
rect 151200 22900 151300 23000
rect 151200 23000 151300 23100
rect 151200 23100 151300 23200
rect 151200 23200 151300 23300
rect 151200 23300 151300 23400
rect 151200 23400 151300 23500
rect 151200 23500 151300 23600
rect 151200 23600 151300 23700
rect 151200 23700 151300 23800
rect 151200 23800 151300 23900
rect 151200 23900 151300 24000
rect 151200 24000 151300 24100
rect 151200 24100 151300 24200
rect 151200 24200 151300 24300
rect 151200 24300 151300 24400
rect 151200 24400 151300 24500
rect 151200 24500 151300 24600
rect 151200 24600 151300 24700
rect 151200 24700 151300 24800
rect 151200 24800 151300 24900
rect 151200 24900 151300 25000
rect 151200 25000 151300 25100
rect 151200 25100 151300 25200
rect 151200 25200 151300 25300
rect 151200 25300 151300 25400
rect 151200 25400 151300 25500
rect 151200 25500 151300 25600
rect 151200 25600 151300 25700
rect 151200 25700 151300 25800
rect 151200 25800 151300 25900
rect 151200 25900 151300 26000
rect 151200 26000 151300 26100
rect 151200 26100 151300 26200
rect 151200 26200 151300 26300
rect 151200 26300 151300 26400
rect 151200 26400 151300 26500
rect 151200 26500 151300 26600
rect 151200 26600 151300 26700
rect 151200 26700 151300 26800
rect 151200 26800 151300 26900
rect 151200 26900 151300 27000
rect 151200 27000 151300 27100
rect 151200 27100 151300 27200
rect 151200 27200 151300 27300
rect 151200 27300 151300 27400
rect 151200 27400 151300 27500
rect 151200 27500 151300 27600
rect 151200 27600 151300 27700
rect 151200 27700 151300 27800
rect 151200 27800 151300 27900
rect 151200 27900 151300 28000
rect 151200 28000 151300 28100
rect 151200 28100 151300 28200
rect 151200 28200 151300 28300
rect 151200 28300 151300 28400
rect 151200 28400 151300 28500
rect 151200 28500 151300 28600
rect 151200 28600 151300 28700
rect 151200 28700 151300 28800
rect 151200 28800 151300 28900
rect 151200 28900 151300 29000
rect 151200 29000 151300 29100
rect 151200 29100 151300 29200
rect 151200 29200 151300 29300
rect 151200 29300 151300 29400
rect 151200 29400 151300 29500
rect 151200 29500 151300 29600
rect 151200 29600 151300 29700
rect 151200 29700 151300 29800
rect 151200 29800 151300 29900
rect 151200 29900 151300 30000
rect 151200 30000 151300 30100
rect 151200 30100 151300 30200
rect 151200 30200 151300 30300
rect 151200 30300 151300 30400
rect 151200 30400 151300 30500
rect 151200 30500 151300 30600
rect 151200 30600 151300 30700
rect 151200 30700 151300 30800
rect 151200 30800 151300 30900
rect 151200 30900 151300 31000
rect 151200 31000 151300 31100
rect 151200 31100 151300 31200
rect 151200 31200 151300 31300
rect 151200 31300 151300 31400
rect 151200 31400 151300 31500
rect 151200 31500 151300 31600
rect 151200 31600 151300 31700
rect 151200 31700 151300 31800
rect 151200 31800 151300 31900
rect 151200 31900 151300 32000
rect 151200 32000 151300 32100
rect 151200 32100 151300 32200
rect 151200 32200 151300 32300
rect 151200 32300 151300 32400
rect 151200 32400 151300 32500
rect 151200 32500 151300 32600
rect 151200 32600 151300 32700
rect 151200 32700 151300 32800
rect 151200 32800 151300 32900
rect 151200 32900 151300 33000
rect 151200 33000 151300 33100
rect 151200 33100 151300 33200
rect 151200 33200 151300 33300
rect 151200 33300 151300 33400
rect 151200 33400 151300 33500
rect 151200 33500 151300 33600
rect 151200 33600 151300 33700
rect 151200 33700 151300 33800
rect 151200 33800 151300 33900
rect 151200 33900 151300 34000
rect 151200 34000 151300 34100
rect 151200 34100 151300 34200
rect 151200 34200 151300 34300
rect 151200 34300 151300 34400
rect 151200 34400 151300 34500
rect 151200 34500 151300 34600
rect 151200 34600 151300 34700
rect 151200 34700 151300 34800
rect 151200 34800 151300 34900
rect 151200 34900 151300 35000
rect 151200 35000 151300 35100
rect 151200 35100 151300 35200
rect 151200 35200 151300 35300
rect 151200 35300 151300 35400
rect 151200 35400 151300 35500
rect 151200 35500 151300 35600
rect 151200 35600 151300 35700
rect 151200 35700 151300 35800
rect 151200 35800 151300 35900
rect 151200 35900 151300 36000
rect 151200 36000 151300 36100
rect 151200 36100 151300 36200
rect 151200 36200 151300 36300
rect 151200 36300 151300 36400
rect 151200 36400 151300 36500
rect 151200 36500 151300 36600
rect 151200 36600 151300 36700
rect 151200 36700 151300 36800
rect 151200 36800 151300 36900
rect 151200 36900 151300 37000
rect 151200 37000 151300 37100
rect 151200 37100 151300 37200
rect 151200 37200 151300 37300
rect 151200 37300 151300 37400
rect 151200 37400 151300 37500
rect 151200 37500 151300 37600
rect 151200 37600 151300 37700
rect 151200 37700 151300 37800
rect 151200 37800 151300 37900
rect 151200 37900 151300 38000
rect 151200 38000 151300 38100
rect 151200 38100 151300 38200
rect 151200 38200 151300 38300
rect 151300 21100 151400 21200
rect 151300 21200 151400 21300
rect 151300 21300 151400 21400
rect 151300 21400 151400 21500
rect 151300 21500 151400 21600
rect 151300 21600 151400 21700
rect 151300 21700 151400 21800
rect 151300 21800 151400 21900
rect 151300 21900 151400 22000
rect 151300 22000 151400 22100
rect 151300 22100 151400 22200
rect 151300 22200 151400 22300
rect 151300 22300 151400 22400
rect 151300 22400 151400 22500
rect 151300 22500 151400 22600
rect 151300 22600 151400 22700
rect 151300 22700 151400 22800
rect 151300 22800 151400 22900
rect 151300 22900 151400 23000
rect 151300 23000 151400 23100
rect 151300 23100 151400 23200
rect 151300 23200 151400 23300
rect 151300 23300 151400 23400
rect 151300 23400 151400 23500
rect 151300 23500 151400 23600
rect 151300 23600 151400 23700
rect 151300 23700 151400 23800
rect 151300 23800 151400 23900
rect 151300 23900 151400 24000
rect 151300 24000 151400 24100
rect 151300 24100 151400 24200
rect 151300 24200 151400 24300
rect 151300 24300 151400 24400
rect 151300 24400 151400 24500
rect 151300 24500 151400 24600
rect 151300 24600 151400 24700
rect 151300 24700 151400 24800
rect 151300 24800 151400 24900
rect 151300 24900 151400 25000
rect 151300 25000 151400 25100
rect 151300 25100 151400 25200
rect 151300 25200 151400 25300
rect 151300 25300 151400 25400
rect 151300 25400 151400 25500
rect 151300 25500 151400 25600
rect 151300 25600 151400 25700
rect 151300 25700 151400 25800
rect 151300 25800 151400 25900
rect 151300 25900 151400 26000
rect 151300 26000 151400 26100
rect 151300 26100 151400 26200
rect 151300 26200 151400 26300
rect 151300 26300 151400 26400
rect 151300 26400 151400 26500
rect 151300 26500 151400 26600
rect 151300 26600 151400 26700
rect 151300 26700 151400 26800
rect 151300 26800 151400 26900
rect 151300 26900 151400 27000
rect 151300 27000 151400 27100
rect 151300 27100 151400 27200
rect 151300 27200 151400 27300
rect 151300 27300 151400 27400
rect 151300 27400 151400 27500
rect 151300 27500 151400 27600
rect 151300 27600 151400 27700
rect 151300 27700 151400 27800
rect 151300 27800 151400 27900
rect 151300 27900 151400 28000
rect 151300 28000 151400 28100
rect 151300 28100 151400 28200
rect 151300 28200 151400 28300
rect 151300 28300 151400 28400
rect 151300 28400 151400 28500
rect 151300 28500 151400 28600
rect 151300 28600 151400 28700
rect 151300 28700 151400 28800
rect 151300 28800 151400 28900
rect 151300 28900 151400 29000
rect 151300 29000 151400 29100
rect 151300 29100 151400 29200
rect 151300 29200 151400 29300
rect 151300 29300 151400 29400
rect 151300 29400 151400 29500
rect 151300 29500 151400 29600
rect 151300 29600 151400 29700
rect 151300 29700 151400 29800
rect 151300 29800 151400 29900
rect 151300 29900 151400 30000
rect 151300 30000 151400 30100
rect 151300 30100 151400 30200
rect 151300 30200 151400 30300
rect 151300 30300 151400 30400
rect 151300 30400 151400 30500
rect 151300 30500 151400 30600
rect 151300 30600 151400 30700
rect 151300 30700 151400 30800
rect 151300 30800 151400 30900
rect 151300 30900 151400 31000
rect 151300 31000 151400 31100
rect 151300 31100 151400 31200
rect 151300 31200 151400 31300
rect 151300 31300 151400 31400
rect 151300 31400 151400 31500
rect 151300 31500 151400 31600
rect 151300 31600 151400 31700
rect 151300 31700 151400 31800
rect 151300 31800 151400 31900
rect 151300 31900 151400 32000
rect 151300 32000 151400 32100
rect 151300 32100 151400 32200
rect 151300 32200 151400 32300
rect 151300 32300 151400 32400
rect 151300 32400 151400 32500
rect 151300 32500 151400 32600
rect 151300 32600 151400 32700
rect 151300 32700 151400 32800
rect 151300 32800 151400 32900
rect 151300 32900 151400 33000
rect 151300 33000 151400 33100
rect 151300 33100 151400 33200
rect 151300 33200 151400 33300
rect 151300 33300 151400 33400
rect 151300 33400 151400 33500
rect 151300 33500 151400 33600
rect 151300 33600 151400 33700
rect 151300 33700 151400 33800
rect 151300 33800 151400 33900
rect 151300 33900 151400 34000
rect 151300 34000 151400 34100
rect 151300 34100 151400 34200
rect 151300 34200 151400 34300
rect 151300 34300 151400 34400
rect 151300 34400 151400 34500
rect 151300 34500 151400 34600
rect 151300 34600 151400 34700
rect 151300 34700 151400 34800
rect 151300 34800 151400 34900
rect 151300 34900 151400 35000
rect 151300 35000 151400 35100
rect 151300 35100 151400 35200
rect 151300 35200 151400 35300
rect 151300 35300 151400 35400
rect 151300 35400 151400 35500
rect 151300 35500 151400 35600
rect 151300 35600 151400 35700
rect 151300 35700 151400 35800
rect 151300 35800 151400 35900
rect 151300 35900 151400 36000
rect 151300 36000 151400 36100
rect 151300 36100 151400 36200
rect 151300 36200 151400 36300
rect 151300 36300 151400 36400
rect 151300 36400 151400 36500
rect 151300 36500 151400 36600
rect 151300 36600 151400 36700
rect 151300 36700 151400 36800
rect 151300 36800 151400 36900
rect 151300 36900 151400 37000
rect 151300 37000 151400 37100
rect 151300 37100 151400 37200
rect 151300 37200 151400 37300
rect 151300 37300 151400 37400
rect 151300 37400 151400 37500
rect 151300 37500 151400 37600
rect 151300 37600 151400 37700
rect 151300 37700 151400 37800
rect 151300 37800 151400 37900
rect 151300 37900 151400 38000
rect 151300 38000 151400 38100
rect 151300 38100 151400 38200
rect 151300 38200 151400 38300
rect 151400 21100 151500 21200
rect 151400 21200 151500 21300
rect 151400 21300 151500 21400
rect 151400 21400 151500 21500
rect 151400 21500 151500 21600
rect 151400 21600 151500 21700
rect 151400 21700 151500 21800
rect 151400 21800 151500 21900
rect 151400 21900 151500 22000
rect 151400 22000 151500 22100
rect 151400 22100 151500 22200
rect 151400 22200 151500 22300
rect 151400 22300 151500 22400
rect 151400 22400 151500 22500
rect 151400 22500 151500 22600
rect 151400 22600 151500 22700
rect 151400 22700 151500 22800
rect 151400 22800 151500 22900
rect 151400 22900 151500 23000
rect 151400 23000 151500 23100
rect 151400 23100 151500 23200
rect 151400 23200 151500 23300
rect 151400 23300 151500 23400
rect 151400 23400 151500 23500
rect 151400 23500 151500 23600
rect 151400 23600 151500 23700
rect 151400 23700 151500 23800
rect 151400 23800 151500 23900
rect 151400 23900 151500 24000
rect 151400 24000 151500 24100
rect 151400 24100 151500 24200
rect 151400 24200 151500 24300
rect 151400 24300 151500 24400
rect 151400 24400 151500 24500
rect 151400 24500 151500 24600
rect 151400 24600 151500 24700
rect 151400 24700 151500 24800
rect 151400 24800 151500 24900
rect 151400 24900 151500 25000
rect 151400 25000 151500 25100
rect 151400 25100 151500 25200
rect 151400 25200 151500 25300
rect 151400 25300 151500 25400
rect 151400 25400 151500 25500
rect 151400 25500 151500 25600
rect 151400 25600 151500 25700
rect 151400 25700 151500 25800
rect 151400 25800 151500 25900
rect 151400 25900 151500 26000
rect 151400 26000 151500 26100
rect 151400 26100 151500 26200
rect 151400 26200 151500 26300
rect 151400 26300 151500 26400
rect 151400 26400 151500 26500
rect 151400 26500 151500 26600
rect 151400 26600 151500 26700
rect 151400 26700 151500 26800
rect 151400 26800 151500 26900
rect 151400 26900 151500 27000
rect 151400 27000 151500 27100
rect 151400 27100 151500 27200
rect 151400 27200 151500 27300
rect 151400 27300 151500 27400
rect 151400 27400 151500 27500
rect 151400 27500 151500 27600
rect 151400 27600 151500 27700
rect 151400 27700 151500 27800
rect 151400 27800 151500 27900
rect 151400 27900 151500 28000
rect 151400 28000 151500 28100
rect 151400 28100 151500 28200
rect 151400 28200 151500 28300
rect 151400 28300 151500 28400
rect 151400 28400 151500 28500
rect 151400 28500 151500 28600
rect 151400 28600 151500 28700
rect 151400 28700 151500 28800
rect 151400 28800 151500 28900
rect 151400 28900 151500 29000
rect 151400 29000 151500 29100
rect 151400 29100 151500 29200
rect 151400 29200 151500 29300
rect 151400 29300 151500 29400
rect 151400 29400 151500 29500
rect 151400 29500 151500 29600
rect 151400 29600 151500 29700
rect 151400 29700 151500 29800
rect 151400 29800 151500 29900
rect 151400 29900 151500 30000
rect 151400 30000 151500 30100
rect 151400 30100 151500 30200
rect 151400 30200 151500 30300
rect 151400 30300 151500 30400
rect 151400 30400 151500 30500
rect 151400 30500 151500 30600
rect 151400 30600 151500 30700
rect 151400 30700 151500 30800
rect 151400 30800 151500 30900
rect 151400 30900 151500 31000
rect 151400 31000 151500 31100
rect 151400 31100 151500 31200
rect 151400 31200 151500 31300
rect 151400 31300 151500 31400
rect 151400 31400 151500 31500
rect 151400 31500 151500 31600
rect 151400 31600 151500 31700
rect 151400 31700 151500 31800
rect 151400 31800 151500 31900
rect 151400 31900 151500 32000
rect 151400 32000 151500 32100
rect 151400 32100 151500 32200
rect 151400 32200 151500 32300
rect 151400 32300 151500 32400
rect 151400 32400 151500 32500
rect 151400 32500 151500 32600
rect 151400 32600 151500 32700
rect 151400 32700 151500 32800
rect 151400 32800 151500 32900
rect 151400 32900 151500 33000
rect 151400 33000 151500 33100
rect 151400 33100 151500 33200
rect 151400 33200 151500 33300
rect 151400 33300 151500 33400
rect 151400 33400 151500 33500
rect 151400 33500 151500 33600
rect 151400 33600 151500 33700
rect 151400 33700 151500 33800
rect 151400 33800 151500 33900
rect 151400 33900 151500 34000
rect 151400 34000 151500 34100
rect 151400 34100 151500 34200
rect 151400 34200 151500 34300
rect 151400 34300 151500 34400
rect 151400 34400 151500 34500
rect 151400 34500 151500 34600
rect 151400 34600 151500 34700
rect 151400 34700 151500 34800
rect 151400 34800 151500 34900
rect 151400 34900 151500 35000
rect 151400 35000 151500 35100
rect 151400 35100 151500 35200
rect 151400 35200 151500 35300
rect 151400 35300 151500 35400
rect 151400 35400 151500 35500
rect 151400 35500 151500 35600
rect 151400 35600 151500 35700
rect 151400 35700 151500 35800
rect 151400 35800 151500 35900
rect 151400 35900 151500 36000
rect 151400 36000 151500 36100
rect 151400 36100 151500 36200
rect 151400 36200 151500 36300
rect 151400 36300 151500 36400
rect 151400 36400 151500 36500
rect 151400 36500 151500 36600
rect 151400 36600 151500 36700
rect 151400 36700 151500 36800
rect 151400 36800 151500 36900
rect 151400 36900 151500 37000
rect 151400 37000 151500 37100
rect 151400 37100 151500 37200
rect 151400 37200 151500 37300
rect 151400 37300 151500 37400
rect 151400 37400 151500 37500
rect 151400 37500 151500 37600
rect 151400 37600 151500 37700
rect 151400 37700 151500 37800
rect 151400 37800 151500 37900
rect 151400 37900 151500 38000
rect 151400 38000 151500 38100
rect 151400 38100 151500 38200
rect 151400 38200 151500 38300
rect 151500 21100 151600 21200
rect 151500 21200 151600 21300
rect 151500 21300 151600 21400
rect 151500 21400 151600 21500
rect 151500 21500 151600 21600
rect 151500 21600 151600 21700
rect 151500 21700 151600 21800
rect 151500 21800 151600 21900
rect 151500 21900 151600 22000
rect 151500 22000 151600 22100
rect 151500 22100 151600 22200
rect 151500 22200 151600 22300
rect 151500 22300 151600 22400
rect 151500 22400 151600 22500
rect 151500 22500 151600 22600
rect 151500 22600 151600 22700
rect 151500 22700 151600 22800
rect 151500 22800 151600 22900
rect 151500 22900 151600 23000
rect 151500 23000 151600 23100
rect 151500 23100 151600 23200
rect 151500 23200 151600 23300
rect 151500 23300 151600 23400
rect 151500 23400 151600 23500
rect 151500 23500 151600 23600
rect 151500 23600 151600 23700
rect 151500 23700 151600 23800
rect 151500 23800 151600 23900
rect 151500 23900 151600 24000
rect 151500 24000 151600 24100
rect 151500 24100 151600 24200
rect 151500 24200 151600 24300
rect 151500 24300 151600 24400
rect 151500 24400 151600 24500
rect 151500 24500 151600 24600
rect 151500 24600 151600 24700
rect 151500 24700 151600 24800
rect 151500 24800 151600 24900
rect 151500 24900 151600 25000
rect 151500 25000 151600 25100
rect 151500 25100 151600 25200
rect 151500 25200 151600 25300
rect 151500 25300 151600 25400
rect 151500 25400 151600 25500
rect 151500 25500 151600 25600
rect 151500 25600 151600 25700
rect 151500 25700 151600 25800
rect 151500 25800 151600 25900
rect 151500 25900 151600 26000
rect 151500 26000 151600 26100
rect 151500 26100 151600 26200
rect 151500 26200 151600 26300
rect 151500 26300 151600 26400
rect 151500 26400 151600 26500
rect 151500 26500 151600 26600
rect 151500 26600 151600 26700
rect 151500 26700 151600 26800
rect 151500 26800 151600 26900
rect 151500 26900 151600 27000
rect 151500 27000 151600 27100
rect 151500 27100 151600 27200
rect 151500 27200 151600 27300
rect 151500 27300 151600 27400
rect 151500 27400 151600 27500
rect 151500 27500 151600 27600
rect 151500 27600 151600 27700
rect 151500 27700 151600 27800
rect 151500 27800 151600 27900
rect 151500 27900 151600 28000
rect 151500 28000 151600 28100
rect 151500 28100 151600 28200
rect 151500 28200 151600 28300
rect 151500 28300 151600 28400
rect 151500 28400 151600 28500
rect 151500 28500 151600 28600
rect 151500 28600 151600 28700
rect 151500 28700 151600 28800
rect 151500 28800 151600 28900
rect 151500 28900 151600 29000
rect 151500 29000 151600 29100
rect 151500 29100 151600 29200
rect 151500 29200 151600 29300
rect 151500 29300 151600 29400
rect 151500 29400 151600 29500
rect 151500 29900 151600 30000
rect 151500 30000 151600 30100
rect 151500 30100 151600 30200
rect 151500 30200 151600 30300
rect 151500 30300 151600 30400
rect 151500 30400 151600 30500
rect 151500 30500 151600 30600
rect 151500 30600 151600 30700
rect 151500 30700 151600 30800
rect 151500 30800 151600 30900
rect 151500 30900 151600 31000
rect 151500 31000 151600 31100
rect 151500 31100 151600 31200
rect 151500 31200 151600 31300
rect 151500 31300 151600 31400
rect 151500 31400 151600 31500
rect 151500 31500 151600 31600
rect 151500 31600 151600 31700
rect 151500 31700 151600 31800
rect 151500 31800 151600 31900
rect 151500 31900 151600 32000
rect 151500 32000 151600 32100
rect 151500 32100 151600 32200
rect 151500 32200 151600 32300
rect 151500 32300 151600 32400
rect 151500 32400 151600 32500
rect 151500 32500 151600 32600
rect 151500 32600 151600 32700
rect 151500 32700 151600 32800
rect 151500 32800 151600 32900
rect 151500 32900 151600 33000
rect 151500 33000 151600 33100
rect 151500 33100 151600 33200
rect 151500 33200 151600 33300
rect 151500 33300 151600 33400
rect 151500 33400 151600 33500
rect 151500 33500 151600 33600
rect 151500 33600 151600 33700
rect 151500 33700 151600 33800
rect 151500 33800 151600 33900
rect 151500 33900 151600 34000
rect 151500 34000 151600 34100
rect 151500 34100 151600 34200
rect 151500 34200 151600 34300
rect 151500 34300 151600 34400
rect 151500 34400 151600 34500
rect 151500 34500 151600 34600
rect 151500 34600 151600 34700
rect 151500 34700 151600 34800
rect 151500 34800 151600 34900
rect 151500 34900 151600 35000
rect 151500 35000 151600 35100
rect 151500 35100 151600 35200
rect 151500 35200 151600 35300
rect 151500 35300 151600 35400
rect 151500 35400 151600 35500
rect 151500 35500 151600 35600
rect 151500 35600 151600 35700
rect 151500 35700 151600 35800
rect 151500 35800 151600 35900
rect 151500 35900 151600 36000
rect 151500 36000 151600 36100
rect 151500 36100 151600 36200
rect 151500 36200 151600 36300
rect 151500 36300 151600 36400
rect 151500 36400 151600 36500
rect 151500 36500 151600 36600
rect 151500 36600 151600 36700
rect 151500 36700 151600 36800
rect 151500 36800 151600 36900
rect 151500 36900 151600 37000
rect 151500 37000 151600 37100
rect 151500 37100 151600 37200
rect 151500 37200 151600 37300
rect 151500 37300 151600 37400
rect 151500 37400 151600 37500
rect 151500 37500 151600 37600
rect 151500 37600 151600 37700
rect 151500 37700 151600 37800
rect 151500 37800 151600 37900
rect 151500 37900 151600 38000
rect 151500 38000 151600 38100
rect 151500 38100 151600 38200
rect 151500 38200 151600 38300
rect 151500 38300 151600 38400
rect 151600 21200 151700 21300
rect 151600 21300 151700 21400
rect 151600 21400 151700 21500
rect 151600 21500 151700 21600
rect 151600 21600 151700 21700
rect 151600 21700 151700 21800
rect 151600 21800 151700 21900
rect 151600 21900 151700 22000
rect 151600 22000 151700 22100
rect 151600 22100 151700 22200
rect 151600 22200 151700 22300
rect 151600 22300 151700 22400
rect 151600 22400 151700 22500
rect 151600 22500 151700 22600
rect 151600 22600 151700 22700
rect 151600 22700 151700 22800
rect 151600 22800 151700 22900
rect 151600 22900 151700 23000
rect 151600 23000 151700 23100
rect 151600 23100 151700 23200
rect 151600 23200 151700 23300
rect 151600 23300 151700 23400
rect 151600 23400 151700 23500
rect 151600 23500 151700 23600
rect 151600 23600 151700 23700
rect 151600 23700 151700 23800
rect 151600 23800 151700 23900
rect 151600 23900 151700 24000
rect 151600 24000 151700 24100
rect 151600 24100 151700 24200
rect 151600 24200 151700 24300
rect 151600 24300 151700 24400
rect 151600 24400 151700 24500
rect 151600 24500 151700 24600
rect 151600 24600 151700 24700
rect 151600 24700 151700 24800
rect 151600 24800 151700 24900
rect 151600 24900 151700 25000
rect 151600 25000 151700 25100
rect 151600 25100 151700 25200
rect 151600 25200 151700 25300
rect 151600 25300 151700 25400
rect 151600 25400 151700 25500
rect 151600 25500 151700 25600
rect 151600 25600 151700 25700
rect 151600 25700 151700 25800
rect 151600 25800 151700 25900
rect 151600 25900 151700 26000
rect 151600 26000 151700 26100
rect 151600 26100 151700 26200
rect 151600 26200 151700 26300
rect 151600 26300 151700 26400
rect 151600 26400 151700 26500
rect 151600 26500 151700 26600
rect 151600 26600 151700 26700
rect 151600 26700 151700 26800
rect 151600 26800 151700 26900
rect 151600 26900 151700 27000
rect 151600 27000 151700 27100
rect 151600 27100 151700 27200
rect 151600 27200 151700 27300
rect 151600 27300 151700 27400
rect 151600 27400 151700 27500
rect 151600 27500 151700 27600
rect 151600 27600 151700 27700
rect 151600 27700 151700 27800
rect 151600 27800 151700 27900
rect 151600 27900 151700 28000
rect 151600 28000 151700 28100
rect 151600 28100 151700 28200
rect 151600 28200 151700 28300
rect 151600 28300 151700 28400
rect 151600 28400 151700 28500
rect 151600 28500 151700 28600
rect 151600 28600 151700 28700
rect 151600 28700 151700 28800
rect 151600 28800 151700 28900
rect 151600 28900 151700 29000
rect 151600 29000 151700 29100
rect 151600 29100 151700 29200
rect 151600 29200 151700 29300
rect 151600 30100 151700 30200
rect 151600 30200 151700 30300
rect 151600 30300 151700 30400
rect 151600 30400 151700 30500
rect 151600 30500 151700 30600
rect 151600 30600 151700 30700
rect 151600 30700 151700 30800
rect 151600 30800 151700 30900
rect 151600 30900 151700 31000
rect 151600 31000 151700 31100
rect 151600 31100 151700 31200
rect 151600 31200 151700 31300
rect 151600 31300 151700 31400
rect 151600 31400 151700 31500
rect 151600 31500 151700 31600
rect 151600 31600 151700 31700
rect 151600 31700 151700 31800
rect 151600 31800 151700 31900
rect 151600 31900 151700 32000
rect 151600 32000 151700 32100
rect 151600 32100 151700 32200
rect 151600 32200 151700 32300
rect 151600 32300 151700 32400
rect 151600 32400 151700 32500
rect 151600 32500 151700 32600
rect 151600 32600 151700 32700
rect 151600 32700 151700 32800
rect 151600 32800 151700 32900
rect 151600 32900 151700 33000
rect 151600 33000 151700 33100
rect 151600 33100 151700 33200
rect 151600 33200 151700 33300
rect 151600 33300 151700 33400
rect 151600 33400 151700 33500
rect 151600 33500 151700 33600
rect 151600 33600 151700 33700
rect 151600 33700 151700 33800
rect 151600 33800 151700 33900
rect 151600 33900 151700 34000
rect 151600 34000 151700 34100
rect 151600 34100 151700 34200
rect 151600 34200 151700 34300
rect 151600 34300 151700 34400
rect 151600 34400 151700 34500
rect 151600 34500 151700 34600
rect 151600 34600 151700 34700
rect 151600 34700 151700 34800
rect 151600 34800 151700 34900
rect 151600 34900 151700 35000
rect 151600 35000 151700 35100
rect 151600 35100 151700 35200
rect 151600 35200 151700 35300
rect 151600 35300 151700 35400
rect 151600 35400 151700 35500
rect 151600 35500 151700 35600
rect 151600 35600 151700 35700
rect 151600 35700 151700 35800
rect 151600 35800 151700 35900
rect 151600 35900 151700 36000
rect 151600 36000 151700 36100
rect 151600 36100 151700 36200
rect 151600 36200 151700 36300
rect 151600 36300 151700 36400
rect 151600 36400 151700 36500
rect 151600 36500 151700 36600
rect 151600 36600 151700 36700
rect 151600 36700 151700 36800
rect 151600 36800 151700 36900
rect 151600 36900 151700 37000
rect 151600 37000 151700 37100
rect 151600 37100 151700 37200
rect 151600 37200 151700 37300
rect 151600 37300 151700 37400
rect 151600 37400 151700 37500
rect 151600 37500 151700 37600
rect 151600 37600 151700 37700
rect 151600 37700 151700 37800
rect 151600 37800 151700 37900
rect 151600 37900 151700 38000
rect 151600 38000 151700 38100
rect 151600 38100 151700 38200
rect 151600 38200 151700 38300
rect 151700 21200 151800 21300
rect 151700 21300 151800 21400
rect 151700 21400 151800 21500
rect 151700 21500 151800 21600
rect 151700 21600 151800 21700
rect 151700 21700 151800 21800
rect 151700 21800 151800 21900
rect 151700 21900 151800 22000
rect 151700 22000 151800 22100
rect 151700 22100 151800 22200
rect 151700 22200 151800 22300
rect 151700 22300 151800 22400
rect 151700 22400 151800 22500
rect 151700 22500 151800 22600
rect 151700 22600 151800 22700
rect 151700 22700 151800 22800
rect 151700 22800 151800 22900
rect 151700 22900 151800 23000
rect 151700 23000 151800 23100
rect 151700 23100 151800 23200
rect 151700 23200 151800 23300
rect 151700 23300 151800 23400
rect 151700 23400 151800 23500
rect 151700 23500 151800 23600
rect 151700 23600 151800 23700
rect 151700 23700 151800 23800
rect 151700 23800 151800 23900
rect 151700 23900 151800 24000
rect 151700 24000 151800 24100
rect 151700 24100 151800 24200
rect 151700 24200 151800 24300
rect 151700 24300 151800 24400
rect 151700 24400 151800 24500
rect 151700 24500 151800 24600
rect 151700 24600 151800 24700
rect 151700 24700 151800 24800
rect 151700 24800 151800 24900
rect 151700 24900 151800 25000
rect 151700 25000 151800 25100
rect 151700 25100 151800 25200
rect 151700 25200 151800 25300
rect 151700 25300 151800 25400
rect 151700 25400 151800 25500
rect 151700 25500 151800 25600
rect 151700 25600 151800 25700
rect 151700 25700 151800 25800
rect 151700 25800 151800 25900
rect 151700 25900 151800 26000
rect 151700 26000 151800 26100
rect 151700 26100 151800 26200
rect 151700 26200 151800 26300
rect 151700 26300 151800 26400
rect 151700 26400 151800 26500
rect 151700 26500 151800 26600
rect 151700 26600 151800 26700
rect 151700 26700 151800 26800
rect 151700 26800 151800 26900
rect 151700 26900 151800 27000
rect 151700 27000 151800 27100
rect 151700 27100 151800 27200
rect 151700 27200 151800 27300
rect 151700 27300 151800 27400
rect 151700 27400 151800 27500
rect 151700 27500 151800 27600
rect 151700 27600 151800 27700
rect 151700 27700 151800 27800
rect 151700 27800 151800 27900
rect 151700 27900 151800 28000
rect 151700 28000 151800 28100
rect 151700 28100 151800 28200
rect 151700 28200 151800 28300
rect 151700 28300 151800 28400
rect 151700 28400 151800 28500
rect 151700 28500 151800 28600
rect 151700 28600 151800 28700
rect 151700 28700 151800 28800
rect 151700 28800 151800 28900
rect 151700 28900 151800 29000
rect 151700 29000 151800 29100
rect 151700 30300 151800 30400
rect 151700 30400 151800 30500
rect 151700 30500 151800 30600
rect 151700 30600 151800 30700
rect 151700 30700 151800 30800
rect 151700 30800 151800 30900
rect 151700 30900 151800 31000
rect 151700 31000 151800 31100
rect 151700 31100 151800 31200
rect 151700 31200 151800 31300
rect 151700 31300 151800 31400
rect 151700 31400 151800 31500
rect 151700 31500 151800 31600
rect 151700 31600 151800 31700
rect 151700 31700 151800 31800
rect 151700 31800 151800 31900
rect 151700 31900 151800 32000
rect 151700 32000 151800 32100
rect 151700 32100 151800 32200
rect 151700 32200 151800 32300
rect 151700 32300 151800 32400
rect 151700 32400 151800 32500
rect 151700 32500 151800 32600
rect 151700 32600 151800 32700
rect 151700 32700 151800 32800
rect 151700 32800 151800 32900
rect 151700 32900 151800 33000
rect 151700 33000 151800 33100
rect 151700 33100 151800 33200
rect 151700 33200 151800 33300
rect 151700 33300 151800 33400
rect 151700 33400 151800 33500
rect 151700 33500 151800 33600
rect 151700 33600 151800 33700
rect 151700 33700 151800 33800
rect 151700 33800 151800 33900
rect 151700 33900 151800 34000
rect 151700 34000 151800 34100
rect 151700 34100 151800 34200
rect 151700 34200 151800 34300
rect 151700 34300 151800 34400
rect 151700 34400 151800 34500
rect 151700 34500 151800 34600
rect 151700 34600 151800 34700
rect 151700 34700 151800 34800
rect 151700 34800 151800 34900
rect 151700 34900 151800 35000
rect 151700 35000 151800 35100
rect 151700 35100 151800 35200
rect 151700 35200 151800 35300
rect 151700 35300 151800 35400
rect 151700 35400 151800 35500
rect 151700 35500 151800 35600
rect 151700 35600 151800 35700
rect 151700 35700 151800 35800
rect 151700 35800 151800 35900
rect 151700 35900 151800 36000
rect 151700 36000 151800 36100
rect 151700 36100 151800 36200
rect 151700 36200 151800 36300
rect 151700 36300 151800 36400
rect 151700 36400 151800 36500
rect 151700 36500 151800 36600
rect 151700 36600 151800 36700
rect 151700 36700 151800 36800
rect 151700 36800 151800 36900
rect 151700 36900 151800 37000
rect 151700 37000 151800 37100
rect 151700 37100 151800 37200
rect 151700 37200 151800 37300
rect 151700 37300 151800 37400
rect 151700 37400 151800 37500
rect 151700 37500 151800 37600
rect 151700 37600 151800 37700
rect 151700 37700 151800 37800
rect 151700 37800 151800 37900
rect 151700 37900 151800 38000
rect 151700 38000 151800 38100
rect 151700 38100 151800 38200
rect 151700 38200 151800 38300
rect 151800 21200 151900 21300
rect 151800 21300 151900 21400
rect 151800 21400 151900 21500
rect 151800 21500 151900 21600
rect 151800 21600 151900 21700
rect 151800 21700 151900 21800
rect 151800 21800 151900 21900
rect 151800 21900 151900 22000
rect 151800 22000 151900 22100
rect 151800 22100 151900 22200
rect 151800 22200 151900 22300
rect 151800 22300 151900 22400
rect 151800 22400 151900 22500
rect 151800 22500 151900 22600
rect 151800 22600 151900 22700
rect 151800 22700 151900 22800
rect 151800 22800 151900 22900
rect 151800 22900 151900 23000
rect 151800 23000 151900 23100
rect 151800 23100 151900 23200
rect 151800 23200 151900 23300
rect 151800 23300 151900 23400
rect 151800 23400 151900 23500
rect 151800 23500 151900 23600
rect 151800 23600 151900 23700
rect 151800 23700 151900 23800
rect 151800 23800 151900 23900
rect 151800 23900 151900 24000
rect 151800 24000 151900 24100
rect 151800 24100 151900 24200
rect 151800 24200 151900 24300
rect 151800 24300 151900 24400
rect 151800 24400 151900 24500
rect 151800 24500 151900 24600
rect 151800 24600 151900 24700
rect 151800 24700 151900 24800
rect 151800 24800 151900 24900
rect 151800 24900 151900 25000
rect 151800 25000 151900 25100
rect 151800 25100 151900 25200
rect 151800 25200 151900 25300
rect 151800 25300 151900 25400
rect 151800 25400 151900 25500
rect 151800 25500 151900 25600
rect 151800 25600 151900 25700
rect 151800 25700 151900 25800
rect 151800 25800 151900 25900
rect 151800 25900 151900 26000
rect 151800 26000 151900 26100
rect 151800 26100 151900 26200
rect 151800 26200 151900 26300
rect 151800 26300 151900 26400
rect 151800 26400 151900 26500
rect 151800 26500 151900 26600
rect 151800 26600 151900 26700
rect 151800 26700 151900 26800
rect 151800 26800 151900 26900
rect 151800 26900 151900 27000
rect 151800 27000 151900 27100
rect 151800 27100 151900 27200
rect 151800 27200 151900 27300
rect 151800 27300 151900 27400
rect 151800 27400 151900 27500
rect 151800 27500 151900 27600
rect 151800 27600 151900 27700
rect 151800 27700 151900 27800
rect 151800 27800 151900 27900
rect 151800 27900 151900 28000
rect 151800 28000 151900 28100
rect 151800 28100 151900 28200
rect 151800 28200 151900 28300
rect 151800 28300 151900 28400
rect 151800 28400 151900 28500
rect 151800 28500 151900 28600
rect 151800 28600 151900 28700
rect 151800 28700 151900 28800
rect 151800 28800 151900 28900
rect 151800 28900 151900 29000
rect 151800 30400 151900 30500
rect 151800 30500 151900 30600
rect 151800 30600 151900 30700
rect 151800 30700 151900 30800
rect 151800 30800 151900 30900
rect 151800 30900 151900 31000
rect 151800 31000 151900 31100
rect 151800 31100 151900 31200
rect 151800 31200 151900 31300
rect 151800 31300 151900 31400
rect 151800 31400 151900 31500
rect 151800 31500 151900 31600
rect 151800 31600 151900 31700
rect 151800 31700 151900 31800
rect 151800 31800 151900 31900
rect 151800 31900 151900 32000
rect 151800 32000 151900 32100
rect 151800 32100 151900 32200
rect 151800 32200 151900 32300
rect 151800 32300 151900 32400
rect 151800 32400 151900 32500
rect 151800 32500 151900 32600
rect 151800 32600 151900 32700
rect 151800 32700 151900 32800
rect 151800 32800 151900 32900
rect 151800 32900 151900 33000
rect 151800 33000 151900 33100
rect 151800 33100 151900 33200
rect 151800 33200 151900 33300
rect 151800 33300 151900 33400
rect 151800 33400 151900 33500
rect 151800 33500 151900 33600
rect 151800 33600 151900 33700
rect 151800 33700 151900 33800
rect 151800 33800 151900 33900
rect 151800 33900 151900 34000
rect 151800 34000 151900 34100
rect 151800 34100 151900 34200
rect 151800 34200 151900 34300
rect 151800 34300 151900 34400
rect 151800 34400 151900 34500
rect 151800 34500 151900 34600
rect 151800 34600 151900 34700
rect 151800 34700 151900 34800
rect 151800 34800 151900 34900
rect 151800 34900 151900 35000
rect 151800 35000 151900 35100
rect 151800 35100 151900 35200
rect 151800 35200 151900 35300
rect 151800 35300 151900 35400
rect 151800 35400 151900 35500
rect 151800 35500 151900 35600
rect 151800 35600 151900 35700
rect 151800 35700 151900 35800
rect 151800 35800 151900 35900
rect 151800 35900 151900 36000
rect 151800 36000 151900 36100
rect 151800 36100 151900 36200
rect 151800 36200 151900 36300
rect 151800 36300 151900 36400
rect 151800 36400 151900 36500
rect 151800 36500 151900 36600
rect 151800 36600 151900 36700
rect 151800 36700 151900 36800
rect 151800 36800 151900 36900
rect 151800 36900 151900 37000
rect 151800 37000 151900 37100
rect 151800 37100 151900 37200
rect 151800 37200 151900 37300
rect 151800 37300 151900 37400
rect 151800 37400 151900 37500
rect 151800 37500 151900 37600
rect 151800 37600 151900 37700
rect 151800 37700 151900 37800
rect 151800 37800 151900 37900
rect 151800 37900 151900 38000
rect 151800 38000 151900 38100
rect 151800 38100 151900 38200
rect 151800 38200 151900 38300
rect 151900 21200 152000 21300
rect 151900 21300 152000 21400
rect 151900 21400 152000 21500
rect 151900 21500 152000 21600
rect 151900 21600 152000 21700
rect 151900 21700 152000 21800
rect 151900 21800 152000 21900
rect 151900 21900 152000 22000
rect 151900 22000 152000 22100
rect 151900 22100 152000 22200
rect 151900 22200 152000 22300
rect 151900 22300 152000 22400
rect 151900 22400 152000 22500
rect 151900 22500 152000 22600
rect 151900 22600 152000 22700
rect 151900 22700 152000 22800
rect 151900 22800 152000 22900
rect 151900 22900 152000 23000
rect 151900 23000 152000 23100
rect 151900 23100 152000 23200
rect 151900 23200 152000 23300
rect 151900 23300 152000 23400
rect 151900 23400 152000 23500
rect 151900 23500 152000 23600
rect 151900 23600 152000 23700
rect 151900 23700 152000 23800
rect 151900 23800 152000 23900
rect 151900 23900 152000 24000
rect 151900 24000 152000 24100
rect 151900 24100 152000 24200
rect 151900 24200 152000 24300
rect 151900 24300 152000 24400
rect 151900 24400 152000 24500
rect 151900 24500 152000 24600
rect 151900 24600 152000 24700
rect 151900 24700 152000 24800
rect 151900 24800 152000 24900
rect 151900 24900 152000 25000
rect 151900 25000 152000 25100
rect 151900 25100 152000 25200
rect 151900 25200 152000 25300
rect 151900 25300 152000 25400
rect 151900 25400 152000 25500
rect 151900 25500 152000 25600
rect 151900 25600 152000 25700
rect 151900 25700 152000 25800
rect 151900 25800 152000 25900
rect 151900 25900 152000 26000
rect 151900 26000 152000 26100
rect 151900 26100 152000 26200
rect 151900 26200 152000 26300
rect 151900 26300 152000 26400
rect 151900 26400 152000 26500
rect 151900 26500 152000 26600
rect 151900 26600 152000 26700
rect 151900 26700 152000 26800
rect 151900 26800 152000 26900
rect 151900 26900 152000 27000
rect 151900 27000 152000 27100
rect 151900 27100 152000 27200
rect 151900 27200 152000 27300
rect 151900 27300 152000 27400
rect 151900 27400 152000 27500
rect 151900 27500 152000 27600
rect 151900 27600 152000 27700
rect 151900 27700 152000 27800
rect 151900 27800 152000 27900
rect 151900 27900 152000 28000
rect 151900 28000 152000 28100
rect 151900 28100 152000 28200
rect 151900 28200 152000 28300
rect 151900 28300 152000 28400
rect 151900 28400 152000 28500
rect 151900 28500 152000 28600
rect 151900 28600 152000 28700
rect 151900 28700 152000 28800
rect 151900 28800 152000 28900
rect 151900 28900 152000 29000
rect 151900 30400 152000 30500
rect 151900 30500 152000 30600
rect 151900 30600 152000 30700
rect 151900 30700 152000 30800
rect 151900 30800 152000 30900
rect 151900 30900 152000 31000
rect 151900 31000 152000 31100
rect 151900 31100 152000 31200
rect 151900 31200 152000 31300
rect 151900 31300 152000 31400
rect 151900 31400 152000 31500
rect 151900 31500 152000 31600
rect 151900 31600 152000 31700
rect 151900 31700 152000 31800
rect 151900 31800 152000 31900
rect 151900 31900 152000 32000
rect 151900 32000 152000 32100
rect 151900 32100 152000 32200
rect 151900 32200 152000 32300
rect 151900 32300 152000 32400
rect 151900 32400 152000 32500
rect 151900 32500 152000 32600
rect 151900 32600 152000 32700
rect 151900 32700 152000 32800
rect 151900 32800 152000 32900
rect 151900 32900 152000 33000
rect 151900 33000 152000 33100
rect 151900 33100 152000 33200
rect 151900 33200 152000 33300
rect 151900 33300 152000 33400
rect 151900 33400 152000 33500
rect 151900 33500 152000 33600
rect 151900 33600 152000 33700
rect 151900 33700 152000 33800
rect 151900 33800 152000 33900
rect 151900 33900 152000 34000
rect 151900 34000 152000 34100
rect 151900 34100 152000 34200
rect 151900 34200 152000 34300
rect 151900 34300 152000 34400
rect 151900 34400 152000 34500
rect 151900 34500 152000 34600
rect 151900 34600 152000 34700
rect 151900 34700 152000 34800
rect 151900 34800 152000 34900
rect 151900 34900 152000 35000
rect 151900 35000 152000 35100
rect 151900 35100 152000 35200
rect 151900 35200 152000 35300
rect 151900 35300 152000 35400
rect 151900 35400 152000 35500
rect 151900 35500 152000 35600
rect 151900 35600 152000 35700
rect 151900 35700 152000 35800
rect 151900 35800 152000 35900
rect 151900 35900 152000 36000
rect 151900 36000 152000 36100
rect 151900 36100 152000 36200
rect 151900 36200 152000 36300
rect 151900 36300 152000 36400
rect 151900 36400 152000 36500
rect 151900 36500 152000 36600
rect 151900 36600 152000 36700
rect 151900 36700 152000 36800
rect 151900 36800 152000 36900
rect 151900 36900 152000 37000
rect 151900 37000 152000 37100
rect 151900 37100 152000 37200
rect 151900 37200 152000 37300
rect 151900 37300 152000 37400
rect 151900 37400 152000 37500
rect 151900 37500 152000 37600
rect 151900 37600 152000 37700
rect 151900 37700 152000 37800
rect 151900 37800 152000 37900
rect 151900 37900 152000 38000
rect 151900 38000 152000 38100
rect 151900 38100 152000 38200
rect 151900 38200 152000 38300
rect 152000 21300 152100 21400
rect 152000 21400 152100 21500
rect 152000 21500 152100 21600
rect 152000 21600 152100 21700
rect 152000 21700 152100 21800
rect 152000 21800 152100 21900
rect 152000 21900 152100 22000
rect 152000 22000 152100 22100
rect 152000 22100 152100 22200
rect 152000 22200 152100 22300
rect 152000 22300 152100 22400
rect 152000 22400 152100 22500
rect 152000 22500 152100 22600
rect 152000 22600 152100 22700
rect 152000 22700 152100 22800
rect 152000 22800 152100 22900
rect 152000 22900 152100 23000
rect 152000 23000 152100 23100
rect 152000 23100 152100 23200
rect 152000 23200 152100 23300
rect 152000 23300 152100 23400
rect 152000 23400 152100 23500
rect 152000 23500 152100 23600
rect 152000 23600 152100 23700
rect 152000 23700 152100 23800
rect 152000 23800 152100 23900
rect 152000 23900 152100 24000
rect 152000 24000 152100 24100
rect 152000 24100 152100 24200
rect 152000 24200 152100 24300
rect 152000 24300 152100 24400
rect 152000 24400 152100 24500
rect 152000 24500 152100 24600
rect 152000 24600 152100 24700
rect 152000 24700 152100 24800
rect 152000 24800 152100 24900
rect 152000 24900 152100 25000
rect 152000 25000 152100 25100
rect 152000 25100 152100 25200
rect 152000 25200 152100 25300
rect 152000 25300 152100 25400
rect 152000 25400 152100 25500
rect 152000 25500 152100 25600
rect 152000 25600 152100 25700
rect 152000 25700 152100 25800
rect 152000 25800 152100 25900
rect 152000 25900 152100 26000
rect 152000 26000 152100 26100
rect 152000 26100 152100 26200
rect 152000 26200 152100 26300
rect 152000 26300 152100 26400
rect 152000 26400 152100 26500
rect 152000 26500 152100 26600
rect 152000 26600 152100 26700
rect 152000 26700 152100 26800
rect 152000 26800 152100 26900
rect 152000 26900 152100 27000
rect 152000 27000 152100 27100
rect 152000 27100 152100 27200
rect 152000 27200 152100 27300
rect 152000 27300 152100 27400
rect 152000 27400 152100 27500
rect 152000 27500 152100 27600
rect 152000 27600 152100 27700
rect 152000 27700 152100 27800
rect 152000 27800 152100 27900
rect 152000 27900 152100 28000
rect 152000 28000 152100 28100
rect 152000 28100 152100 28200
rect 152000 28200 152100 28300
rect 152000 28300 152100 28400
rect 152000 28400 152100 28500
rect 152000 28500 152100 28600
rect 152000 28600 152100 28700
rect 152000 28700 152100 28800
rect 152000 28800 152100 28900
rect 152000 28900 152100 29000
rect 152000 30500 152100 30600
rect 152000 30600 152100 30700
rect 152000 30700 152100 30800
rect 152000 30800 152100 30900
rect 152000 30900 152100 31000
rect 152000 31000 152100 31100
rect 152000 31100 152100 31200
rect 152000 31200 152100 31300
rect 152000 31300 152100 31400
rect 152000 31400 152100 31500
rect 152000 31500 152100 31600
rect 152000 31600 152100 31700
rect 152000 31700 152100 31800
rect 152000 31800 152100 31900
rect 152000 31900 152100 32000
rect 152000 32000 152100 32100
rect 152000 32100 152100 32200
rect 152000 32200 152100 32300
rect 152000 32300 152100 32400
rect 152000 32400 152100 32500
rect 152000 32500 152100 32600
rect 152000 32600 152100 32700
rect 152000 32700 152100 32800
rect 152000 32800 152100 32900
rect 152000 32900 152100 33000
rect 152000 33000 152100 33100
rect 152000 33100 152100 33200
rect 152000 33200 152100 33300
rect 152000 33300 152100 33400
rect 152000 33400 152100 33500
rect 152000 33500 152100 33600
rect 152000 33600 152100 33700
rect 152000 33700 152100 33800
rect 152000 33800 152100 33900
rect 152000 33900 152100 34000
rect 152000 34000 152100 34100
rect 152000 34100 152100 34200
rect 152000 34200 152100 34300
rect 152000 34300 152100 34400
rect 152000 34400 152100 34500
rect 152000 34500 152100 34600
rect 152000 34600 152100 34700
rect 152000 34700 152100 34800
rect 152000 34800 152100 34900
rect 152000 34900 152100 35000
rect 152000 35000 152100 35100
rect 152000 35100 152100 35200
rect 152000 35200 152100 35300
rect 152000 35300 152100 35400
rect 152000 35400 152100 35500
rect 152000 35500 152100 35600
rect 152000 35600 152100 35700
rect 152000 35700 152100 35800
rect 152000 35800 152100 35900
rect 152000 35900 152100 36000
rect 152000 36000 152100 36100
rect 152000 36100 152100 36200
rect 152000 36200 152100 36300
rect 152000 36300 152100 36400
rect 152000 36400 152100 36500
rect 152000 36500 152100 36600
rect 152000 36600 152100 36700
rect 152000 36700 152100 36800
rect 152000 36800 152100 36900
rect 152000 36900 152100 37000
rect 152000 37000 152100 37100
rect 152000 37100 152100 37200
rect 152000 37200 152100 37300
rect 152000 37300 152100 37400
rect 152000 37400 152100 37500
rect 152000 37500 152100 37600
rect 152000 37600 152100 37700
rect 152000 37700 152100 37800
rect 152000 37800 152100 37900
rect 152000 37900 152100 38000
rect 152000 38000 152100 38100
rect 152000 38100 152100 38200
rect 152100 21400 152200 21500
rect 152100 21500 152200 21600
rect 152100 21600 152200 21700
rect 152100 21700 152200 21800
rect 152100 21800 152200 21900
rect 152100 21900 152200 22000
rect 152100 22000 152200 22100
rect 152100 22100 152200 22200
rect 152100 22200 152200 22300
rect 152100 22300 152200 22400
rect 152100 22400 152200 22500
rect 152100 22500 152200 22600
rect 152100 22600 152200 22700
rect 152100 22700 152200 22800
rect 152100 22800 152200 22900
rect 152100 22900 152200 23000
rect 152100 23000 152200 23100
rect 152100 23100 152200 23200
rect 152100 23200 152200 23300
rect 152100 23300 152200 23400
rect 152100 23400 152200 23500
rect 152100 23500 152200 23600
rect 152100 23600 152200 23700
rect 152100 23700 152200 23800
rect 152100 23800 152200 23900
rect 152100 23900 152200 24000
rect 152100 24000 152200 24100
rect 152100 24100 152200 24200
rect 152100 24200 152200 24300
rect 152100 24300 152200 24400
rect 152100 24400 152200 24500
rect 152100 24500 152200 24600
rect 152100 24600 152200 24700
rect 152100 24700 152200 24800
rect 152100 24800 152200 24900
rect 152100 24900 152200 25000
rect 152100 25000 152200 25100
rect 152100 25100 152200 25200
rect 152100 25200 152200 25300
rect 152100 25300 152200 25400
rect 152100 25400 152200 25500
rect 152100 25500 152200 25600
rect 152100 25600 152200 25700
rect 152100 25700 152200 25800
rect 152100 25800 152200 25900
rect 152100 25900 152200 26000
rect 152100 26000 152200 26100
rect 152100 26100 152200 26200
rect 152100 26200 152200 26300
rect 152100 26300 152200 26400
rect 152100 26400 152200 26500
rect 152100 26500 152200 26600
rect 152100 26600 152200 26700
rect 152100 26700 152200 26800
rect 152100 26800 152200 26900
rect 152100 26900 152200 27000
rect 152100 27000 152200 27100
rect 152100 27100 152200 27200
rect 152100 27200 152200 27300
rect 152100 27300 152200 27400
rect 152100 27400 152200 27500
rect 152100 27500 152200 27600
rect 152100 27600 152200 27700
rect 152100 27700 152200 27800
rect 152100 27800 152200 27900
rect 152100 27900 152200 28000
rect 152100 28000 152200 28100
rect 152100 28100 152200 28200
rect 152100 28200 152200 28300
rect 152100 28300 152200 28400
rect 152100 28400 152200 28500
rect 152100 28500 152200 28600
rect 152100 28600 152200 28700
rect 152100 28700 152200 28800
rect 152100 28800 152200 28900
rect 152100 30500 152200 30600
rect 152100 30600 152200 30700
rect 152100 30700 152200 30800
rect 152100 30800 152200 30900
rect 152100 30900 152200 31000
rect 152100 31000 152200 31100
rect 152100 31100 152200 31200
rect 152100 31200 152200 31300
rect 152100 31300 152200 31400
rect 152100 31400 152200 31500
rect 152100 31500 152200 31600
rect 152100 31600 152200 31700
rect 152100 31700 152200 31800
rect 152100 31800 152200 31900
rect 152100 31900 152200 32000
rect 152100 32000 152200 32100
rect 152100 32100 152200 32200
rect 152100 32200 152200 32300
rect 152100 32300 152200 32400
rect 152100 32400 152200 32500
rect 152100 32500 152200 32600
rect 152100 32600 152200 32700
rect 152100 32700 152200 32800
rect 152100 32800 152200 32900
rect 152100 32900 152200 33000
rect 152100 33000 152200 33100
rect 152100 33100 152200 33200
rect 152100 33200 152200 33300
rect 152100 33300 152200 33400
rect 152100 33400 152200 33500
rect 152100 33500 152200 33600
rect 152100 33600 152200 33700
rect 152100 33700 152200 33800
rect 152100 33800 152200 33900
rect 152100 33900 152200 34000
rect 152100 34000 152200 34100
rect 152100 34100 152200 34200
rect 152100 34200 152200 34300
rect 152100 34300 152200 34400
rect 152100 34400 152200 34500
rect 152100 34500 152200 34600
rect 152100 34600 152200 34700
rect 152100 34700 152200 34800
rect 152100 34800 152200 34900
rect 152100 34900 152200 35000
rect 152100 35000 152200 35100
rect 152100 35100 152200 35200
rect 152100 35200 152200 35300
rect 152100 35300 152200 35400
rect 152100 35400 152200 35500
rect 152100 35500 152200 35600
rect 152100 35600 152200 35700
rect 152100 35700 152200 35800
rect 152100 35800 152200 35900
rect 152100 35900 152200 36000
rect 152100 36000 152200 36100
rect 152100 36100 152200 36200
rect 152100 36200 152200 36300
rect 152100 36300 152200 36400
rect 152100 36400 152200 36500
rect 152100 36500 152200 36600
rect 152100 36600 152200 36700
rect 152100 36700 152200 36800
rect 152100 36800 152200 36900
rect 152100 36900 152200 37000
rect 152100 37000 152200 37100
rect 152100 37100 152200 37200
rect 152100 37200 152200 37300
rect 152100 37300 152200 37400
rect 152100 37400 152200 37500
rect 152100 37500 152200 37600
rect 152100 37600 152200 37700
rect 152100 37700 152200 37800
rect 152100 37800 152200 37900
rect 152100 37900 152200 38000
rect 152100 38000 152200 38100
rect 152100 38100 152200 38200
rect 152200 21600 152300 21700
rect 152200 21700 152300 21800
rect 152200 21800 152300 21900
rect 152200 21900 152300 22000
rect 152200 22000 152300 22100
rect 152200 22100 152300 22200
rect 152200 22200 152300 22300
rect 152200 22300 152300 22400
rect 152200 22400 152300 22500
rect 152200 22500 152300 22600
rect 152200 22600 152300 22700
rect 152200 22700 152300 22800
rect 152200 22800 152300 22900
rect 152200 22900 152300 23000
rect 152200 23000 152300 23100
rect 152200 23100 152300 23200
rect 152200 23200 152300 23300
rect 152200 23300 152300 23400
rect 152200 23400 152300 23500
rect 152200 23500 152300 23600
rect 152200 23600 152300 23700
rect 152200 23700 152300 23800
rect 152200 23800 152300 23900
rect 152200 23900 152300 24000
rect 152200 24000 152300 24100
rect 152200 24100 152300 24200
rect 152200 24200 152300 24300
rect 152200 24300 152300 24400
rect 152200 24400 152300 24500
rect 152200 24500 152300 24600
rect 152200 24600 152300 24700
rect 152200 24700 152300 24800
rect 152200 24800 152300 24900
rect 152200 24900 152300 25000
rect 152200 25000 152300 25100
rect 152200 25100 152300 25200
rect 152200 25200 152300 25300
rect 152200 25300 152300 25400
rect 152200 25400 152300 25500
rect 152200 25500 152300 25600
rect 152200 25600 152300 25700
rect 152200 25700 152300 25800
rect 152200 25800 152300 25900
rect 152200 25900 152300 26000
rect 152200 26000 152300 26100
rect 152200 26100 152300 26200
rect 152200 26200 152300 26300
rect 152200 26300 152300 26400
rect 152200 26400 152300 26500
rect 152200 26500 152300 26600
rect 152200 26600 152300 26700
rect 152200 26700 152300 26800
rect 152200 26800 152300 26900
rect 152200 26900 152300 27000
rect 152200 27000 152300 27100
rect 152200 27100 152300 27200
rect 152200 27200 152300 27300
rect 152200 27300 152300 27400
rect 152200 27400 152300 27500
rect 152200 27500 152300 27600
rect 152200 27600 152300 27700
rect 152200 27700 152300 27800
rect 152200 27800 152300 27900
rect 152200 27900 152300 28000
rect 152200 28000 152300 28100
rect 152200 28100 152300 28200
rect 152200 28200 152300 28300
rect 152200 28300 152300 28400
rect 152200 28400 152300 28500
rect 152200 28500 152300 28600
rect 152200 28600 152300 28700
rect 152200 28700 152300 28800
rect 152200 28800 152300 28900
rect 152200 28900 152300 29000
rect 152200 30600 152300 30700
rect 152200 30700 152300 30800
rect 152200 30800 152300 30900
rect 152200 30900 152300 31000
rect 152200 31000 152300 31100
rect 152200 31100 152300 31200
rect 152200 31200 152300 31300
rect 152200 31300 152300 31400
rect 152200 31400 152300 31500
rect 152200 31500 152300 31600
rect 152200 31600 152300 31700
rect 152200 31700 152300 31800
rect 152200 31800 152300 31900
rect 152200 31900 152300 32000
rect 152200 32000 152300 32100
rect 152200 32100 152300 32200
rect 152200 32200 152300 32300
rect 152200 32300 152300 32400
rect 152200 32400 152300 32500
rect 152200 32500 152300 32600
rect 152200 32600 152300 32700
rect 152200 32700 152300 32800
rect 152200 32800 152300 32900
rect 152200 32900 152300 33000
rect 152200 33000 152300 33100
rect 152200 33100 152300 33200
rect 152200 33200 152300 33300
rect 152200 33300 152300 33400
rect 152200 33400 152300 33500
rect 152200 33500 152300 33600
rect 152200 33600 152300 33700
rect 152200 33700 152300 33800
rect 152200 33800 152300 33900
rect 152200 33900 152300 34000
rect 152200 34000 152300 34100
rect 152200 34100 152300 34200
rect 152200 34200 152300 34300
rect 152200 34300 152300 34400
rect 152200 34400 152300 34500
rect 152200 34500 152300 34600
rect 152200 34600 152300 34700
rect 152200 34700 152300 34800
rect 152200 34800 152300 34900
rect 152200 34900 152300 35000
rect 152200 35000 152300 35100
rect 152200 35100 152300 35200
rect 152200 35200 152300 35300
rect 152200 35300 152300 35400
rect 152200 35400 152300 35500
rect 152200 35500 152300 35600
rect 152200 35600 152300 35700
rect 152200 35700 152300 35800
rect 152200 35800 152300 35900
rect 152200 35900 152300 36000
rect 152200 36000 152300 36100
rect 152200 36100 152300 36200
rect 152200 36200 152300 36300
rect 152200 36300 152300 36400
rect 152200 36400 152300 36500
rect 152200 36500 152300 36600
rect 152200 36600 152300 36700
rect 152200 36700 152300 36800
rect 152200 36800 152300 36900
rect 152200 36900 152300 37000
rect 152200 37000 152300 37100
rect 152200 37100 152300 37200
rect 152200 37200 152300 37300
rect 152200 37300 152300 37400
rect 152200 37400 152300 37500
rect 152200 37500 152300 37600
rect 152200 37600 152300 37700
rect 152200 37700 152300 37800
rect 152200 37800 152300 37900
rect 152200 37900 152300 38000
rect 152200 38000 152300 38100
rect 152300 21900 152400 22000
rect 152300 22000 152400 22100
rect 152300 22100 152400 22200
rect 152300 22200 152400 22300
rect 152300 22300 152400 22400
rect 152300 22400 152400 22500
rect 152300 22500 152400 22600
rect 152300 22600 152400 22700
rect 152300 22700 152400 22800
rect 152300 22800 152400 22900
rect 152300 22900 152400 23000
rect 152300 23000 152400 23100
rect 152300 23100 152400 23200
rect 152300 23200 152400 23300
rect 152300 23300 152400 23400
rect 152300 23400 152400 23500
rect 152300 23500 152400 23600
rect 152300 23600 152400 23700
rect 152300 23700 152400 23800
rect 152300 23800 152400 23900
rect 152300 23900 152400 24000
rect 152300 24000 152400 24100
rect 152300 24100 152400 24200
rect 152300 24200 152400 24300
rect 152300 24300 152400 24400
rect 152300 24400 152400 24500
rect 152300 24500 152400 24600
rect 152300 24600 152400 24700
rect 152300 24700 152400 24800
rect 152300 24800 152400 24900
rect 152300 24900 152400 25000
rect 152300 25000 152400 25100
rect 152300 25100 152400 25200
rect 152300 25200 152400 25300
rect 152300 25300 152400 25400
rect 152300 25400 152400 25500
rect 152300 25500 152400 25600
rect 152300 25600 152400 25700
rect 152300 25700 152400 25800
rect 152300 25800 152400 25900
rect 152300 25900 152400 26000
rect 152300 26000 152400 26100
rect 152300 26100 152400 26200
rect 152300 26200 152400 26300
rect 152300 26300 152400 26400
rect 152300 26400 152400 26500
rect 152300 26500 152400 26600
rect 152300 26600 152400 26700
rect 152300 26700 152400 26800
rect 152300 26800 152400 26900
rect 152300 26900 152400 27000
rect 152300 27000 152400 27100
rect 152300 27100 152400 27200
rect 152300 27200 152400 27300
rect 152300 27300 152400 27400
rect 152300 27400 152400 27500
rect 152300 27500 152400 27600
rect 152300 27600 152400 27700
rect 152300 27700 152400 27800
rect 152300 27800 152400 27900
rect 152300 27900 152400 28000
rect 152300 28000 152400 28100
rect 152300 28100 152400 28200
rect 152300 28200 152400 28300
rect 152300 28300 152400 28400
rect 152300 28400 152400 28500
rect 152300 28500 152400 28600
rect 152300 28600 152400 28700
rect 152300 28700 152400 28800
rect 152300 28800 152400 28900
rect 152300 28900 152400 29000
rect 152300 30600 152400 30700
rect 152300 30700 152400 30800
rect 152300 30800 152400 30900
rect 152300 30900 152400 31000
rect 152300 31000 152400 31100
rect 152300 31100 152400 31200
rect 152300 31200 152400 31300
rect 152300 31300 152400 31400
rect 152300 31400 152400 31500
rect 152300 31500 152400 31600
rect 152300 31600 152400 31700
rect 152300 31700 152400 31800
rect 152300 31800 152400 31900
rect 152300 31900 152400 32000
rect 152300 32000 152400 32100
rect 152300 32100 152400 32200
rect 152300 32200 152400 32300
rect 152300 32300 152400 32400
rect 152300 32400 152400 32500
rect 152300 32500 152400 32600
rect 152300 32600 152400 32700
rect 152300 32700 152400 32800
rect 152300 32800 152400 32900
rect 152300 32900 152400 33000
rect 152300 33000 152400 33100
rect 152300 33100 152400 33200
rect 152300 33200 152400 33300
rect 152300 33300 152400 33400
rect 152300 33400 152400 33500
rect 152300 33500 152400 33600
rect 152300 33600 152400 33700
rect 152300 33700 152400 33800
rect 152300 33800 152400 33900
rect 152300 33900 152400 34000
rect 152300 34000 152400 34100
rect 152300 34100 152400 34200
rect 152300 34200 152400 34300
rect 152300 34300 152400 34400
rect 152300 34400 152400 34500
rect 152300 34500 152400 34600
rect 152300 34600 152400 34700
rect 152300 34700 152400 34800
rect 152300 34800 152400 34900
rect 152300 34900 152400 35000
rect 152300 35000 152400 35100
rect 152300 35100 152400 35200
rect 152300 35200 152400 35300
rect 152300 35300 152400 35400
rect 152300 35400 152400 35500
rect 152300 35500 152400 35600
rect 152300 35600 152400 35700
rect 152300 35700 152400 35800
rect 152300 35800 152400 35900
rect 152300 35900 152400 36000
rect 152300 36000 152400 36100
rect 152300 36100 152400 36200
rect 152300 36200 152400 36300
rect 152300 36300 152400 36400
rect 152300 36400 152400 36500
rect 152300 36500 152400 36600
rect 152300 36600 152400 36700
rect 152300 36700 152400 36800
rect 152300 36800 152400 36900
rect 152300 36900 152400 37000
rect 152300 37000 152400 37100
rect 152300 37100 152400 37200
rect 152300 37200 152400 37300
rect 152300 37300 152400 37400
rect 152300 37400 152400 37500
rect 152300 37500 152400 37600
rect 152300 37600 152400 37700
rect 152300 37700 152400 37800
rect 152300 37800 152400 37900
rect 152300 37900 152400 38000
rect 152400 27300 152500 27400
rect 152400 27400 152500 27500
rect 152400 27500 152500 27600
rect 152400 27600 152500 27700
rect 152400 27700 152500 27800
rect 152400 27800 152500 27900
rect 152400 27900 152500 28000
rect 152400 28000 152500 28100
rect 152400 28100 152500 28200
rect 152400 28200 152500 28300
rect 152400 28300 152500 28400
rect 152400 28400 152500 28500
rect 152400 28500 152500 28600
rect 152400 28600 152500 28700
rect 152400 28700 152500 28800
rect 152400 28800 152500 28900
rect 152400 28900 152500 29000
rect 152400 30600 152500 30700
rect 152400 30700 152500 30800
rect 152400 30800 152500 30900
rect 152400 30900 152500 31000
rect 152400 31000 152500 31100
rect 152400 31100 152500 31200
rect 152400 31200 152500 31300
rect 152400 31300 152500 31400
rect 152400 31400 152500 31500
rect 152400 31500 152500 31600
rect 152400 31600 152500 31700
rect 152400 31700 152500 31800
rect 152400 31800 152500 31900
rect 152400 31900 152500 32000
rect 152400 32000 152500 32100
rect 152400 32100 152500 32200
rect 152400 33700 152500 33800
rect 152400 33900 152500 34000
rect 152400 34000 152500 34100
rect 152400 34100 152500 34200
rect 152400 34200 152500 34300
rect 152400 34300 152500 34400
rect 152400 34400 152500 34500
rect 152400 34500 152500 34600
rect 152400 34600 152500 34700
rect 152400 34700 152500 34800
rect 152400 34800 152500 34900
rect 152400 34900 152500 35000
rect 152400 35000 152500 35100
rect 152400 35100 152500 35200
rect 152400 35200 152500 35300
rect 152400 35300 152500 35400
rect 152400 35400 152500 35500
rect 152400 35500 152500 35600
rect 152400 35600 152500 35700
rect 152400 35700 152500 35800
rect 152400 35800 152500 35900
rect 152400 35900 152500 36000
rect 152400 36000 152500 36100
rect 152400 36100 152500 36200
rect 152400 36200 152500 36300
rect 152400 36300 152500 36400
rect 152400 36400 152500 36500
rect 152400 36500 152500 36600
rect 152400 36600 152500 36700
rect 152400 36700 152500 36800
rect 152400 36800 152500 36900
rect 152400 36900 152500 37000
rect 152400 37000 152500 37100
rect 152400 37100 152500 37200
rect 152400 37200 152500 37300
rect 152400 37300 152500 37400
rect 152400 37400 152500 37500
rect 152400 37500 152500 37600
rect 152400 37600 152500 37700
rect 152400 37700 152500 37800
rect 152500 27300 152600 27400
rect 152500 27400 152600 27500
rect 152500 27500 152600 27600
rect 152500 27600 152600 27700
rect 152500 27700 152600 27800
rect 152500 27800 152600 27900
rect 152500 27900 152600 28000
rect 152500 28000 152600 28100
rect 152500 28100 152600 28200
rect 152500 28200 152600 28300
rect 152500 28300 152600 28400
rect 152500 28400 152600 28500
rect 152500 28500 152600 28600
rect 152500 28600 152600 28700
rect 152500 28700 152600 28800
rect 152500 28800 152600 28900
rect 152500 28900 152600 29000
rect 152500 29000 152600 29100
rect 152500 30600 152600 30700
rect 152500 30700 152600 30800
rect 152500 30800 152600 30900
rect 152500 30900 152600 31000
rect 152500 31000 152600 31100
rect 152500 31100 152600 31200
rect 152500 31200 152600 31300
rect 152500 31300 152600 31400
rect 152500 31400 152600 31500
rect 152500 31500 152600 31600
rect 152500 31600 152600 31700
rect 152500 31700 152600 31800
rect 152500 31800 152600 31900
rect 152500 31900 152600 32000
rect 152500 32000 152600 32100
rect 152500 32100 152600 32200
rect 152500 35700 152600 35800
rect 152500 35900 152600 36000
rect 152500 36000 152600 36100
rect 152500 36100 152600 36200
rect 152500 36200 152600 36300
rect 152500 36300 152600 36400
rect 152500 36400 152600 36500
rect 152500 36500 152600 36600
rect 152500 36600 152600 36700
rect 152500 36700 152600 36800
rect 152500 36800 152600 36900
rect 152500 36900 152600 37000
rect 152500 37000 152600 37100
rect 152500 37100 152600 37200
rect 152500 37200 152600 37300
rect 152500 37300 152600 37400
rect 152500 37400 152600 37500
rect 152500 37500 152600 37600
rect 152600 27300 152700 27400
rect 152600 27400 152700 27500
rect 152600 27500 152700 27600
rect 152600 27600 152700 27700
rect 152600 27700 152700 27800
rect 152600 27800 152700 27900
rect 152600 27900 152700 28000
rect 152600 28000 152700 28100
rect 152600 28100 152700 28200
rect 152600 28200 152700 28300
rect 152600 28300 152700 28400
rect 152600 28400 152700 28500
rect 152600 28500 152700 28600
rect 152600 28600 152700 28700
rect 152600 28700 152700 28800
rect 152600 28800 152700 28900
rect 152600 28900 152700 29000
rect 152600 29000 152700 29100
rect 152600 30500 152700 30600
rect 152600 30600 152700 30700
rect 152600 30700 152700 30800
rect 152600 30800 152700 30900
rect 152600 30900 152700 31000
rect 152600 31000 152700 31100
rect 152600 31100 152700 31200
rect 152600 31200 152700 31300
rect 152600 31300 152700 31400
rect 152600 31400 152700 31500
rect 152600 31500 152700 31600
rect 152600 31600 152700 31700
rect 152600 31700 152700 31800
rect 152600 31800 152700 31900
rect 152600 31900 152700 32000
rect 152600 32000 152700 32100
rect 152700 27300 152800 27400
rect 152700 27400 152800 27500
rect 152700 27500 152800 27600
rect 152700 27600 152800 27700
rect 152700 27700 152800 27800
rect 152700 27800 152800 27900
rect 152700 27900 152800 28000
rect 152700 28000 152800 28100
rect 152700 28100 152800 28200
rect 152700 28200 152800 28300
rect 152700 28300 152800 28400
rect 152700 28400 152800 28500
rect 152700 28500 152800 28600
rect 152700 28600 152800 28700
rect 152700 28700 152800 28800
rect 152700 28800 152800 28900
rect 152700 28900 152800 29000
rect 152700 29000 152800 29100
rect 152700 29100 152800 29200
rect 152700 30500 152800 30600
rect 152700 30600 152800 30700
rect 152700 30700 152800 30800
rect 152700 30800 152800 30900
rect 152700 30900 152800 31000
rect 152700 31000 152800 31100
rect 152700 31100 152800 31200
rect 152700 31200 152800 31300
rect 152700 31300 152800 31400
rect 152700 31400 152800 31500
rect 152700 31500 152800 31600
rect 152700 31600 152800 31700
rect 152700 31700 152800 31800
rect 152700 31800 152800 31900
rect 152700 31900 152800 32000
rect 152700 32000 152800 32100
rect 152800 27300 152900 27400
rect 152800 27400 152900 27500
rect 152800 27500 152900 27600
rect 152800 27600 152900 27700
rect 152800 27700 152900 27800
rect 152800 27800 152900 27900
rect 152800 27900 152900 28000
rect 152800 28000 152900 28100
rect 152800 28100 152900 28200
rect 152800 28200 152900 28300
rect 152800 28300 152900 28400
rect 152800 28400 152900 28500
rect 152800 28500 152900 28600
rect 152800 28600 152900 28700
rect 152800 28700 152900 28800
rect 152800 28800 152900 28900
rect 152800 28900 152900 29000
rect 152800 29000 152900 29100
rect 152800 29100 152900 29200
rect 152800 29200 152900 29300
rect 152800 30400 152900 30500
rect 152800 30500 152900 30600
rect 152800 30600 152900 30700
rect 152800 30700 152900 30800
rect 152800 30800 152900 30900
rect 152800 30900 152900 31000
rect 152800 31000 152900 31100
rect 152800 31100 152900 31200
rect 152800 31200 152900 31300
rect 152800 31300 152900 31400
rect 152800 31400 152900 31500
rect 152800 31500 152900 31600
rect 152800 31600 152900 31700
rect 152800 31700 152900 31800
rect 152800 31800 152900 31900
rect 152800 31900 152900 32000
rect 152800 32000 152900 32100
rect 152900 27200 153000 27300
rect 152900 27300 153000 27400
rect 152900 27400 153000 27500
rect 152900 27500 153000 27600
rect 152900 27600 153000 27700
rect 152900 27700 153000 27800
rect 152900 27800 153000 27900
rect 152900 27900 153000 28000
rect 152900 28000 153000 28100
rect 152900 28100 153000 28200
rect 152900 28200 153000 28300
rect 152900 28300 153000 28400
rect 152900 28400 153000 28500
rect 152900 28500 153000 28600
rect 152900 28600 153000 28700
rect 152900 28700 153000 28800
rect 152900 28800 153000 28900
rect 152900 28900 153000 29000
rect 152900 29000 153000 29100
rect 152900 29100 153000 29200
rect 152900 29200 153000 29300
rect 152900 29300 153000 29400
rect 152900 30300 153000 30400
rect 152900 30400 153000 30500
rect 152900 30500 153000 30600
rect 152900 30600 153000 30700
rect 152900 30700 153000 30800
rect 152900 30800 153000 30900
rect 152900 30900 153000 31000
rect 152900 31000 153000 31100
rect 152900 31100 153000 31200
rect 152900 31200 153000 31300
rect 152900 31300 153000 31400
rect 152900 31400 153000 31500
rect 152900 31500 153000 31600
rect 152900 31600 153000 31700
rect 152900 31700 153000 31800
rect 152900 31800 153000 31900
rect 152900 31900 153000 32000
rect 153000 27100 153100 27200
rect 153000 27200 153100 27300
rect 153000 27300 153100 27400
rect 153000 27400 153100 27500
rect 153000 27500 153100 27600
rect 153000 27600 153100 27700
rect 153000 27700 153100 27800
rect 153000 27800 153100 27900
rect 153000 27900 153100 28000
rect 153000 28000 153100 28100
rect 153000 28100 153100 28200
rect 153000 28200 153100 28300
rect 153000 28300 153100 28400
rect 153000 28400 153100 28500
rect 153000 28500 153100 28600
rect 153000 28600 153100 28700
rect 153000 28700 153100 28800
rect 153000 28800 153100 28900
rect 153000 28900 153100 29000
rect 153000 29000 153100 29100
rect 153000 29100 153100 29200
rect 153000 29200 153100 29300
rect 153000 29300 153100 29400
rect 153000 29400 153100 29500
rect 153000 30200 153100 30300
rect 153000 30300 153100 30400
rect 153000 30400 153100 30500
rect 153000 30500 153100 30600
rect 153000 30600 153100 30700
rect 153000 30700 153100 30800
rect 153000 30800 153100 30900
rect 153000 30900 153100 31000
rect 153000 31000 153100 31100
rect 153000 31100 153100 31200
rect 153000 31200 153100 31300
rect 153000 31300 153100 31400
rect 153000 31400 153100 31500
rect 153000 31500 153100 31600
rect 153000 31600 153100 31700
rect 153000 31700 153100 31800
rect 153000 31800 153100 31900
rect 153000 31900 153100 32000
rect 153100 27000 153200 27100
rect 153100 27100 153200 27200
rect 153100 27200 153200 27300
rect 153100 27300 153200 27400
rect 153100 27400 153200 27500
rect 153100 27500 153200 27600
rect 153100 27600 153200 27700
rect 153100 27700 153200 27800
rect 153100 27800 153200 27900
rect 153100 27900 153200 28000
rect 153100 28000 153200 28100
rect 153100 28100 153200 28200
rect 153100 28200 153200 28300
rect 153100 28300 153200 28400
rect 153100 28400 153200 28500
rect 153100 28500 153200 28600
rect 153100 28600 153200 28700
rect 153100 28700 153200 28800
rect 153100 28800 153200 28900
rect 153100 28900 153200 29000
rect 153100 29000 153200 29100
rect 153100 29100 153200 29200
rect 153100 29200 153200 29300
rect 153100 29300 153200 29400
rect 153100 29400 153200 29500
rect 153100 29500 153200 29600
rect 153100 29600 153200 29700
rect 153100 29700 153200 29800
rect 153100 29800 153200 29900
rect 153100 29900 153200 30000
rect 153100 30000 153200 30100
rect 153100 30100 153200 30200
rect 153100 30200 153200 30300
rect 153100 30300 153200 30400
rect 153100 30400 153200 30500
rect 153100 30500 153200 30600
rect 153100 30600 153200 30700
rect 153100 30700 153200 30800
rect 153100 30800 153200 30900
rect 153100 30900 153200 31000
rect 153100 31000 153200 31100
rect 153100 31100 153200 31200
rect 153100 31200 153200 31300
rect 153100 31300 153200 31400
rect 153100 31400 153200 31500
rect 153100 31500 153200 31600
rect 153100 31600 153200 31700
rect 153100 31700 153200 31800
rect 153100 31800 153200 31900
rect 153100 31900 153200 32000
rect 153200 26900 153300 27000
rect 153200 27000 153300 27100
rect 153200 27100 153300 27200
rect 153200 27200 153300 27300
rect 153200 27300 153300 27400
rect 153200 27400 153300 27500
rect 153200 27500 153300 27600
rect 153200 27600 153300 27700
rect 153200 27700 153300 27800
rect 153200 27800 153300 27900
rect 153200 27900 153300 28000
rect 153200 28000 153300 28100
rect 153200 28100 153300 28200
rect 153200 28200 153300 28300
rect 153200 28300 153300 28400
rect 153200 28400 153300 28500
rect 153200 28500 153300 28600
rect 153200 28600 153300 28700
rect 153200 28700 153300 28800
rect 153200 28800 153300 28900
rect 153200 28900 153300 29000
rect 153200 29000 153300 29100
rect 153200 29100 153300 29200
rect 153200 29200 153300 29300
rect 153200 29300 153300 29400
rect 153200 29400 153300 29500
rect 153200 29500 153300 29600
rect 153200 29600 153300 29700
rect 153200 29700 153300 29800
rect 153200 29800 153300 29900
rect 153200 29900 153300 30000
rect 153200 30000 153300 30100
rect 153200 30100 153300 30200
rect 153200 30200 153300 30300
rect 153200 30300 153300 30400
rect 153200 30400 153300 30500
rect 153200 30500 153300 30600
rect 153200 30600 153300 30700
rect 153200 30700 153300 30800
rect 153200 30800 153300 30900
rect 153200 30900 153300 31000
rect 153200 31000 153300 31100
rect 153200 31100 153300 31200
rect 153200 31200 153300 31300
rect 153200 31300 153300 31400
rect 153200 31400 153300 31500
rect 153200 31500 153300 31600
rect 153200 31600 153300 31700
rect 153200 31700 153300 31800
rect 153200 31800 153300 31900
rect 153300 26800 153400 26900
rect 153300 26900 153400 27000
rect 153300 27000 153400 27100
rect 153300 27100 153400 27200
rect 153300 27200 153400 27300
rect 153300 27300 153400 27400
rect 153300 27400 153400 27500
rect 153300 27500 153400 27600
rect 153300 27600 153400 27700
rect 153300 27700 153400 27800
rect 153300 27800 153400 27900
rect 153300 27900 153400 28000
rect 153300 28000 153400 28100
rect 153300 28100 153400 28200
rect 153300 28200 153400 28300
rect 153300 28300 153400 28400
rect 153300 28400 153400 28500
rect 153300 28500 153400 28600
rect 153300 28600 153400 28700
rect 153300 28700 153400 28800
rect 153300 28800 153400 28900
rect 153300 28900 153400 29000
rect 153300 29000 153400 29100
rect 153300 29100 153400 29200
rect 153300 29200 153400 29300
rect 153300 29300 153400 29400
rect 153300 29400 153400 29500
rect 153300 29500 153400 29600
rect 153300 29600 153400 29700
rect 153300 29700 153400 29800
rect 153300 29800 153400 29900
rect 153300 29900 153400 30000
rect 153300 30000 153400 30100
rect 153300 30100 153400 30200
rect 153300 30200 153400 30300
rect 153300 30300 153400 30400
rect 153300 30400 153400 30500
rect 153300 30500 153400 30600
rect 153300 30600 153400 30700
rect 153300 30700 153400 30800
rect 153300 30800 153400 30900
rect 153300 30900 153400 31000
rect 153300 31000 153400 31100
rect 153300 31100 153400 31200
rect 153300 31200 153400 31300
rect 153300 31300 153400 31400
rect 153300 31400 153400 31500
rect 153300 31500 153400 31600
rect 153300 31600 153400 31700
rect 153300 31700 153400 31800
rect 153300 31800 153400 31900
rect 153400 26700 153500 26800
rect 153400 26800 153500 26900
rect 153400 26900 153500 27000
rect 153400 27000 153500 27100
rect 153400 27100 153500 27200
rect 153400 27200 153500 27300
rect 153400 27300 153500 27400
rect 153400 27400 153500 27500
rect 153400 27500 153500 27600
rect 153400 27600 153500 27700
rect 153400 27700 153500 27800
rect 153400 27800 153500 27900
rect 153400 27900 153500 28000
rect 153400 28000 153500 28100
rect 153400 28100 153500 28200
rect 153400 28200 153500 28300
rect 153400 28300 153500 28400
rect 153400 28400 153500 28500
rect 153400 28500 153500 28600
rect 153400 28600 153500 28700
rect 153400 28700 153500 28800
rect 153400 28800 153500 28900
rect 153400 28900 153500 29000
rect 153400 29000 153500 29100
rect 153400 29100 153500 29200
rect 153400 29200 153500 29300
rect 153400 29300 153500 29400
rect 153400 29400 153500 29500
rect 153400 29500 153500 29600
rect 153400 29600 153500 29700
rect 153400 29700 153500 29800
rect 153400 29800 153500 29900
rect 153400 29900 153500 30000
rect 153400 30000 153500 30100
rect 153400 30100 153500 30200
rect 153400 30200 153500 30300
rect 153400 30300 153500 30400
rect 153400 30400 153500 30500
rect 153400 30500 153500 30600
rect 153400 30600 153500 30700
rect 153400 30700 153500 30800
rect 153400 30800 153500 30900
rect 153400 30900 153500 31000
rect 153400 31000 153500 31100
rect 153400 31100 153500 31200
rect 153400 31200 153500 31300
rect 153400 31300 153500 31400
rect 153400 31400 153500 31500
rect 153400 31500 153500 31600
rect 153400 31600 153500 31700
rect 153400 31700 153500 31800
rect 153400 31800 153500 31900
rect 153400 31900 153500 32000
rect 153500 26600 153600 26700
rect 153500 26700 153600 26800
rect 153500 26800 153600 26900
rect 153500 26900 153600 27000
rect 153500 27000 153600 27100
rect 153500 27100 153600 27200
rect 153500 27200 153600 27300
rect 153500 27300 153600 27400
rect 153500 27400 153600 27500
rect 153500 27500 153600 27600
rect 153500 27600 153600 27700
rect 153500 27700 153600 27800
rect 153500 27800 153600 27900
rect 153500 27900 153600 28000
rect 153500 28000 153600 28100
rect 153500 28100 153600 28200
rect 153500 28200 153600 28300
rect 153500 28300 153600 28400
rect 153500 28400 153600 28500
rect 153500 28500 153600 28600
rect 153500 28600 153600 28700
rect 153500 28700 153600 28800
rect 153500 28800 153600 28900
rect 153500 28900 153600 29000
rect 153500 29000 153600 29100
rect 153500 29100 153600 29200
rect 153500 29200 153600 29300
rect 153500 29300 153600 29400
rect 153500 29400 153600 29500
rect 153500 29500 153600 29600
rect 153500 29600 153600 29700
rect 153500 29700 153600 29800
rect 153500 29800 153600 29900
rect 153500 29900 153600 30000
rect 153500 30000 153600 30100
rect 153500 30100 153600 30200
rect 153500 30200 153600 30300
rect 153500 30300 153600 30400
rect 153500 30400 153600 30500
rect 153500 30500 153600 30600
rect 153500 30600 153600 30700
rect 153500 30700 153600 30800
rect 153500 30800 153600 30900
rect 153500 30900 153600 31000
rect 153500 31000 153600 31100
rect 153500 31100 153600 31200
rect 153500 31200 153600 31300
rect 153500 31300 153600 31400
rect 153500 31400 153600 31500
rect 153500 31500 153600 31600
rect 153500 31600 153600 31700
rect 153500 31700 153600 31800
rect 153500 31800 153600 31900
rect 153500 31900 153600 32000
rect 153500 32000 153600 32100
rect 153600 26500 153700 26600
rect 153600 26600 153700 26700
rect 153600 26700 153700 26800
rect 153600 26800 153700 26900
rect 153600 26900 153700 27000
rect 153600 27000 153700 27100
rect 153600 27100 153700 27200
rect 153600 27200 153700 27300
rect 153600 27300 153700 27400
rect 153600 27400 153700 27500
rect 153600 27500 153700 27600
rect 153600 27600 153700 27700
rect 153600 27700 153700 27800
rect 153600 27800 153700 27900
rect 153600 27900 153700 28000
rect 153600 28000 153700 28100
rect 153600 28100 153700 28200
rect 153600 28200 153700 28300
rect 153600 28300 153700 28400
rect 153600 28400 153700 28500
rect 153600 28500 153700 28600
rect 153600 28600 153700 28700
rect 153600 28700 153700 28800
rect 153600 28800 153700 28900
rect 153600 28900 153700 29000
rect 153600 29000 153700 29100
rect 153600 29100 153700 29200
rect 153600 29200 153700 29300
rect 153600 29300 153700 29400
rect 153600 29400 153700 29500
rect 153600 29500 153700 29600
rect 153600 29600 153700 29700
rect 153600 29700 153700 29800
rect 153600 29800 153700 29900
rect 153600 29900 153700 30000
rect 153600 30000 153700 30100
rect 153600 30100 153700 30200
rect 153600 30200 153700 30300
rect 153600 30300 153700 30400
rect 153600 30400 153700 30500
rect 153600 30500 153700 30600
rect 153600 30600 153700 30700
rect 153600 30700 153700 30800
rect 153600 30800 153700 30900
rect 153600 30900 153700 31000
rect 153600 31000 153700 31100
rect 153600 31100 153700 31200
rect 153600 31200 153700 31300
rect 153600 31300 153700 31400
rect 153600 31400 153700 31500
rect 153600 31500 153700 31600
rect 153600 31600 153700 31700
rect 153600 31700 153700 31800
rect 153600 31800 153700 31900
rect 153600 31900 153700 32000
rect 153600 32000 153700 32100
rect 153600 32100 153700 32200
rect 153700 26400 153800 26500
rect 153700 26500 153800 26600
rect 153700 26600 153800 26700
rect 153700 26700 153800 26800
rect 153700 26800 153800 26900
rect 153700 26900 153800 27000
rect 153700 27000 153800 27100
rect 153700 27100 153800 27200
rect 153700 27200 153800 27300
rect 153700 27300 153800 27400
rect 153700 27400 153800 27500
rect 153700 27500 153800 27600
rect 153700 27600 153800 27700
rect 153700 27700 153800 27800
rect 153700 27800 153800 27900
rect 153700 27900 153800 28000
rect 153700 28000 153800 28100
rect 153700 28100 153800 28200
rect 153700 28200 153800 28300
rect 153700 28300 153800 28400
rect 153700 28400 153800 28500
rect 153700 28500 153800 28600
rect 153700 28600 153800 28700
rect 153700 28700 153800 28800
rect 153700 28800 153800 28900
rect 153700 28900 153800 29000
rect 153700 29000 153800 29100
rect 153700 29100 153800 29200
rect 153700 29200 153800 29300
rect 153700 29300 153800 29400
rect 153700 29400 153800 29500
rect 153700 29500 153800 29600
rect 153700 29600 153800 29700
rect 153700 29700 153800 29800
rect 153700 29800 153800 29900
rect 153700 29900 153800 30000
rect 153700 30000 153800 30100
rect 153700 30100 153800 30200
rect 153700 30200 153800 30300
rect 153700 30300 153800 30400
rect 153700 30400 153800 30500
rect 153700 30500 153800 30600
rect 153700 30600 153800 30700
rect 153700 30700 153800 30800
rect 153700 30800 153800 30900
rect 153700 30900 153800 31000
rect 153700 31000 153800 31100
rect 153700 31100 153800 31200
rect 153700 31200 153800 31300
rect 153700 31300 153800 31400
rect 153700 31400 153800 31500
rect 153700 31500 153800 31600
rect 153700 31600 153800 31700
rect 153700 31700 153800 31800
rect 153700 31800 153800 31900
rect 153700 31900 153800 32000
rect 153700 32000 153800 32100
rect 153700 32100 153800 32200
rect 153700 32200 153800 32300
rect 153700 32300 153800 32400
rect 153800 26300 153900 26400
rect 153800 26400 153900 26500
rect 153800 26500 153900 26600
rect 153800 26600 153900 26700
rect 153800 26700 153900 26800
rect 153800 26800 153900 26900
rect 153800 26900 153900 27000
rect 153800 27000 153900 27100
rect 153800 27100 153900 27200
rect 153800 27200 153900 27300
rect 153800 27300 153900 27400
rect 153800 27400 153900 27500
rect 153800 27500 153900 27600
rect 153800 27600 153900 27700
rect 153800 27700 153900 27800
rect 153800 27800 153900 27900
rect 153800 27900 153900 28000
rect 153800 28000 153900 28100
rect 153800 28100 153900 28200
rect 153800 28200 153900 28300
rect 153800 28300 153900 28400
rect 153800 28400 153900 28500
rect 153800 28500 153900 28600
rect 153800 28600 153900 28700
rect 153800 28700 153900 28800
rect 153800 28800 153900 28900
rect 153800 28900 153900 29000
rect 153800 29000 153900 29100
rect 153800 29100 153900 29200
rect 153800 29200 153900 29300
rect 153800 29300 153900 29400
rect 153800 29400 153900 29500
rect 153800 29500 153900 29600
rect 153800 29600 153900 29700
rect 153800 29700 153900 29800
rect 153800 29800 153900 29900
rect 153800 29900 153900 30000
rect 153800 30000 153900 30100
rect 153800 30100 153900 30200
rect 153800 30200 153900 30300
rect 153800 30300 153900 30400
rect 153800 30400 153900 30500
rect 153800 30500 153900 30600
rect 153800 30600 153900 30700
rect 153800 30700 153900 30800
rect 153800 30800 153900 30900
rect 153800 30900 153900 31000
rect 153800 31000 153900 31100
rect 153800 31100 153900 31200
rect 153800 31200 153900 31300
rect 153800 31300 153900 31400
rect 153800 31400 153900 31500
rect 153800 31500 153900 31600
rect 153800 31600 153900 31700
rect 153800 31700 153900 31800
rect 153800 31800 153900 31900
rect 153800 31900 153900 32000
rect 153800 32000 153900 32100
rect 153800 32100 153900 32200
rect 153800 32200 153900 32300
rect 153800 32300 153900 32400
rect 153900 26200 154000 26300
rect 153900 26300 154000 26400
rect 153900 26400 154000 26500
rect 153900 26500 154000 26600
rect 153900 26600 154000 26700
rect 153900 26700 154000 26800
rect 153900 26800 154000 26900
rect 153900 26900 154000 27000
rect 153900 27000 154000 27100
rect 153900 27100 154000 27200
rect 153900 27200 154000 27300
rect 153900 27300 154000 27400
rect 153900 27400 154000 27500
rect 153900 27500 154000 27600
rect 153900 27600 154000 27700
rect 153900 27700 154000 27800
rect 153900 27800 154000 27900
rect 153900 27900 154000 28000
rect 153900 28000 154000 28100
rect 153900 28100 154000 28200
rect 153900 28200 154000 28300
rect 153900 28300 154000 28400
rect 153900 28400 154000 28500
rect 153900 28500 154000 28600
rect 153900 28600 154000 28700
rect 153900 28700 154000 28800
rect 153900 28800 154000 28900
rect 153900 28900 154000 29000
rect 153900 29000 154000 29100
rect 153900 29100 154000 29200
rect 153900 29200 154000 29300
rect 153900 29300 154000 29400
rect 153900 29400 154000 29500
rect 153900 29500 154000 29600
rect 153900 29600 154000 29700
rect 153900 29700 154000 29800
rect 153900 29800 154000 29900
rect 153900 29900 154000 30000
rect 153900 30000 154000 30100
rect 153900 30100 154000 30200
rect 153900 30200 154000 30300
rect 153900 30300 154000 30400
rect 153900 30400 154000 30500
rect 153900 30500 154000 30600
rect 153900 30600 154000 30700
rect 153900 30700 154000 30800
rect 153900 30800 154000 30900
rect 153900 30900 154000 31000
rect 153900 31000 154000 31100
rect 153900 31100 154000 31200
rect 153900 31200 154000 31300
rect 153900 31300 154000 31400
rect 153900 31400 154000 31500
rect 153900 31500 154000 31600
rect 153900 31600 154000 31700
rect 153900 31700 154000 31800
rect 153900 31800 154000 31900
rect 153900 31900 154000 32000
rect 153900 32000 154000 32100
rect 153900 32100 154000 32200
rect 153900 32200 154000 32300
rect 153900 32300 154000 32400
rect 153900 32400 154000 32500
rect 153900 32500 154000 32600
rect 154000 26100 154100 26200
rect 154000 26200 154100 26300
rect 154000 26300 154100 26400
rect 154000 26400 154100 26500
rect 154000 26500 154100 26600
rect 154000 26600 154100 26700
rect 154000 26700 154100 26800
rect 154000 26800 154100 26900
rect 154000 26900 154100 27000
rect 154000 27000 154100 27100
rect 154000 27100 154100 27200
rect 154000 27200 154100 27300
rect 154000 27300 154100 27400
rect 154000 27400 154100 27500
rect 154000 27500 154100 27600
rect 154000 27600 154100 27700
rect 154000 27700 154100 27800
rect 154000 27800 154100 27900
rect 154000 27900 154100 28000
rect 154000 28000 154100 28100
rect 154000 28100 154100 28200
rect 154000 28200 154100 28300
rect 154000 28300 154100 28400
rect 154000 28400 154100 28500
rect 154000 28500 154100 28600
rect 154000 28600 154100 28700
rect 154000 28700 154100 28800
rect 154000 28800 154100 28900
rect 154000 28900 154100 29000
rect 154000 29000 154100 29100
rect 154000 29100 154100 29200
rect 154000 29200 154100 29300
rect 154000 29300 154100 29400
rect 154000 29400 154100 29500
rect 154000 29500 154100 29600
rect 154000 29600 154100 29700
rect 154000 29700 154100 29800
rect 154000 29800 154100 29900
rect 154000 29900 154100 30000
rect 154000 30000 154100 30100
rect 154000 30100 154100 30200
rect 154000 30200 154100 30300
rect 154000 30300 154100 30400
rect 154000 30400 154100 30500
rect 154000 30500 154100 30600
rect 154000 30600 154100 30700
rect 154000 30700 154100 30800
rect 154000 30800 154100 30900
rect 154000 30900 154100 31000
rect 154000 31000 154100 31100
rect 154000 31100 154100 31200
rect 154000 31200 154100 31300
rect 154000 31300 154100 31400
rect 154000 31400 154100 31500
rect 154000 31500 154100 31600
rect 154000 31600 154100 31700
rect 154000 31700 154100 31800
rect 154000 31800 154100 31900
rect 154000 31900 154100 32000
rect 154000 32000 154100 32100
rect 154000 32100 154100 32200
rect 154000 32200 154100 32300
rect 154000 32300 154100 32400
rect 154000 32400 154100 32500
rect 154000 32500 154100 32600
rect 154000 32600 154100 32700
rect 154100 26000 154200 26100
rect 154100 26100 154200 26200
rect 154100 26200 154200 26300
rect 154100 26300 154200 26400
rect 154100 26400 154200 26500
rect 154100 26500 154200 26600
rect 154100 26600 154200 26700
rect 154100 26700 154200 26800
rect 154100 26800 154200 26900
rect 154100 26900 154200 27000
rect 154100 27000 154200 27100
rect 154100 27100 154200 27200
rect 154100 27200 154200 27300
rect 154100 27300 154200 27400
rect 154100 27400 154200 27500
rect 154100 27500 154200 27600
rect 154100 27600 154200 27700
rect 154100 27700 154200 27800
rect 154100 27800 154200 27900
rect 154100 27900 154200 28000
rect 154100 28000 154200 28100
rect 154100 28100 154200 28200
rect 154100 28200 154200 28300
rect 154100 28300 154200 28400
rect 154100 28400 154200 28500
rect 154100 28500 154200 28600
rect 154100 28600 154200 28700
rect 154100 28700 154200 28800
rect 154100 28800 154200 28900
rect 154100 28900 154200 29000
rect 154100 29000 154200 29100
rect 154100 29100 154200 29200
rect 154100 29200 154200 29300
rect 154100 29300 154200 29400
rect 154100 29400 154200 29500
rect 154100 29500 154200 29600
rect 154100 29600 154200 29700
rect 154100 29700 154200 29800
rect 154100 29800 154200 29900
rect 154100 29900 154200 30000
rect 154100 30000 154200 30100
rect 154100 30100 154200 30200
rect 154100 30200 154200 30300
rect 154100 30300 154200 30400
rect 154100 30400 154200 30500
rect 154100 30500 154200 30600
rect 154100 30600 154200 30700
rect 154100 30700 154200 30800
rect 154100 30800 154200 30900
rect 154100 30900 154200 31000
rect 154100 31000 154200 31100
rect 154100 31100 154200 31200
rect 154100 31200 154200 31300
rect 154100 31300 154200 31400
rect 154100 31400 154200 31500
rect 154100 31500 154200 31600
rect 154100 31600 154200 31700
rect 154100 31700 154200 31800
rect 154100 31800 154200 31900
rect 154100 31900 154200 32000
rect 154100 32000 154200 32100
rect 154100 32100 154200 32200
rect 154100 32200 154200 32300
rect 154100 32300 154200 32400
rect 154100 32400 154200 32500
rect 154100 32500 154200 32600
rect 154100 32600 154200 32700
rect 154100 32700 154200 32800
rect 154200 25900 154300 26000
rect 154200 26000 154300 26100
rect 154200 26100 154300 26200
rect 154200 26200 154300 26300
rect 154200 26300 154300 26400
rect 154200 26400 154300 26500
rect 154200 26500 154300 26600
rect 154200 26600 154300 26700
rect 154200 26700 154300 26800
rect 154200 26800 154300 26900
rect 154200 26900 154300 27000
rect 154200 27000 154300 27100
rect 154200 27100 154300 27200
rect 154200 27200 154300 27300
rect 154200 27300 154300 27400
rect 154200 27400 154300 27500
rect 154200 27500 154300 27600
rect 154200 27600 154300 27700
rect 154200 27700 154300 27800
rect 154200 27800 154300 27900
rect 154200 27900 154300 28000
rect 154200 28000 154300 28100
rect 154200 28100 154300 28200
rect 154200 28200 154300 28300
rect 154200 28300 154300 28400
rect 154200 28400 154300 28500
rect 154200 28500 154300 28600
rect 154200 28600 154300 28700
rect 154200 28700 154300 28800
rect 154200 28800 154300 28900
rect 154200 28900 154300 29000
rect 154200 29000 154300 29100
rect 154200 29100 154300 29200
rect 154200 29200 154300 29300
rect 154200 29300 154300 29400
rect 154200 29400 154300 29500
rect 154200 29500 154300 29600
rect 154200 29600 154300 29700
rect 154200 29700 154300 29800
rect 154200 29800 154300 29900
rect 154200 29900 154300 30000
rect 154200 30000 154300 30100
rect 154200 30100 154300 30200
rect 154200 30200 154300 30300
rect 154200 30300 154300 30400
rect 154200 30400 154300 30500
rect 154200 30500 154300 30600
rect 154200 30600 154300 30700
rect 154200 30700 154300 30800
rect 154200 30800 154300 30900
rect 154200 30900 154300 31000
rect 154200 31000 154300 31100
rect 154200 31100 154300 31200
rect 154200 31200 154300 31300
rect 154200 31300 154300 31400
rect 154200 31400 154300 31500
rect 154200 31500 154300 31600
rect 154200 31600 154300 31700
rect 154200 31700 154300 31800
rect 154200 31800 154300 31900
rect 154200 31900 154300 32000
rect 154200 32000 154300 32100
rect 154200 32100 154300 32200
rect 154200 32200 154300 32300
rect 154200 32300 154300 32400
rect 154200 32400 154300 32500
rect 154200 32500 154300 32600
rect 154200 32600 154300 32700
rect 154200 32700 154300 32800
rect 154200 32800 154300 32900
rect 154300 25800 154400 25900
rect 154300 25900 154400 26000
rect 154300 26000 154400 26100
rect 154300 26100 154400 26200
rect 154300 26200 154400 26300
rect 154300 26300 154400 26400
rect 154300 26400 154400 26500
rect 154300 26500 154400 26600
rect 154300 26600 154400 26700
rect 154300 26700 154400 26800
rect 154300 26800 154400 26900
rect 154300 26900 154400 27000
rect 154300 27000 154400 27100
rect 154300 27100 154400 27200
rect 154300 27200 154400 27300
rect 154300 27300 154400 27400
rect 154300 27400 154400 27500
rect 154300 27500 154400 27600
rect 154300 27600 154400 27700
rect 154300 27700 154400 27800
rect 154300 27800 154400 27900
rect 154300 27900 154400 28000
rect 154300 28000 154400 28100
rect 154300 28100 154400 28200
rect 154300 28200 154400 28300
rect 154300 28300 154400 28400
rect 154300 28400 154400 28500
rect 154300 28500 154400 28600
rect 154300 28600 154400 28700
rect 154300 28700 154400 28800
rect 154300 28800 154400 28900
rect 154300 28900 154400 29000
rect 154300 29000 154400 29100
rect 154300 29100 154400 29200
rect 154300 29200 154400 29300
rect 154300 29300 154400 29400
rect 154300 29400 154400 29500
rect 154300 29500 154400 29600
rect 154300 29600 154400 29700
rect 154300 29700 154400 29800
rect 154300 29800 154400 29900
rect 154300 29900 154400 30000
rect 154300 30000 154400 30100
rect 154300 30100 154400 30200
rect 154300 30200 154400 30300
rect 154300 30300 154400 30400
rect 154300 30400 154400 30500
rect 154300 30500 154400 30600
rect 154300 30600 154400 30700
rect 154300 30700 154400 30800
rect 154300 30800 154400 30900
rect 154300 30900 154400 31000
rect 154300 31000 154400 31100
rect 154300 31100 154400 31200
rect 154300 31200 154400 31300
rect 154300 31300 154400 31400
rect 154300 31400 154400 31500
rect 154300 31500 154400 31600
rect 154300 31600 154400 31700
rect 154300 31700 154400 31800
rect 154300 31800 154400 31900
rect 154300 31900 154400 32000
rect 154300 32000 154400 32100
rect 154300 32100 154400 32200
rect 154300 32200 154400 32300
rect 154300 32300 154400 32400
rect 154300 32400 154400 32500
rect 154300 32500 154400 32600
rect 154300 32600 154400 32700
rect 154300 32700 154400 32800
rect 154300 32800 154400 32900
rect 154300 32900 154400 33000
rect 154400 25700 154500 25800
rect 154400 25800 154500 25900
rect 154400 25900 154500 26000
rect 154400 26000 154500 26100
rect 154400 26100 154500 26200
rect 154400 26200 154500 26300
rect 154400 26300 154500 26400
rect 154400 26400 154500 26500
rect 154400 26500 154500 26600
rect 154400 26600 154500 26700
rect 154400 26700 154500 26800
rect 154400 26800 154500 26900
rect 154400 26900 154500 27000
rect 154400 27000 154500 27100
rect 154400 27100 154500 27200
rect 154400 27200 154500 27300
rect 154400 27300 154500 27400
rect 154400 27400 154500 27500
rect 154400 27500 154500 27600
rect 154400 27600 154500 27700
rect 154400 27700 154500 27800
rect 154400 27800 154500 27900
rect 154400 27900 154500 28000
rect 154400 28000 154500 28100
rect 154400 28100 154500 28200
rect 154400 28200 154500 28300
rect 154400 28300 154500 28400
rect 154400 28400 154500 28500
rect 154400 28500 154500 28600
rect 154400 28600 154500 28700
rect 154400 28700 154500 28800
rect 154400 28800 154500 28900
rect 154400 28900 154500 29000
rect 154400 29000 154500 29100
rect 154400 29100 154500 29200
rect 154400 29200 154500 29300
rect 154400 29300 154500 29400
rect 154400 29400 154500 29500
rect 154400 29500 154500 29600
rect 154400 29600 154500 29700
rect 154400 29700 154500 29800
rect 154400 29800 154500 29900
rect 154400 29900 154500 30000
rect 154400 30000 154500 30100
rect 154400 30100 154500 30200
rect 154400 30200 154500 30300
rect 154400 30300 154500 30400
rect 154400 30400 154500 30500
rect 154400 30500 154500 30600
rect 154400 30600 154500 30700
rect 154400 30700 154500 30800
rect 154400 30800 154500 30900
rect 154400 30900 154500 31000
rect 154400 31000 154500 31100
rect 154400 31100 154500 31200
rect 154400 31200 154500 31300
rect 154400 31300 154500 31400
rect 154400 31400 154500 31500
rect 154400 31500 154500 31600
rect 154400 31600 154500 31700
rect 154400 31700 154500 31800
rect 154400 31800 154500 31900
rect 154400 31900 154500 32000
rect 154400 32000 154500 32100
rect 154400 32100 154500 32200
rect 154400 32200 154500 32300
rect 154400 32300 154500 32400
rect 154400 32400 154500 32500
rect 154400 32500 154500 32600
rect 154400 32600 154500 32700
rect 154400 32700 154500 32800
rect 154400 32800 154500 32900
rect 154400 32900 154500 33000
rect 154400 33000 154500 33100
rect 154500 25600 154600 25700
rect 154500 25700 154600 25800
rect 154500 25800 154600 25900
rect 154500 25900 154600 26000
rect 154500 26000 154600 26100
rect 154500 26100 154600 26200
rect 154500 26200 154600 26300
rect 154500 26300 154600 26400
rect 154500 26400 154600 26500
rect 154500 26500 154600 26600
rect 154500 26600 154600 26700
rect 154500 26700 154600 26800
rect 154500 26800 154600 26900
rect 154500 26900 154600 27000
rect 154500 27000 154600 27100
rect 154500 27100 154600 27200
rect 154500 27200 154600 27300
rect 154500 27300 154600 27400
rect 154500 27400 154600 27500
rect 154500 27500 154600 27600
rect 154500 27600 154600 27700
rect 154500 27700 154600 27800
rect 154500 27800 154600 27900
rect 154500 27900 154600 28000
rect 154500 28000 154600 28100
rect 154500 28100 154600 28200
rect 154500 28200 154600 28300
rect 154500 28300 154600 28400
rect 154500 28400 154600 28500
rect 154500 28500 154600 28600
rect 154500 28600 154600 28700
rect 154500 28800 154600 28900
rect 154500 28900 154600 29000
rect 154500 29000 154600 29100
rect 154500 29100 154600 29200
rect 154500 29200 154600 29300
rect 154500 29300 154600 29400
rect 154500 29400 154600 29500
rect 154500 29500 154600 29600
rect 154500 29600 154600 29700
rect 154500 29700 154600 29800
rect 154500 29800 154600 29900
rect 154500 29900 154600 30000
rect 154500 30000 154600 30100
rect 154500 30200 154600 30300
rect 154500 30300 154600 30400
rect 154500 30400 154600 30500
rect 154500 30500 154600 30600
rect 154500 30600 154600 30700
rect 154500 30700 154600 30800
rect 154500 30800 154600 30900
rect 154500 30900 154600 31000
rect 154500 31000 154600 31100
rect 154500 31100 154600 31200
rect 154500 31200 154600 31300
rect 154500 31300 154600 31400
rect 154500 31400 154600 31500
rect 154500 31500 154600 31600
rect 154500 31600 154600 31700
rect 154500 31700 154600 31800
rect 154500 31800 154600 31900
rect 154500 31900 154600 32000
rect 154500 32000 154600 32100
rect 154500 32100 154600 32200
rect 154500 32200 154600 32300
rect 154500 32300 154600 32400
rect 154500 32400 154600 32500
rect 154500 32500 154600 32600
rect 154500 32600 154600 32700
rect 154500 32700 154600 32800
rect 154500 32800 154600 32900
rect 154500 32900 154600 33000
rect 154500 33000 154600 33100
rect 154500 33100 154600 33200
rect 154600 25500 154700 25600
rect 154600 25600 154700 25700
rect 154600 25700 154700 25800
rect 154600 25800 154700 25900
rect 154600 25900 154700 26000
rect 154600 26000 154700 26100
rect 154600 26100 154700 26200
rect 154600 26200 154700 26300
rect 154600 26300 154700 26400
rect 154600 26400 154700 26500
rect 154600 26500 154700 26600
rect 154600 26600 154700 26700
rect 154600 26700 154700 26800
rect 154600 26800 154700 26900
rect 154600 26900 154700 27000
rect 154600 27000 154700 27100
rect 154600 27100 154700 27200
rect 154600 27200 154700 27300
rect 154600 27300 154700 27400
rect 154600 27400 154700 27500
rect 154600 27500 154700 27600
rect 154600 27600 154700 27700
rect 154600 27700 154700 27800
rect 154600 27800 154700 27900
rect 154600 27900 154700 28000
rect 154600 28000 154700 28100
rect 154600 28100 154700 28200
rect 154600 28200 154700 28300
rect 154600 28300 154700 28400
rect 154600 28400 154700 28500
rect 154600 28500 154700 28600
rect 154600 30300 154700 30400
rect 154600 30400 154700 30500
rect 154600 30500 154700 30600
rect 154600 30600 154700 30700
rect 154600 30700 154700 30800
rect 154600 30800 154700 30900
rect 154600 30900 154700 31000
rect 154600 31000 154700 31100
rect 154600 31100 154700 31200
rect 154600 31200 154700 31300
rect 154600 31300 154700 31400
rect 154600 31400 154700 31500
rect 154600 31500 154700 31600
rect 154600 31600 154700 31700
rect 154600 31700 154700 31800
rect 154600 31800 154700 31900
rect 154600 31900 154700 32000
rect 154600 32000 154700 32100
rect 154600 32100 154700 32200
rect 154600 32200 154700 32300
rect 154600 32300 154700 32400
rect 154600 32400 154700 32500
rect 154600 32500 154700 32600
rect 154600 32600 154700 32700
rect 154600 32700 154700 32800
rect 154600 32800 154700 32900
rect 154600 32900 154700 33000
rect 154600 33000 154700 33100
rect 154600 33100 154700 33200
rect 154600 33200 154700 33300
rect 154700 25400 154800 25500
rect 154700 25500 154800 25600
rect 154700 25600 154800 25700
rect 154700 25700 154800 25800
rect 154700 25800 154800 25900
rect 154700 25900 154800 26000
rect 154700 26000 154800 26100
rect 154700 26100 154800 26200
rect 154700 26200 154800 26300
rect 154700 26300 154800 26400
rect 154700 26400 154800 26500
rect 154700 26500 154800 26600
rect 154700 26600 154800 26700
rect 154700 26700 154800 26800
rect 154700 26800 154800 26900
rect 154700 26900 154800 27000
rect 154700 27000 154800 27100
rect 154700 27100 154800 27200
rect 154700 27200 154800 27300
rect 154700 27300 154800 27400
rect 154700 27400 154800 27500
rect 154700 27500 154800 27600
rect 154700 27600 154800 27700
rect 154700 27700 154800 27800
rect 154700 27800 154800 27900
rect 154700 27900 154800 28000
rect 154700 28000 154800 28100
rect 154700 28100 154800 28200
rect 154700 28200 154800 28300
rect 154700 28300 154800 28400
rect 154700 28400 154800 28500
rect 154700 30400 154800 30500
rect 154700 30500 154800 30600
rect 154700 30600 154800 30700
rect 154700 30700 154800 30800
rect 154700 30800 154800 30900
rect 154700 30900 154800 31000
rect 154700 31000 154800 31100
rect 154700 31100 154800 31200
rect 154700 31200 154800 31300
rect 154700 31300 154800 31400
rect 154700 31400 154800 31500
rect 154700 31500 154800 31600
rect 154700 31600 154800 31700
rect 154700 31700 154800 31800
rect 154700 31800 154800 31900
rect 154700 31900 154800 32000
rect 154700 32000 154800 32100
rect 154700 32100 154800 32200
rect 154700 32200 154800 32300
rect 154700 32300 154800 32400
rect 154700 32400 154800 32500
rect 154700 32500 154800 32600
rect 154700 32600 154800 32700
rect 154700 32700 154800 32800
rect 154700 32800 154800 32900
rect 154700 32900 154800 33000
rect 154700 33000 154800 33100
rect 154700 33100 154800 33200
rect 154700 33200 154800 33300
rect 154700 33300 154800 33400
rect 154800 25300 154900 25400
rect 154800 25400 154900 25500
rect 154800 25500 154900 25600
rect 154800 25600 154900 25700
rect 154800 25700 154900 25800
rect 154800 25800 154900 25900
rect 154800 25900 154900 26000
rect 154800 26000 154900 26100
rect 154800 26100 154900 26200
rect 154800 26200 154900 26300
rect 154800 26300 154900 26400
rect 154800 26400 154900 26500
rect 154800 26500 154900 26600
rect 154800 26600 154900 26700
rect 154800 26700 154900 26800
rect 154800 26800 154900 26900
rect 154800 26900 154900 27000
rect 154800 27000 154900 27100
rect 154800 27100 154900 27200
rect 154800 27200 154900 27300
rect 154800 27300 154900 27400
rect 154800 27400 154900 27500
rect 154800 27500 154900 27600
rect 154800 27600 154900 27700
rect 154800 27700 154900 27800
rect 154800 27800 154900 27900
rect 154800 27900 154900 28000
rect 154800 28000 154900 28100
rect 154800 28100 154900 28200
rect 154800 28200 154900 28300
rect 154800 28300 154900 28400
rect 154800 30500 154900 30600
rect 154800 30600 154900 30700
rect 154800 30700 154900 30800
rect 154800 30800 154900 30900
rect 154800 30900 154900 31000
rect 154800 31000 154900 31100
rect 154800 31100 154900 31200
rect 154800 31200 154900 31300
rect 154800 31300 154900 31400
rect 154800 31400 154900 31500
rect 154800 31500 154900 31600
rect 154800 31600 154900 31700
rect 154800 31700 154900 31800
rect 154800 31800 154900 31900
rect 154800 31900 154900 32000
rect 154800 32000 154900 32100
rect 154800 32100 154900 32200
rect 154800 32200 154900 32300
rect 154800 32300 154900 32400
rect 154800 32400 154900 32500
rect 154800 32500 154900 32600
rect 154800 32600 154900 32700
rect 154800 32700 154900 32800
rect 154800 32800 154900 32900
rect 154800 32900 154900 33000
rect 154800 33000 154900 33100
rect 154800 33100 154900 33200
rect 154800 33200 154900 33300
rect 154800 33300 154900 33400
rect 154800 33400 154900 33500
rect 154900 25200 155000 25300
rect 154900 25300 155000 25400
rect 154900 25400 155000 25500
rect 154900 25500 155000 25600
rect 154900 25600 155000 25700
rect 154900 25700 155000 25800
rect 154900 25800 155000 25900
rect 154900 25900 155000 26000
rect 154900 26000 155000 26100
rect 154900 26100 155000 26200
rect 154900 26200 155000 26300
rect 154900 26300 155000 26400
rect 154900 26400 155000 26500
rect 154900 26500 155000 26600
rect 154900 26600 155000 26700
rect 154900 26700 155000 26800
rect 154900 26800 155000 26900
rect 154900 26900 155000 27000
rect 154900 27000 155000 27100
rect 154900 27100 155000 27200
rect 154900 27200 155000 27300
rect 154900 27300 155000 27400
rect 154900 27400 155000 27500
rect 154900 27500 155000 27600
rect 154900 27600 155000 27700
rect 154900 27700 155000 27800
rect 154900 27800 155000 27900
rect 154900 27900 155000 28000
rect 154900 28000 155000 28100
rect 154900 28100 155000 28200
rect 154900 28200 155000 28300
rect 154900 30600 155000 30700
rect 154900 30700 155000 30800
rect 154900 30800 155000 30900
rect 154900 30900 155000 31000
rect 154900 31000 155000 31100
rect 154900 31100 155000 31200
rect 154900 31200 155000 31300
rect 154900 31300 155000 31400
rect 154900 31400 155000 31500
rect 154900 31500 155000 31600
rect 154900 31600 155000 31700
rect 154900 31700 155000 31800
rect 154900 31800 155000 31900
rect 154900 31900 155000 32000
rect 154900 32000 155000 32100
rect 154900 32100 155000 32200
rect 154900 32200 155000 32300
rect 154900 32300 155000 32400
rect 154900 32400 155000 32500
rect 154900 32500 155000 32600
rect 154900 32600 155000 32700
rect 154900 32700 155000 32800
rect 154900 32800 155000 32900
rect 154900 32900 155000 33000
rect 154900 33000 155000 33100
rect 154900 33100 155000 33200
rect 154900 33200 155000 33300
rect 154900 33300 155000 33400
rect 154900 33400 155000 33500
rect 154900 33500 155000 33600
rect 155000 25100 155100 25200
rect 155000 25200 155100 25300
rect 155000 25300 155100 25400
rect 155000 25400 155100 25500
rect 155000 25500 155100 25600
rect 155000 25600 155100 25700
rect 155000 25700 155100 25800
rect 155000 25800 155100 25900
rect 155000 25900 155100 26000
rect 155000 26000 155100 26100
rect 155000 26100 155100 26200
rect 155000 26200 155100 26300
rect 155000 26300 155100 26400
rect 155000 26400 155100 26500
rect 155000 26500 155100 26600
rect 155000 26600 155100 26700
rect 155000 26700 155100 26800
rect 155000 26800 155100 26900
rect 155000 26900 155100 27000
rect 155000 27000 155100 27100
rect 155000 27100 155100 27200
rect 155000 27200 155100 27300
rect 155000 27300 155100 27400
rect 155000 27400 155100 27500
rect 155000 27500 155100 27600
rect 155000 27600 155100 27700
rect 155000 27700 155100 27800
rect 155000 27800 155100 27900
rect 155000 27900 155100 28000
rect 155000 28000 155100 28100
rect 155000 28100 155100 28200
rect 155000 30700 155100 30800
rect 155000 30800 155100 30900
rect 155000 30900 155100 31000
rect 155000 31000 155100 31100
rect 155000 31100 155100 31200
rect 155000 31200 155100 31300
rect 155000 31300 155100 31400
rect 155000 31400 155100 31500
rect 155000 31500 155100 31600
rect 155000 31600 155100 31700
rect 155000 31700 155100 31800
rect 155000 31800 155100 31900
rect 155000 31900 155100 32000
rect 155000 32000 155100 32100
rect 155000 32100 155100 32200
rect 155000 32200 155100 32300
rect 155000 32300 155100 32400
rect 155000 32400 155100 32500
rect 155000 32500 155100 32600
rect 155000 32600 155100 32700
rect 155000 32700 155100 32800
rect 155000 32800 155100 32900
rect 155000 32900 155100 33000
rect 155000 33000 155100 33100
rect 155000 33100 155100 33200
rect 155000 33200 155100 33300
rect 155000 33300 155100 33400
rect 155000 33400 155100 33500
rect 155000 33500 155100 33600
rect 155000 33600 155100 33700
rect 155000 33700 155100 33800
rect 155100 25000 155200 25100
rect 155100 25100 155200 25200
rect 155100 25200 155200 25300
rect 155100 25300 155200 25400
rect 155100 25400 155200 25500
rect 155100 25500 155200 25600
rect 155100 25600 155200 25700
rect 155100 25700 155200 25800
rect 155100 25800 155200 25900
rect 155100 25900 155200 26000
rect 155100 26000 155200 26100
rect 155100 26100 155200 26200
rect 155100 26200 155200 26300
rect 155100 26300 155200 26400
rect 155100 26400 155200 26500
rect 155100 26500 155200 26600
rect 155100 26600 155200 26700
rect 155100 26700 155200 26800
rect 155100 26800 155200 26900
rect 155100 26900 155200 27000
rect 155100 27000 155200 27100
rect 155100 27100 155200 27200
rect 155100 27200 155200 27300
rect 155100 27300 155200 27400
rect 155100 27400 155200 27500
rect 155100 27500 155200 27600
rect 155100 27600 155200 27700
rect 155100 27700 155200 27800
rect 155100 27800 155200 27900
rect 155100 27900 155200 28000
rect 155100 28000 155200 28100
rect 155100 30800 155200 30900
rect 155100 30900 155200 31000
rect 155100 31000 155200 31100
rect 155100 31100 155200 31200
rect 155100 31200 155200 31300
rect 155100 31300 155200 31400
rect 155100 31400 155200 31500
rect 155100 31500 155200 31600
rect 155100 31600 155200 31700
rect 155100 31700 155200 31800
rect 155100 31800 155200 31900
rect 155100 31900 155200 32000
rect 155100 32000 155200 32100
rect 155100 32100 155200 32200
rect 155100 32200 155200 32300
rect 155100 32300 155200 32400
rect 155100 32400 155200 32500
rect 155100 32500 155200 32600
rect 155100 32600 155200 32700
rect 155100 32700 155200 32800
rect 155100 32800 155200 32900
rect 155100 32900 155200 33000
rect 155100 33000 155200 33100
rect 155100 33100 155200 33200
rect 155100 33200 155200 33300
rect 155100 33300 155200 33400
rect 155100 33400 155200 33500
rect 155100 33500 155200 33600
rect 155100 33600 155200 33700
rect 155100 33700 155200 33800
rect 155100 33800 155200 33900
rect 155200 24900 155300 25000
rect 155200 25000 155300 25100
rect 155200 25100 155300 25200
rect 155200 25200 155300 25300
rect 155200 25300 155300 25400
rect 155200 25400 155300 25500
rect 155200 25500 155300 25600
rect 155200 25600 155300 25700
rect 155200 25700 155300 25800
rect 155200 25800 155300 25900
rect 155200 25900 155300 26000
rect 155200 26000 155300 26100
rect 155200 26100 155300 26200
rect 155200 26200 155300 26300
rect 155200 26300 155300 26400
rect 155200 26400 155300 26500
rect 155200 26500 155300 26600
rect 155200 26600 155300 26700
rect 155200 26700 155300 26800
rect 155200 26800 155300 26900
rect 155200 26900 155300 27000
rect 155200 27000 155300 27100
rect 155200 27100 155300 27200
rect 155200 27200 155300 27300
rect 155200 27300 155300 27400
rect 155200 27400 155300 27500
rect 155200 27500 155300 27600
rect 155200 27600 155300 27700
rect 155200 27700 155300 27800
rect 155200 27800 155300 27900
rect 155200 27900 155300 28000
rect 155200 30900 155300 31000
rect 155200 31000 155300 31100
rect 155200 31100 155300 31200
rect 155200 31200 155300 31300
rect 155200 31300 155300 31400
rect 155200 31400 155300 31500
rect 155200 31500 155300 31600
rect 155200 31600 155300 31700
rect 155200 31700 155300 31800
rect 155200 31800 155300 31900
rect 155200 31900 155300 32000
rect 155200 32000 155300 32100
rect 155200 32100 155300 32200
rect 155200 32200 155300 32300
rect 155200 32300 155300 32400
rect 155200 32400 155300 32500
rect 155200 32500 155300 32600
rect 155200 32600 155300 32700
rect 155200 32700 155300 32800
rect 155200 32800 155300 32900
rect 155200 32900 155300 33000
rect 155200 33000 155300 33100
rect 155200 33100 155300 33200
rect 155200 33200 155300 33300
rect 155200 33300 155300 33400
rect 155200 33400 155300 33500
rect 155200 33500 155300 33600
rect 155200 33600 155300 33700
rect 155200 33700 155300 33800
rect 155200 33800 155300 33900
rect 155200 33900 155300 34000
rect 155300 24800 155400 24900
rect 155300 24900 155400 25000
rect 155300 25000 155400 25100
rect 155300 25100 155400 25200
rect 155300 25200 155400 25300
rect 155300 25300 155400 25400
rect 155300 25400 155400 25500
rect 155300 25500 155400 25600
rect 155300 25600 155400 25700
rect 155300 25700 155400 25800
rect 155300 25800 155400 25900
rect 155300 25900 155400 26000
rect 155300 26000 155400 26100
rect 155300 26100 155400 26200
rect 155300 26200 155400 26300
rect 155300 26300 155400 26400
rect 155300 26400 155400 26500
rect 155300 26500 155400 26600
rect 155300 26600 155400 26700
rect 155300 26700 155400 26800
rect 155300 26800 155400 26900
rect 155300 26900 155400 27000
rect 155300 27000 155400 27100
rect 155300 27100 155400 27200
rect 155300 27200 155400 27300
rect 155300 27300 155400 27400
rect 155300 27400 155400 27500
rect 155300 27500 155400 27600
rect 155300 27600 155400 27700
rect 155300 27700 155400 27800
rect 155300 27800 155400 27900
rect 155300 31000 155400 31100
rect 155300 31100 155400 31200
rect 155300 31200 155400 31300
rect 155300 31300 155400 31400
rect 155300 31400 155400 31500
rect 155300 31500 155400 31600
rect 155300 31600 155400 31700
rect 155300 31700 155400 31800
rect 155300 31800 155400 31900
rect 155300 31900 155400 32000
rect 155300 32000 155400 32100
rect 155300 32100 155400 32200
rect 155300 32200 155400 32300
rect 155300 32300 155400 32400
rect 155300 32400 155400 32500
rect 155300 32500 155400 32600
rect 155300 32600 155400 32700
rect 155300 32700 155400 32800
rect 155300 32800 155400 32900
rect 155300 32900 155400 33000
rect 155300 33000 155400 33100
rect 155300 33100 155400 33200
rect 155300 33200 155400 33300
rect 155300 33300 155400 33400
rect 155300 33400 155400 33500
rect 155300 33500 155400 33600
rect 155300 33600 155400 33700
rect 155300 33700 155400 33800
rect 155300 33800 155400 33900
rect 155300 33900 155400 34000
rect 155300 34000 155400 34100
rect 155400 24700 155500 24800
rect 155400 24800 155500 24900
rect 155400 24900 155500 25000
rect 155400 25000 155500 25100
rect 155400 25100 155500 25200
rect 155400 25200 155500 25300
rect 155400 25300 155500 25400
rect 155400 25400 155500 25500
rect 155400 25500 155500 25600
rect 155400 25600 155500 25700
rect 155400 25700 155500 25800
rect 155400 25800 155500 25900
rect 155400 25900 155500 26000
rect 155400 26000 155500 26100
rect 155400 26100 155500 26200
rect 155400 26200 155500 26300
rect 155400 26300 155500 26400
rect 155400 26400 155500 26500
rect 155400 26500 155500 26600
rect 155400 26600 155500 26700
rect 155400 26700 155500 26800
rect 155400 26800 155500 26900
rect 155400 26900 155500 27000
rect 155400 27000 155500 27100
rect 155400 27100 155500 27200
rect 155400 27200 155500 27300
rect 155400 27300 155500 27400
rect 155400 27400 155500 27500
rect 155400 27500 155500 27600
rect 155400 27600 155500 27700
rect 155400 27700 155500 27800
rect 155400 31100 155500 31200
rect 155400 31200 155500 31300
rect 155400 31300 155500 31400
rect 155400 31400 155500 31500
rect 155400 31500 155500 31600
rect 155400 31600 155500 31700
rect 155400 31700 155500 31800
rect 155400 31800 155500 31900
rect 155400 31900 155500 32000
rect 155400 32000 155500 32100
rect 155400 32100 155500 32200
rect 155400 32200 155500 32300
rect 155400 32300 155500 32400
rect 155400 32400 155500 32500
rect 155400 32500 155500 32600
rect 155400 32600 155500 32700
rect 155400 32700 155500 32800
rect 155400 32800 155500 32900
rect 155400 32900 155500 33000
rect 155400 33000 155500 33100
rect 155400 33100 155500 33200
rect 155400 33200 155500 33300
rect 155400 33300 155500 33400
rect 155400 33400 155500 33500
rect 155400 33500 155500 33600
rect 155400 33600 155500 33700
rect 155400 33700 155500 33800
rect 155400 33800 155500 33900
rect 155400 33900 155500 34000
rect 155400 34000 155500 34100
rect 155400 34100 155500 34200
rect 155500 24600 155600 24700
rect 155500 24700 155600 24800
rect 155500 24800 155600 24900
rect 155500 24900 155600 25000
rect 155500 25000 155600 25100
rect 155500 25100 155600 25200
rect 155500 25200 155600 25300
rect 155500 25300 155600 25400
rect 155500 25400 155600 25500
rect 155500 25500 155600 25600
rect 155500 25600 155600 25700
rect 155500 25700 155600 25800
rect 155500 25800 155600 25900
rect 155500 25900 155600 26000
rect 155500 26000 155600 26100
rect 155500 26100 155600 26200
rect 155500 26200 155600 26300
rect 155500 26300 155600 26400
rect 155500 26400 155600 26500
rect 155500 26500 155600 26600
rect 155500 26600 155600 26700
rect 155500 26700 155600 26800
rect 155500 26800 155600 26900
rect 155500 26900 155600 27000
rect 155500 27000 155600 27100
rect 155500 27100 155600 27200
rect 155500 27200 155600 27300
rect 155500 27300 155600 27400
rect 155500 27400 155600 27500
rect 155500 27500 155600 27600
rect 155500 27600 155600 27700
rect 155500 31200 155600 31300
rect 155500 31300 155600 31400
rect 155500 31400 155600 31500
rect 155500 31500 155600 31600
rect 155500 31600 155600 31700
rect 155500 31700 155600 31800
rect 155500 31800 155600 31900
rect 155500 31900 155600 32000
rect 155500 32000 155600 32100
rect 155500 32100 155600 32200
rect 155500 32200 155600 32300
rect 155500 32300 155600 32400
rect 155500 32400 155600 32500
rect 155500 32500 155600 32600
rect 155500 32600 155600 32700
rect 155500 32700 155600 32800
rect 155500 32800 155600 32900
rect 155500 32900 155600 33000
rect 155500 33000 155600 33100
rect 155500 33100 155600 33200
rect 155500 33200 155600 33300
rect 155500 33300 155600 33400
rect 155500 33400 155600 33500
rect 155500 33500 155600 33600
rect 155500 33600 155600 33700
rect 155500 33700 155600 33800
rect 155500 33800 155600 33900
rect 155500 33900 155600 34000
rect 155500 34000 155600 34100
rect 155500 34100 155600 34200
rect 155500 34200 155600 34300
rect 155600 24500 155700 24600
rect 155600 24600 155700 24700
rect 155600 24700 155700 24800
rect 155600 24800 155700 24900
rect 155600 24900 155700 25000
rect 155600 25000 155700 25100
rect 155600 25100 155700 25200
rect 155600 25200 155700 25300
rect 155600 25300 155700 25400
rect 155600 25400 155700 25500
rect 155600 25500 155700 25600
rect 155600 25600 155700 25700
rect 155600 25700 155700 25800
rect 155600 25800 155700 25900
rect 155600 25900 155700 26000
rect 155600 26000 155700 26100
rect 155600 26100 155700 26200
rect 155600 26200 155700 26300
rect 155600 26300 155700 26400
rect 155600 26400 155700 26500
rect 155600 26500 155700 26600
rect 155600 26600 155700 26700
rect 155600 26700 155700 26800
rect 155600 26800 155700 26900
rect 155600 26900 155700 27000
rect 155600 27000 155700 27100
rect 155600 27100 155700 27200
rect 155600 27200 155700 27300
rect 155600 27300 155700 27400
rect 155600 27400 155700 27500
rect 155600 27500 155700 27600
rect 155600 31300 155700 31400
rect 155600 31400 155700 31500
rect 155600 31500 155700 31600
rect 155600 31600 155700 31700
rect 155600 31700 155700 31800
rect 155600 31800 155700 31900
rect 155600 31900 155700 32000
rect 155600 32000 155700 32100
rect 155600 32100 155700 32200
rect 155600 32200 155700 32300
rect 155600 32300 155700 32400
rect 155600 32400 155700 32500
rect 155600 32500 155700 32600
rect 155600 32600 155700 32700
rect 155600 32700 155700 32800
rect 155600 32800 155700 32900
rect 155600 32900 155700 33000
rect 155600 33000 155700 33100
rect 155600 33100 155700 33200
rect 155600 33200 155700 33300
rect 155600 33300 155700 33400
rect 155600 33400 155700 33500
rect 155600 33500 155700 33600
rect 155600 33600 155700 33700
rect 155600 33700 155700 33800
rect 155600 33800 155700 33900
rect 155600 33900 155700 34000
rect 155600 34000 155700 34100
rect 155600 34100 155700 34200
rect 155600 34200 155700 34300
rect 155600 34300 155700 34400
rect 155700 24400 155800 24500
rect 155700 24500 155800 24600
rect 155700 24600 155800 24700
rect 155700 24700 155800 24800
rect 155700 24800 155800 24900
rect 155700 24900 155800 25000
rect 155700 25000 155800 25100
rect 155700 25100 155800 25200
rect 155700 25200 155800 25300
rect 155700 25300 155800 25400
rect 155700 25400 155800 25500
rect 155700 25500 155800 25600
rect 155700 25600 155800 25700
rect 155700 25700 155800 25800
rect 155700 25800 155800 25900
rect 155700 25900 155800 26000
rect 155700 26000 155800 26100
rect 155700 26100 155800 26200
rect 155700 26200 155800 26300
rect 155700 26300 155800 26400
rect 155700 26400 155800 26500
rect 155700 26500 155800 26600
rect 155700 26600 155800 26700
rect 155700 26700 155800 26800
rect 155700 26800 155800 26900
rect 155700 26900 155800 27000
rect 155700 27000 155800 27100
rect 155700 27100 155800 27200
rect 155700 27200 155800 27300
rect 155700 27300 155800 27400
rect 155700 27400 155800 27500
rect 155700 31400 155800 31500
rect 155700 31500 155800 31600
rect 155700 31600 155800 31700
rect 155700 31700 155800 31800
rect 155700 31800 155800 31900
rect 155700 31900 155800 32000
rect 155700 32000 155800 32100
rect 155700 32100 155800 32200
rect 155700 32200 155800 32300
rect 155700 32300 155800 32400
rect 155700 32400 155800 32500
rect 155700 32500 155800 32600
rect 155700 32600 155800 32700
rect 155700 32700 155800 32800
rect 155700 32800 155800 32900
rect 155700 32900 155800 33000
rect 155700 33000 155800 33100
rect 155700 33100 155800 33200
rect 155700 33200 155800 33300
rect 155700 33300 155800 33400
rect 155700 33400 155800 33500
rect 155700 33500 155800 33600
rect 155700 33600 155800 33700
rect 155700 33700 155800 33800
rect 155700 33800 155800 33900
rect 155700 33900 155800 34000
rect 155700 34000 155800 34100
rect 155700 34100 155800 34200
rect 155700 34200 155800 34300
rect 155700 34300 155800 34400
rect 155700 34400 155800 34500
rect 155800 24300 155900 24400
rect 155800 24400 155900 24500
rect 155800 24500 155900 24600
rect 155800 24600 155900 24700
rect 155800 24700 155900 24800
rect 155800 24800 155900 24900
rect 155800 24900 155900 25000
rect 155800 25000 155900 25100
rect 155800 25100 155900 25200
rect 155800 25200 155900 25300
rect 155800 25300 155900 25400
rect 155800 25400 155900 25500
rect 155800 25500 155900 25600
rect 155800 25600 155900 25700
rect 155800 25700 155900 25800
rect 155800 25800 155900 25900
rect 155800 25900 155900 26000
rect 155800 26000 155900 26100
rect 155800 26100 155900 26200
rect 155800 26200 155900 26300
rect 155800 26300 155900 26400
rect 155800 26400 155900 26500
rect 155800 26500 155900 26600
rect 155800 26600 155900 26700
rect 155800 26700 155900 26800
rect 155800 26800 155900 26900
rect 155800 26900 155900 27000
rect 155800 27000 155900 27100
rect 155800 27100 155900 27200
rect 155800 27200 155900 27300
rect 155800 27300 155900 27400
rect 155800 31500 155900 31600
rect 155800 31600 155900 31700
rect 155800 31700 155900 31800
rect 155800 31800 155900 31900
rect 155800 31900 155900 32000
rect 155800 32000 155900 32100
rect 155800 32100 155900 32200
rect 155800 32200 155900 32300
rect 155800 32300 155900 32400
rect 155800 32400 155900 32500
rect 155800 32500 155900 32600
rect 155800 32600 155900 32700
rect 155800 32700 155900 32800
rect 155800 32800 155900 32900
rect 155800 32900 155900 33000
rect 155800 33000 155900 33100
rect 155800 33100 155900 33200
rect 155800 33200 155900 33300
rect 155800 33300 155900 33400
rect 155800 33400 155900 33500
rect 155800 33500 155900 33600
rect 155800 33600 155900 33700
rect 155800 33700 155900 33800
rect 155800 33800 155900 33900
rect 155800 33900 155900 34000
rect 155800 34000 155900 34100
rect 155800 34100 155900 34200
rect 155800 34200 155900 34300
rect 155800 34300 155900 34400
rect 155800 34400 155900 34500
rect 155800 34500 155900 34600
rect 155800 34600 155900 34700
rect 155900 24300 156000 24400
rect 155900 24400 156000 24500
rect 155900 24500 156000 24600
rect 155900 24600 156000 24700
rect 155900 24700 156000 24800
rect 155900 24800 156000 24900
rect 155900 24900 156000 25000
rect 155900 25000 156000 25100
rect 155900 25100 156000 25200
rect 155900 25200 156000 25300
rect 155900 25300 156000 25400
rect 155900 25400 156000 25500
rect 155900 25500 156000 25600
rect 155900 25600 156000 25700
rect 155900 25700 156000 25800
rect 155900 25800 156000 25900
rect 155900 25900 156000 26000
rect 155900 26000 156000 26100
rect 155900 26100 156000 26200
rect 155900 26200 156000 26300
rect 155900 26300 156000 26400
rect 155900 26400 156000 26500
rect 155900 26500 156000 26600
rect 155900 26600 156000 26700
rect 155900 26700 156000 26800
rect 155900 26800 156000 26900
rect 155900 26900 156000 27000
rect 155900 27000 156000 27100
rect 155900 27100 156000 27200
rect 155900 27200 156000 27300
rect 155900 31600 156000 31700
rect 155900 31700 156000 31800
rect 155900 31800 156000 31900
rect 155900 31900 156000 32000
rect 155900 32000 156000 32100
rect 155900 32100 156000 32200
rect 155900 32200 156000 32300
rect 155900 32300 156000 32400
rect 155900 32400 156000 32500
rect 155900 32500 156000 32600
rect 155900 32600 156000 32700
rect 155900 32700 156000 32800
rect 155900 32800 156000 32900
rect 155900 32900 156000 33000
rect 155900 33000 156000 33100
rect 155900 33100 156000 33200
rect 155900 33200 156000 33300
rect 155900 33300 156000 33400
rect 155900 33400 156000 33500
rect 155900 33500 156000 33600
rect 155900 33600 156000 33700
rect 155900 33700 156000 33800
rect 155900 33800 156000 33900
rect 155900 33900 156000 34000
rect 155900 34000 156000 34100
rect 155900 34100 156000 34200
rect 155900 34200 156000 34300
rect 155900 34300 156000 34400
rect 155900 34400 156000 34500
rect 155900 34500 156000 34600
rect 155900 34600 156000 34700
rect 155900 34700 156000 34800
rect 156000 24200 156100 24300
rect 156000 24300 156100 24400
rect 156000 24400 156100 24500
rect 156000 24500 156100 24600
rect 156000 24600 156100 24700
rect 156000 24700 156100 24800
rect 156000 24800 156100 24900
rect 156000 24900 156100 25000
rect 156000 25000 156100 25100
rect 156000 25100 156100 25200
rect 156000 25200 156100 25300
rect 156000 25300 156100 25400
rect 156000 25400 156100 25500
rect 156000 25500 156100 25600
rect 156000 25600 156100 25700
rect 156000 25700 156100 25800
rect 156000 25800 156100 25900
rect 156000 25900 156100 26000
rect 156000 26000 156100 26100
rect 156000 26100 156100 26200
rect 156000 26200 156100 26300
rect 156000 26300 156100 26400
rect 156000 26400 156100 26500
rect 156000 26500 156100 26600
rect 156000 26600 156100 26700
rect 156000 26700 156100 26800
rect 156000 26800 156100 26900
rect 156000 26900 156100 27000
rect 156000 27000 156100 27100
rect 156000 27100 156100 27200
rect 156000 31700 156100 31800
rect 156000 31800 156100 31900
rect 156000 31900 156100 32000
rect 156000 32000 156100 32100
rect 156000 32100 156100 32200
rect 156000 32200 156100 32300
rect 156000 32300 156100 32400
rect 156000 32400 156100 32500
rect 156000 32500 156100 32600
rect 156000 32600 156100 32700
rect 156000 32700 156100 32800
rect 156000 32800 156100 32900
rect 156000 32900 156100 33000
rect 156000 33000 156100 33100
rect 156000 33100 156100 33200
rect 156000 33200 156100 33300
rect 156000 33300 156100 33400
rect 156000 33400 156100 33500
rect 156000 33500 156100 33600
rect 156000 33600 156100 33700
rect 156000 33700 156100 33800
rect 156000 33800 156100 33900
rect 156000 33900 156100 34000
rect 156000 34000 156100 34100
rect 156000 34100 156100 34200
rect 156000 34200 156100 34300
rect 156000 34300 156100 34400
rect 156000 34400 156100 34500
rect 156000 34500 156100 34600
rect 156000 34600 156100 34700
rect 156000 34700 156100 34800
rect 156000 34800 156100 34900
rect 156100 24100 156200 24200
rect 156100 24200 156200 24300
rect 156100 24300 156200 24400
rect 156100 24400 156200 24500
rect 156100 24500 156200 24600
rect 156100 24600 156200 24700
rect 156100 24700 156200 24800
rect 156100 24800 156200 24900
rect 156100 24900 156200 25000
rect 156100 25000 156200 25100
rect 156100 25100 156200 25200
rect 156100 25200 156200 25300
rect 156100 25300 156200 25400
rect 156100 25400 156200 25500
rect 156100 25500 156200 25600
rect 156100 25600 156200 25700
rect 156100 25700 156200 25800
rect 156100 25800 156200 25900
rect 156100 25900 156200 26000
rect 156100 26000 156200 26100
rect 156100 26100 156200 26200
rect 156100 26200 156200 26300
rect 156100 26300 156200 26400
rect 156100 26400 156200 26500
rect 156100 26500 156200 26600
rect 156100 26600 156200 26700
rect 156100 26700 156200 26800
rect 156100 26800 156200 26900
rect 156100 26900 156200 27000
rect 156100 27000 156200 27100
rect 156100 31800 156200 31900
rect 156100 31900 156200 32000
rect 156100 32000 156200 32100
rect 156100 32100 156200 32200
rect 156100 32200 156200 32300
rect 156100 32300 156200 32400
rect 156100 32400 156200 32500
rect 156100 32500 156200 32600
rect 156100 32600 156200 32700
rect 156100 32700 156200 32800
rect 156100 32800 156200 32900
rect 156100 32900 156200 33000
rect 156100 33000 156200 33100
rect 156100 33100 156200 33200
rect 156100 33200 156200 33300
rect 156100 33300 156200 33400
rect 156100 33400 156200 33500
rect 156100 33500 156200 33600
rect 156100 33600 156200 33700
rect 156100 33700 156200 33800
rect 156100 33800 156200 33900
rect 156100 33900 156200 34000
rect 156100 34000 156200 34100
rect 156100 34100 156200 34200
rect 156100 34200 156200 34300
rect 156100 34300 156200 34400
rect 156100 34400 156200 34500
rect 156100 34500 156200 34600
rect 156100 34600 156200 34700
rect 156100 34700 156200 34800
rect 156100 34800 156200 34900
rect 156100 34900 156200 35000
rect 156200 24000 156300 24100
rect 156200 24100 156300 24200
rect 156200 24200 156300 24300
rect 156200 24300 156300 24400
rect 156200 24400 156300 24500
rect 156200 24500 156300 24600
rect 156200 24600 156300 24700
rect 156200 24700 156300 24800
rect 156200 24800 156300 24900
rect 156200 24900 156300 25000
rect 156200 25000 156300 25100
rect 156200 25100 156300 25200
rect 156200 25200 156300 25300
rect 156200 25300 156300 25400
rect 156200 25400 156300 25500
rect 156200 25500 156300 25600
rect 156200 25600 156300 25700
rect 156200 25700 156300 25800
rect 156200 25800 156300 25900
rect 156200 25900 156300 26000
rect 156200 26000 156300 26100
rect 156200 26100 156300 26200
rect 156200 26200 156300 26300
rect 156200 26300 156300 26400
rect 156200 26400 156300 26500
rect 156200 26500 156300 26600
rect 156200 26600 156300 26700
rect 156200 26700 156300 26800
rect 156200 26800 156300 26900
rect 156200 26900 156300 27000
rect 156200 31900 156300 32000
rect 156200 32000 156300 32100
rect 156200 32100 156300 32200
rect 156200 32200 156300 32300
rect 156200 32300 156300 32400
rect 156200 32400 156300 32500
rect 156200 32500 156300 32600
rect 156200 32600 156300 32700
rect 156200 32700 156300 32800
rect 156200 32800 156300 32900
rect 156200 32900 156300 33000
rect 156200 33000 156300 33100
rect 156200 33100 156300 33200
rect 156200 33200 156300 33300
rect 156200 33300 156300 33400
rect 156200 33400 156300 33500
rect 156200 33500 156300 33600
rect 156200 33600 156300 33700
rect 156200 33700 156300 33800
rect 156200 33800 156300 33900
rect 156200 33900 156300 34000
rect 156200 34000 156300 34100
rect 156200 34100 156300 34200
rect 156200 34200 156300 34300
rect 156200 34300 156300 34400
rect 156200 34400 156300 34500
rect 156200 34500 156300 34600
rect 156200 34600 156300 34700
rect 156200 34700 156300 34800
rect 156200 34800 156300 34900
rect 156200 34900 156300 35000
rect 156200 35000 156300 35100
rect 156300 23900 156400 24000
rect 156300 24000 156400 24100
rect 156300 24100 156400 24200
rect 156300 24200 156400 24300
rect 156300 24300 156400 24400
rect 156300 24400 156400 24500
rect 156300 24500 156400 24600
rect 156300 24600 156400 24700
rect 156300 24700 156400 24800
rect 156300 24800 156400 24900
rect 156300 24900 156400 25000
rect 156300 25000 156400 25100
rect 156300 25100 156400 25200
rect 156300 25200 156400 25300
rect 156300 25300 156400 25400
rect 156300 25400 156400 25500
rect 156300 25500 156400 25600
rect 156300 25600 156400 25700
rect 156300 25700 156400 25800
rect 156300 25800 156400 25900
rect 156300 25900 156400 26000
rect 156300 26000 156400 26100
rect 156300 26100 156400 26200
rect 156300 26200 156400 26300
rect 156300 26300 156400 26400
rect 156300 26400 156400 26500
rect 156300 26500 156400 26600
rect 156300 26600 156400 26700
rect 156300 26700 156400 26800
rect 156300 26800 156400 26900
rect 156300 32000 156400 32100
rect 156300 32100 156400 32200
rect 156300 32200 156400 32300
rect 156300 32300 156400 32400
rect 156300 32400 156400 32500
rect 156300 32500 156400 32600
rect 156300 32600 156400 32700
rect 156300 32700 156400 32800
rect 156300 32800 156400 32900
rect 156300 32900 156400 33000
rect 156300 33000 156400 33100
rect 156300 33100 156400 33200
rect 156300 33200 156400 33300
rect 156300 33300 156400 33400
rect 156300 33400 156400 33500
rect 156300 33500 156400 33600
rect 156300 33600 156400 33700
rect 156300 33700 156400 33800
rect 156300 33800 156400 33900
rect 156300 33900 156400 34000
rect 156300 34000 156400 34100
rect 156300 34100 156400 34200
rect 156300 34200 156400 34300
rect 156300 34300 156400 34400
rect 156300 34400 156400 34500
rect 156300 34500 156400 34600
rect 156300 34600 156400 34700
rect 156300 34700 156400 34800
rect 156300 34800 156400 34900
rect 156300 34900 156400 35000
rect 156300 35000 156400 35100
rect 156300 35100 156400 35200
rect 156400 23800 156500 23900
rect 156400 23900 156500 24000
rect 156400 24000 156500 24100
rect 156400 24100 156500 24200
rect 156400 24200 156500 24300
rect 156400 24300 156500 24400
rect 156400 24400 156500 24500
rect 156400 24500 156500 24600
rect 156400 24600 156500 24700
rect 156400 24700 156500 24800
rect 156400 24800 156500 24900
rect 156400 24900 156500 25000
rect 156400 25000 156500 25100
rect 156400 25100 156500 25200
rect 156400 25200 156500 25300
rect 156400 25300 156500 25400
rect 156400 25400 156500 25500
rect 156400 25500 156500 25600
rect 156400 25600 156500 25700
rect 156400 25700 156500 25800
rect 156400 25800 156500 25900
rect 156400 25900 156500 26000
rect 156400 26000 156500 26100
rect 156400 26100 156500 26200
rect 156400 26200 156500 26300
rect 156400 26300 156500 26400
rect 156400 26400 156500 26500
rect 156400 26500 156500 26600
rect 156400 26600 156500 26700
rect 156400 26700 156500 26800
rect 156400 32100 156500 32200
rect 156400 32200 156500 32300
rect 156400 32300 156500 32400
rect 156400 32400 156500 32500
rect 156400 32500 156500 32600
rect 156400 32600 156500 32700
rect 156400 32700 156500 32800
rect 156400 32800 156500 32900
rect 156400 32900 156500 33000
rect 156400 33000 156500 33100
rect 156400 33100 156500 33200
rect 156400 33200 156500 33300
rect 156400 33300 156500 33400
rect 156400 33400 156500 33500
rect 156400 33500 156500 33600
rect 156400 33600 156500 33700
rect 156400 33700 156500 33800
rect 156400 33800 156500 33900
rect 156400 33900 156500 34000
rect 156400 34000 156500 34100
rect 156400 34100 156500 34200
rect 156400 34200 156500 34300
rect 156400 34300 156500 34400
rect 156400 34400 156500 34500
rect 156400 34500 156500 34600
rect 156400 34600 156500 34700
rect 156400 34700 156500 34800
rect 156400 34800 156500 34900
rect 156400 34900 156500 35000
rect 156400 35000 156500 35100
rect 156400 35100 156500 35200
rect 156400 35200 156500 35300
rect 156400 35300 156500 35400
rect 156500 23700 156600 23800
rect 156500 23800 156600 23900
rect 156500 23900 156600 24000
rect 156500 24000 156600 24100
rect 156500 24100 156600 24200
rect 156500 24200 156600 24300
rect 156500 24300 156600 24400
rect 156500 24400 156600 24500
rect 156500 24500 156600 24600
rect 156500 24600 156600 24700
rect 156500 24700 156600 24800
rect 156500 24800 156600 24900
rect 156500 24900 156600 25000
rect 156500 25000 156600 25100
rect 156500 25100 156600 25200
rect 156500 25200 156600 25300
rect 156500 25300 156600 25400
rect 156500 25400 156600 25500
rect 156500 25500 156600 25600
rect 156500 25600 156600 25700
rect 156500 25700 156600 25800
rect 156500 25800 156600 25900
rect 156500 25900 156600 26000
rect 156500 26000 156600 26100
rect 156500 26100 156600 26200
rect 156500 26200 156600 26300
rect 156500 26300 156600 26400
rect 156500 26400 156600 26500
rect 156500 26500 156600 26600
rect 156500 26600 156600 26700
rect 156500 32200 156600 32300
rect 156500 32300 156600 32400
rect 156500 32400 156600 32500
rect 156500 32500 156600 32600
rect 156500 32600 156600 32700
rect 156500 32700 156600 32800
rect 156500 32800 156600 32900
rect 156500 32900 156600 33000
rect 156500 33000 156600 33100
rect 156500 33100 156600 33200
rect 156500 33200 156600 33300
rect 156500 33300 156600 33400
rect 156500 33400 156600 33500
rect 156500 33500 156600 33600
rect 156500 33600 156600 33700
rect 156500 33700 156600 33800
rect 156500 33800 156600 33900
rect 156500 33900 156600 34000
rect 156500 34000 156600 34100
rect 156500 34100 156600 34200
rect 156500 34200 156600 34300
rect 156500 34300 156600 34400
rect 156500 34400 156600 34500
rect 156500 34500 156600 34600
rect 156500 34600 156600 34700
rect 156500 34700 156600 34800
rect 156500 34800 156600 34900
rect 156500 34900 156600 35000
rect 156500 35000 156600 35100
rect 156500 35100 156600 35200
rect 156500 35200 156600 35300
rect 156500 35300 156600 35400
rect 156500 35400 156600 35500
rect 156600 23600 156700 23700
rect 156600 23700 156700 23800
rect 156600 23800 156700 23900
rect 156600 23900 156700 24000
rect 156600 24000 156700 24100
rect 156600 24100 156700 24200
rect 156600 24200 156700 24300
rect 156600 24300 156700 24400
rect 156600 24400 156700 24500
rect 156600 24500 156700 24600
rect 156600 24600 156700 24700
rect 156600 24700 156700 24800
rect 156600 24800 156700 24900
rect 156600 24900 156700 25000
rect 156600 25000 156700 25100
rect 156600 25100 156700 25200
rect 156600 25200 156700 25300
rect 156600 25300 156700 25400
rect 156600 25400 156700 25500
rect 156600 25500 156700 25600
rect 156600 25600 156700 25700
rect 156600 25700 156700 25800
rect 156600 25800 156700 25900
rect 156600 25900 156700 26000
rect 156600 26000 156700 26100
rect 156600 26100 156700 26200
rect 156600 26200 156700 26300
rect 156600 26300 156700 26400
rect 156600 26400 156700 26500
rect 156600 26500 156700 26600
rect 156600 26600 156700 26700
rect 156600 32300 156700 32400
rect 156600 32400 156700 32500
rect 156600 32500 156700 32600
rect 156600 32600 156700 32700
rect 156600 32700 156700 32800
rect 156600 32800 156700 32900
rect 156600 32900 156700 33000
rect 156600 33000 156700 33100
rect 156600 33100 156700 33200
rect 156600 33200 156700 33300
rect 156600 33300 156700 33400
rect 156600 33400 156700 33500
rect 156600 33500 156700 33600
rect 156600 33600 156700 33700
rect 156600 33700 156700 33800
rect 156600 33800 156700 33900
rect 156600 33900 156700 34000
rect 156600 34000 156700 34100
rect 156600 34100 156700 34200
rect 156600 34200 156700 34300
rect 156600 34300 156700 34400
rect 156600 34400 156700 34500
rect 156600 34500 156700 34600
rect 156600 34600 156700 34700
rect 156600 34700 156700 34800
rect 156600 34800 156700 34900
rect 156600 34900 156700 35000
rect 156600 35000 156700 35100
rect 156600 35100 156700 35200
rect 156600 35200 156700 35300
rect 156600 35300 156700 35400
rect 156600 35400 156700 35500
rect 156600 35500 156700 35600
rect 156700 23600 156800 23700
rect 156700 23700 156800 23800
rect 156700 23800 156800 23900
rect 156700 23900 156800 24000
rect 156700 24000 156800 24100
rect 156700 24100 156800 24200
rect 156700 24200 156800 24300
rect 156700 24300 156800 24400
rect 156700 24400 156800 24500
rect 156700 24500 156800 24600
rect 156700 24600 156800 24700
rect 156700 24700 156800 24800
rect 156700 24800 156800 24900
rect 156700 24900 156800 25000
rect 156700 25000 156800 25100
rect 156700 25100 156800 25200
rect 156700 25200 156800 25300
rect 156700 25300 156800 25400
rect 156700 25400 156800 25500
rect 156700 25500 156800 25600
rect 156700 25600 156800 25700
rect 156700 25700 156800 25800
rect 156700 25800 156800 25900
rect 156700 25900 156800 26000
rect 156700 26000 156800 26100
rect 156700 26100 156800 26200
rect 156700 26200 156800 26300
rect 156700 26300 156800 26400
rect 156700 26400 156800 26500
rect 156700 26500 156800 26600
rect 156700 32400 156800 32500
rect 156700 32500 156800 32600
rect 156700 32600 156800 32700
rect 156700 32700 156800 32800
rect 156700 32800 156800 32900
rect 156700 32900 156800 33000
rect 156700 33000 156800 33100
rect 156700 33100 156800 33200
rect 156700 33200 156800 33300
rect 156700 33300 156800 33400
rect 156700 33400 156800 33500
rect 156700 33500 156800 33600
rect 156700 33600 156800 33700
rect 156700 33700 156800 33800
rect 156700 33800 156800 33900
rect 156700 33900 156800 34000
rect 156700 34000 156800 34100
rect 156700 34100 156800 34200
rect 156700 34200 156800 34300
rect 156700 34300 156800 34400
rect 156700 34400 156800 34500
rect 156700 34500 156800 34600
rect 156700 34600 156800 34700
rect 156700 34700 156800 34800
rect 156700 34800 156800 34900
rect 156700 34900 156800 35000
rect 156700 35000 156800 35100
rect 156700 35100 156800 35200
rect 156700 35200 156800 35300
rect 156700 35300 156800 35400
rect 156700 35400 156800 35500
rect 156700 35500 156800 35600
rect 156700 35600 156800 35700
rect 156800 23500 156900 23600
rect 156800 23600 156900 23700
rect 156800 23700 156900 23800
rect 156800 23800 156900 23900
rect 156800 23900 156900 24000
rect 156800 24000 156900 24100
rect 156800 24100 156900 24200
rect 156800 24200 156900 24300
rect 156800 24300 156900 24400
rect 156800 24400 156900 24500
rect 156800 24500 156900 24600
rect 156800 24600 156900 24700
rect 156800 24700 156900 24800
rect 156800 24800 156900 24900
rect 156800 24900 156900 25000
rect 156800 25000 156900 25100
rect 156800 25100 156900 25200
rect 156800 25200 156900 25300
rect 156800 25300 156900 25400
rect 156800 25400 156900 25500
rect 156800 25500 156900 25600
rect 156800 25600 156900 25700
rect 156800 25700 156900 25800
rect 156800 25800 156900 25900
rect 156800 25900 156900 26000
rect 156800 26000 156900 26100
rect 156800 26100 156900 26200
rect 156800 26200 156900 26300
rect 156800 26300 156900 26400
rect 156800 26400 156900 26500
rect 156800 32500 156900 32600
rect 156800 32600 156900 32700
rect 156800 32700 156900 32800
rect 156800 32800 156900 32900
rect 156800 32900 156900 33000
rect 156800 33000 156900 33100
rect 156800 33100 156900 33200
rect 156800 33200 156900 33300
rect 156800 33300 156900 33400
rect 156800 33400 156900 33500
rect 156800 33500 156900 33600
rect 156800 33600 156900 33700
rect 156800 33700 156900 33800
rect 156800 33800 156900 33900
rect 156800 33900 156900 34000
rect 156800 34000 156900 34100
rect 156800 34100 156900 34200
rect 156800 34200 156900 34300
rect 156800 34300 156900 34400
rect 156800 34400 156900 34500
rect 156800 34500 156900 34600
rect 156800 34600 156900 34700
rect 156800 34700 156900 34800
rect 156800 34800 156900 34900
rect 156800 34900 156900 35000
rect 156800 35000 156900 35100
rect 156800 35100 156900 35200
rect 156800 35200 156900 35300
rect 156800 35300 156900 35400
rect 156800 35400 156900 35500
rect 156800 35500 156900 35600
rect 156800 35600 156900 35700
rect 156800 35700 156900 35800
rect 156900 23400 157000 23500
rect 156900 23500 157000 23600
rect 156900 23600 157000 23700
rect 156900 23700 157000 23800
rect 156900 23800 157000 23900
rect 156900 23900 157000 24000
rect 156900 24000 157000 24100
rect 156900 24100 157000 24200
rect 156900 24200 157000 24300
rect 156900 24300 157000 24400
rect 156900 24400 157000 24500
rect 156900 24500 157000 24600
rect 156900 24600 157000 24700
rect 156900 24700 157000 24800
rect 156900 24800 157000 24900
rect 156900 24900 157000 25000
rect 156900 25000 157000 25100
rect 156900 25100 157000 25200
rect 156900 25200 157000 25300
rect 156900 25300 157000 25400
rect 156900 25400 157000 25500
rect 156900 25500 157000 25600
rect 156900 25600 157000 25700
rect 156900 25700 157000 25800
rect 156900 25800 157000 25900
rect 156900 25900 157000 26000
rect 156900 26000 157000 26100
rect 156900 26100 157000 26200
rect 156900 26200 157000 26300
rect 156900 26300 157000 26400
rect 156900 32600 157000 32700
rect 156900 32700 157000 32800
rect 156900 32800 157000 32900
rect 156900 32900 157000 33000
rect 156900 33000 157000 33100
rect 156900 33100 157000 33200
rect 156900 33200 157000 33300
rect 156900 33300 157000 33400
rect 156900 33400 157000 33500
rect 156900 33500 157000 33600
rect 156900 33600 157000 33700
rect 156900 33700 157000 33800
rect 156900 33800 157000 33900
rect 156900 33900 157000 34000
rect 156900 34000 157000 34100
rect 156900 34100 157000 34200
rect 156900 34200 157000 34300
rect 156900 34300 157000 34400
rect 156900 34400 157000 34500
rect 156900 34500 157000 34600
rect 156900 34600 157000 34700
rect 156900 34700 157000 34800
rect 156900 34800 157000 34900
rect 156900 34900 157000 35000
rect 156900 35000 157000 35100
rect 156900 35100 157000 35200
rect 156900 35200 157000 35300
rect 156900 35300 157000 35400
rect 156900 35400 157000 35500
rect 156900 35500 157000 35600
rect 156900 35600 157000 35700
rect 156900 35700 157000 35800
rect 156900 35800 157000 35900
rect 157000 23300 157100 23400
rect 157000 23400 157100 23500
rect 157000 23500 157100 23600
rect 157000 23600 157100 23700
rect 157000 23700 157100 23800
rect 157000 23800 157100 23900
rect 157000 23900 157100 24000
rect 157000 24000 157100 24100
rect 157000 24100 157100 24200
rect 157000 24200 157100 24300
rect 157000 24300 157100 24400
rect 157000 24400 157100 24500
rect 157000 24500 157100 24600
rect 157000 24600 157100 24700
rect 157000 24700 157100 24800
rect 157000 24800 157100 24900
rect 157000 24900 157100 25000
rect 157000 25000 157100 25100
rect 157000 25100 157100 25200
rect 157000 25200 157100 25300
rect 157000 25300 157100 25400
rect 157000 25400 157100 25500
rect 157000 25500 157100 25600
rect 157000 25600 157100 25700
rect 157000 25700 157100 25800
rect 157000 25800 157100 25900
rect 157000 25900 157100 26000
rect 157000 26000 157100 26100
rect 157000 26100 157100 26200
rect 157000 26200 157100 26300
rect 157000 32700 157100 32800
rect 157000 32800 157100 32900
rect 157000 32900 157100 33000
rect 157000 33000 157100 33100
rect 157000 33100 157100 33200
rect 157000 33200 157100 33300
rect 157000 33300 157100 33400
rect 157000 33400 157100 33500
rect 157000 33500 157100 33600
rect 157000 33600 157100 33700
rect 157000 33700 157100 33800
rect 157000 33800 157100 33900
rect 157000 33900 157100 34000
rect 157000 34000 157100 34100
rect 157000 34100 157100 34200
rect 157000 34200 157100 34300
rect 157000 34300 157100 34400
rect 157000 34400 157100 34500
rect 157000 34500 157100 34600
rect 157000 34600 157100 34700
rect 157000 34700 157100 34800
rect 157000 34800 157100 34900
rect 157000 34900 157100 35000
rect 157000 35000 157100 35100
rect 157000 35100 157100 35200
rect 157000 35200 157100 35300
rect 157000 35300 157100 35400
rect 157000 35400 157100 35500
rect 157000 35500 157100 35600
rect 157000 35600 157100 35700
rect 157000 35700 157100 35800
rect 157000 35800 157100 35900
rect 157000 35900 157100 36000
rect 157100 23200 157200 23300
rect 157100 23300 157200 23400
rect 157100 23400 157200 23500
rect 157100 23500 157200 23600
rect 157100 23600 157200 23700
rect 157100 23700 157200 23800
rect 157100 23800 157200 23900
rect 157100 23900 157200 24000
rect 157100 24000 157200 24100
rect 157100 24100 157200 24200
rect 157100 24200 157200 24300
rect 157100 24300 157200 24400
rect 157100 24400 157200 24500
rect 157100 24500 157200 24600
rect 157100 24600 157200 24700
rect 157100 24700 157200 24800
rect 157100 24800 157200 24900
rect 157100 24900 157200 25000
rect 157100 25000 157200 25100
rect 157100 25100 157200 25200
rect 157100 25200 157200 25300
rect 157100 25300 157200 25400
rect 157100 25400 157200 25500
rect 157100 25500 157200 25600
rect 157100 25600 157200 25700
rect 157100 25700 157200 25800
rect 157100 25800 157200 25900
rect 157100 25900 157200 26000
rect 157100 26000 157200 26100
rect 157100 26100 157200 26200
rect 157100 32800 157200 32900
rect 157100 32900 157200 33000
rect 157100 33000 157200 33100
rect 157100 33100 157200 33200
rect 157100 33200 157200 33300
rect 157100 33300 157200 33400
rect 157100 33400 157200 33500
rect 157100 33500 157200 33600
rect 157100 33600 157200 33700
rect 157100 33700 157200 33800
rect 157100 33800 157200 33900
rect 157100 33900 157200 34000
rect 157100 34000 157200 34100
rect 157100 34100 157200 34200
rect 157100 34200 157200 34300
rect 157100 34300 157200 34400
rect 157100 34400 157200 34500
rect 157100 34500 157200 34600
rect 157100 34600 157200 34700
rect 157100 34700 157200 34800
rect 157100 34800 157200 34900
rect 157100 34900 157200 35000
rect 157100 35000 157200 35100
rect 157100 35100 157200 35200
rect 157100 35200 157200 35300
rect 157100 35300 157200 35400
rect 157100 35400 157200 35500
rect 157100 35500 157200 35600
rect 157100 35600 157200 35700
rect 157100 35700 157200 35800
rect 157100 35800 157200 35900
rect 157100 35900 157200 36000
rect 157100 36000 157200 36100
rect 157100 36100 157200 36200
rect 157200 23200 157300 23300
rect 157200 23300 157300 23400
rect 157200 23400 157300 23500
rect 157200 23500 157300 23600
rect 157200 23600 157300 23700
rect 157200 23700 157300 23800
rect 157200 23800 157300 23900
rect 157200 23900 157300 24000
rect 157200 24000 157300 24100
rect 157200 24100 157300 24200
rect 157200 24200 157300 24300
rect 157200 24300 157300 24400
rect 157200 24400 157300 24500
rect 157200 24500 157300 24600
rect 157200 24600 157300 24700
rect 157200 24700 157300 24800
rect 157200 24800 157300 24900
rect 157200 24900 157300 25000
rect 157200 25000 157300 25100
rect 157200 25100 157300 25200
rect 157200 25200 157300 25300
rect 157200 25300 157300 25400
rect 157200 25400 157300 25500
rect 157200 25500 157300 25600
rect 157200 25600 157300 25700
rect 157200 25700 157300 25800
rect 157200 25800 157300 25900
rect 157200 25900 157300 26000
rect 157200 26000 157300 26100
rect 157200 32900 157300 33000
rect 157200 33000 157300 33100
rect 157200 33100 157300 33200
rect 157200 33200 157300 33300
rect 157200 33300 157300 33400
rect 157200 33400 157300 33500
rect 157200 33500 157300 33600
rect 157200 33600 157300 33700
rect 157200 33700 157300 33800
rect 157200 33800 157300 33900
rect 157200 33900 157300 34000
rect 157200 34000 157300 34100
rect 157200 34100 157300 34200
rect 157200 34200 157300 34300
rect 157200 34300 157300 34400
rect 157200 34400 157300 34500
rect 157200 34500 157300 34600
rect 157200 34600 157300 34700
rect 157200 34700 157300 34800
rect 157200 34800 157300 34900
rect 157200 34900 157300 35000
rect 157200 35000 157300 35100
rect 157200 35100 157300 35200
rect 157200 35200 157300 35300
rect 157200 35300 157300 35400
rect 157200 35400 157300 35500
rect 157200 35500 157300 35600
rect 157200 35600 157300 35700
rect 157200 35700 157300 35800
rect 157200 35800 157300 35900
rect 157200 35900 157300 36000
rect 157200 36000 157300 36100
rect 157200 36100 157300 36200
rect 157200 36200 157300 36300
rect 157300 23100 157400 23200
rect 157300 23200 157400 23300
rect 157300 23300 157400 23400
rect 157300 23400 157400 23500
rect 157300 23500 157400 23600
rect 157300 23600 157400 23700
rect 157300 23700 157400 23800
rect 157300 23800 157400 23900
rect 157300 23900 157400 24000
rect 157300 24000 157400 24100
rect 157300 24100 157400 24200
rect 157300 24200 157400 24300
rect 157300 24300 157400 24400
rect 157300 24400 157400 24500
rect 157300 24500 157400 24600
rect 157300 24600 157400 24700
rect 157300 24700 157400 24800
rect 157300 24800 157400 24900
rect 157300 24900 157400 25000
rect 157300 25000 157400 25100
rect 157300 25100 157400 25200
rect 157300 25200 157400 25300
rect 157300 25300 157400 25400
rect 157300 25400 157400 25500
rect 157300 25500 157400 25600
rect 157300 25600 157400 25700
rect 157300 25700 157400 25800
rect 157300 25800 157400 25900
rect 157300 25900 157400 26000
rect 157300 33000 157400 33100
rect 157300 33100 157400 33200
rect 157300 33200 157400 33300
rect 157300 33300 157400 33400
rect 157300 33400 157400 33500
rect 157300 33500 157400 33600
rect 157300 33600 157400 33700
rect 157300 33700 157400 33800
rect 157300 33800 157400 33900
rect 157300 33900 157400 34000
rect 157300 34000 157400 34100
rect 157300 34100 157400 34200
rect 157300 34200 157400 34300
rect 157300 34300 157400 34400
rect 157300 34400 157400 34500
rect 157300 34500 157400 34600
rect 157300 34600 157400 34700
rect 157300 34700 157400 34800
rect 157300 34800 157400 34900
rect 157300 34900 157400 35000
rect 157300 35000 157400 35100
rect 157300 35100 157400 35200
rect 157300 35200 157400 35300
rect 157300 35300 157400 35400
rect 157300 35400 157400 35500
rect 157300 35500 157400 35600
rect 157300 35600 157400 35700
rect 157300 35700 157400 35800
rect 157300 35800 157400 35900
rect 157300 35900 157400 36000
rect 157300 36000 157400 36100
rect 157300 36100 157400 36200
rect 157300 36200 157400 36300
rect 157300 36300 157400 36400
rect 157400 23000 157500 23100
rect 157400 23100 157500 23200
rect 157400 23200 157500 23300
rect 157400 23300 157500 23400
rect 157400 23400 157500 23500
rect 157400 23500 157500 23600
rect 157400 23600 157500 23700
rect 157400 23700 157500 23800
rect 157400 23800 157500 23900
rect 157400 23900 157500 24000
rect 157400 24000 157500 24100
rect 157400 24100 157500 24200
rect 157400 24200 157500 24300
rect 157400 24300 157500 24400
rect 157400 24400 157500 24500
rect 157400 24500 157500 24600
rect 157400 24600 157500 24700
rect 157400 24700 157500 24800
rect 157400 24800 157500 24900
rect 157400 24900 157500 25000
rect 157400 25000 157500 25100
rect 157400 25100 157500 25200
rect 157400 25200 157500 25300
rect 157400 25300 157500 25400
rect 157400 25400 157500 25500
rect 157400 25500 157500 25600
rect 157400 25600 157500 25700
rect 157400 25700 157500 25800
rect 157400 25800 157500 25900
rect 157400 33100 157500 33200
rect 157400 33200 157500 33300
rect 157400 33300 157500 33400
rect 157400 33400 157500 33500
rect 157400 33500 157500 33600
rect 157400 33600 157500 33700
rect 157400 33700 157500 33800
rect 157400 33800 157500 33900
rect 157400 33900 157500 34000
rect 157400 34000 157500 34100
rect 157400 34100 157500 34200
rect 157400 34200 157500 34300
rect 157400 34300 157500 34400
rect 157400 34400 157500 34500
rect 157400 34500 157500 34600
rect 157400 34600 157500 34700
rect 157400 34700 157500 34800
rect 157400 34800 157500 34900
rect 157400 34900 157500 35000
rect 157400 35000 157500 35100
rect 157400 35100 157500 35200
rect 157400 35200 157500 35300
rect 157400 35300 157500 35400
rect 157400 35400 157500 35500
rect 157400 35500 157500 35600
rect 157400 35600 157500 35700
rect 157400 35700 157500 35800
rect 157400 35800 157500 35900
rect 157400 35900 157500 36000
rect 157400 36000 157500 36100
rect 157400 36100 157500 36200
rect 157400 36200 157500 36300
rect 157400 36300 157500 36400
rect 157400 36400 157500 36500
rect 157500 22900 157600 23000
rect 157500 23000 157600 23100
rect 157500 23100 157600 23200
rect 157500 23200 157600 23300
rect 157500 23300 157600 23400
rect 157500 23400 157600 23500
rect 157500 23500 157600 23600
rect 157500 23600 157600 23700
rect 157500 23700 157600 23800
rect 157500 23800 157600 23900
rect 157500 23900 157600 24000
rect 157500 24000 157600 24100
rect 157500 24100 157600 24200
rect 157500 24200 157600 24300
rect 157500 24300 157600 24400
rect 157500 24400 157600 24500
rect 157500 24500 157600 24600
rect 157500 24600 157600 24700
rect 157500 24700 157600 24800
rect 157500 24800 157600 24900
rect 157500 24900 157600 25000
rect 157500 25000 157600 25100
rect 157500 25100 157600 25200
rect 157500 25200 157600 25300
rect 157500 25300 157600 25400
rect 157500 25400 157600 25500
rect 157500 25500 157600 25600
rect 157500 25600 157600 25700
rect 157500 25700 157600 25800
rect 157500 33200 157600 33300
rect 157500 33300 157600 33400
rect 157500 33400 157600 33500
rect 157500 33500 157600 33600
rect 157500 33600 157600 33700
rect 157500 33700 157600 33800
rect 157500 33800 157600 33900
rect 157500 33900 157600 34000
rect 157500 34000 157600 34100
rect 157500 34100 157600 34200
rect 157500 34200 157600 34300
rect 157500 34300 157600 34400
rect 157500 34400 157600 34500
rect 157500 34500 157600 34600
rect 157500 34600 157600 34700
rect 157500 34700 157600 34800
rect 157500 34800 157600 34900
rect 157500 34900 157600 35000
rect 157500 35000 157600 35100
rect 157500 35100 157600 35200
rect 157500 35200 157600 35300
rect 157500 35300 157600 35400
rect 157500 35400 157600 35500
rect 157500 35500 157600 35600
rect 157500 35600 157600 35700
rect 157500 35700 157600 35800
rect 157500 35800 157600 35900
rect 157500 35900 157600 36000
rect 157500 36000 157600 36100
rect 157500 36100 157600 36200
rect 157500 36200 157600 36300
rect 157500 36300 157600 36400
rect 157500 36400 157600 36500
rect 157500 36500 157600 36600
rect 157600 22900 157700 23000
rect 157600 23000 157700 23100
rect 157600 23100 157700 23200
rect 157600 23200 157700 23300
rect 157600 23300 157700 23400
rect 157600 23400 157700 23500
rect 157600 23500 157700 23600
rect 157600 23600 157700 23700
rect 157600 23700 157700 23800
rect 157600 23800 157700 23900
rect 157600 23900 157700 24000
rect 157600 24000 157700 24100
rect 157600 24100 157700 24200
rect 157600 24200 157700 24300
rect 157600 24300 157700 24400
rect 157600 24400 157700 24500
rect 157600 24500 157700 24600
rect 157600 24600 157700 24700
rect 157600 24700 157700 24800
rect 157600 24800 157700 24900
rect 157600 24900 157700 25000
rect 157600 25000 157700 25100
rect 157600 25100 157700 25200
rect 157600 25200 157700 25300
rect 157600 25300 157700 25400
rect 157600 25400 157700 25500
rect 157600 25500 157700 25600
rect 157600 25600 157700 25700
rect 157600 33300 157700 33400
rect 157600 33400 157700 33500
rect 157600 33500 157700 33600
rect 157600 33600 157700 33700
rect 157600 33700 157700 33800
rect 157600 33800 157700 33900
rect 157600 33900 157700 34000
rect 157600 34000 157700 34100
rect 157600 34100 157700 34200
rect 157600 34200 157700 34300
rect 157600 34300 157700 34400
rect 157600 34400 157700 34500
rect 157600 34500 157700 34600
rect 157600 34600 157700 34700
rect 157600 34700 157700 34800
rect 157600 34800 157700 34900
rect 157600 34900 157700 35000
rect 157600 35000 157700 35100
rect 157600 35100 157700 35200
rect 157600 35200 157700 35300
rect 157600 35300 157700 35400
rect 157600 35400 157700 35500
rect 157600 35500 157700 35600
rect 157600 35600 157700 35700
rect 157600 35700 157700 35800
rect 157600 35800 157700 35900
rect 157600 35900 157700 36000
rect 157600 36000 157700 36100
rect 157600 36100 157700 36200
rect 157600 36200 157700 36300
rect 157600 36300 157700 36400
rect 157600 36400 157700 36500
rect 157600 36500 157700 36600
rect 157600 36600 157700 36700
rect 157700 22800 157800 22900
rect 157700 22900 157800 23000
rect 157700 23000 157800 23100
rect 157700 23100 157800 23200
rect 157700 23200 157800 23300
rect 157700 23300 157800 23400
rect 157700 23400 157800 23500
rect 157700 23500 157800 23600
rect 157700 23600 157800 23700
rect 157700 23700 157800 23800
rect 157700 23800 157800 23900
rect 157700 23900 157800 24000
rect 157700 24000 157800 24100
rect 157700 24100 157800 24200
rect 157700 24200 157800 24300
rect 157700 24300 157800 24400
rect 157700 24400 157800 24500
rect 157700 24500 157800 24600
rect 157700 24600 157800 24700
rect 157700 24700 157800 24800
rect 157700 24800 157800 24900
rect 157700 24900 157800 25000
rect 157700 25000 157800 25100
rect 157700 25100 157800 25200
rect 157700 25200 157800 25300
rect 157700 25300 157800 25400
rect 157700 25400 157800 25500
rect 157700 25500 157800 25600
rect 157700 33500 157800 33600
rect 157700 33600 157800 33700
rect 157700 33700 157800 33800
rect 157700 33800 157800 33900
rect 157700 33900 157800 34000
rect 157700 34000 157800 34100
rect 157700 34100 157800 34200
rect 157700 34200 157800 34300
rect 157700 34300 157800 34400
rect 157700 34400 157800 34500
rect 157700 34500 157800 34600
rect 157700 34600 157800 34700
rect 157700 34700 157800 34800
rect 157700 34800 157800 34900
rect 157700 34900 157800 35000
rect 157700 35000 157800 35100
rect 157700 35100 157800 35200
rect 157700 35200 157800 35300
rect 157700 35300 157800 35400
rect 157700 35400 157800 35500
rect 157700 35500 157800 35600
rect 157700 35600 157800 35700
rect 157700 35700 157800 35800
rect 157700 35800 157800 35900
rect 157700 35900 157800 36000
rect 157700 36000 157800 36100
rect 157700 36100 157800 36200
rect 157700 36200 157800 36300
rect 157700 36300 157800 36400
rect 157700 36400 157800 36500
rect 157700 36500 157800 36600
rect 157700 36600 157800 36700
rect 157700 36700 157800 36800
rect 157700 36800 157800 36900
rect 157800 22700 157900 22800
rect 157800 22800 157900 22900
rect 157800 22900 157900 23000
rect 157800 23000 157900 23100
rect 157800 23100 157900 23200
rect 157800 23200 157900 23300
rect 157800 23300 157900 23400
rect 157800 23400 157900 23500
rect 157800 23500 157900 23600
rect 157800 23600 157900 23700
rect 157800 23700 157900 23800
rect 157800 23800 157900 23900
rect 157800 23900 157900 24000
rect 157800 24000 157900 24100
rect 157800 24100 157900 24200
rect 157800 24200 157900 24300
rect 157800 24300 157900 24400
rect 157800 24400 157900 24500
rect 157800 24500 157900 24600
rect 157800 24600 157900 24700
rect 157800 24700 157900 24800
rect 157800 24800 157900 24900
rect 157800 24900 157900 25000
rect 157800 25000 157900 25100
rect 157800 25100 157900 25200
rect 157800 25200 157900 25300
rect 157800 25300 157900 25400
rect 157800 25400 157900 25500
rect 157800 33600 157900 33700
rect 157800 33700 157900 33800
rect 157800 33800 157900 33900
rect 157800 33900 157900 34000
rect 157800 34000 157900 34100
rect 157800 34100 157900 34200
rect 157800 34200 157900 34300
rect 157800 34300 157900 34400
rect 157800 34400 157900 34500
rect 157800 34500 157900 34600
rect 157800 34600 157900 34700
rect 157800 34700 157900 34800
rect 157800 34800 157900 34900
rect 157800 34900 157900 35000
rect 157800 35000 157900 35100
rect 157800 35100 157900 35200
rect 157800 35200 157900 35300
rect 157800 35300 157900 35400
rect 157800 35400 157900 35500
rect 157800 35500 157900 35600
rect 157800 35600 157900 35700
rect 157800 35700 157900 35800
rect 157800 35800 157900 35900
rect 157800 35900 157900 36000
rect 157800 36000 157900 36100
rect 157800 36100 157900 36200
rect 157800 36200 157900 36300
rect 157800 36300 157900 36400
rect 157800 36400 157900 36500
rect 157800 36500 157900 36600
rect 157800 36600 157900 36700
rect 157800 36700 157900 36800
rect 157800 36800 157900 36900
rect 157800 36900 157900 37000
rect 157900 22700 158000 22800
rect 157900 22800 158000 22900
rect 157900 22900 158000 23000
rect 157900 23000 158000 23100
rect 157900 23100 158000 23200
rect 157900 23200 158000 23300
rect 157900 23300 158000 23400
rect 157900 23400 158000 23500
rect 157900 23500 158000 23600
rect 157900 23600 158000 23700
rect 157900 23700 158000 23800
rect 157900 23800 158000 23900
rect 157900 23900 158000 24000
rect 157900 24000 158000 24100
rect 157900 24100 158000 24200
rect 157900 24200 158000 24300
rect 157900 24300 158000 24400
rect 157900 24400 158000 24500
rect 157900 24500 158000 24600
rect 157900 24600 158000 24700
rect 157900 24700 158000 24800
rect 157900 24800 158000 24900
rect 157900 24900 158000 25000
rect 157900 25000 158000 25100
rect 157900 25100 158000 25200
rect 157900 25200 158000 25300
rect 157900 25300 158000 25400
rect 157900 25400 158000 25500
rect 157900 33700 158000 33800
rect 157900 33800 158000 33900
rect 157900 33900 158000 34000
rect 157900 34000 158000 34100
rect 157900 34100 158000 34200
rect 157900 34200 158000 34300
rect 157900 34300 158000 34400
rect 157900 34400 158000 34500
rect 157900 34500 158000 34600
rect 157900 34600 158000 34700
rect 157900 34700 158000 34800
rect 157900 34800 158000 34900
rect 157900 34900 158000 35000
rect 157900 35000 158000 35100
rect 157900 35100 158000 35200
rect 157900 35200 158000 35300
rect 157900 35300 158000 35400
rect 157900 35400 158000 35500
rect 157900 35500 158000 35600
rect 157900 35600 158000 35700
rect 157900 35700 158000 35800
rect 157900 35800 158000 35900
rect 157900 35900 158000 36000
rect 157900 36000 158000 36100
rect 157900 36100 158000 36200
rect 157900 36200 158000 36300
rect 157900 36300 158000 36400
rect 157900 36400 158000 36500
rect 157900 36500 158000 36600
rect 157900 36600 158000 36700
rect 157900 36700 158000 36800
rect 157900 36800 158000 36900
rect 157900 36900 158000 37000
rect 157900 37000 158000 37100
rect 158000 22600 158100 22700
rect 158000 22700 158100 22800
rect 158000 22800 158100 22900
rect 158000 22900 158100 23000
rect 158000 23000 158100 23100
rect 158000 23100 158100 23200
rect 158000 23200 158100 23300
rect 158000 23300 158100 23400
rect 158000 23400 158100 23500
rect 158000 23500 158100 23600
rect 158000 23600 158100 23700
rect 158000 23700 158100 23800
rect 158000 23800 158100 23900
rect 158000 23900 158100 24000
rect 158000 24000 158100 24100
rect 158000 24100 158100 24200
rect 158000 24200 158100 24300
rect 158000 24300 158100 24400
rect 158000 24400 158100 24500
rect 158000 24500 158100 24600
rect 158000 24600 158100 24700
rect 158000 24700 158100 24800
rect 158000 24800 158100 24900
rect 158000 24900 158100 25000
rect 158000 25000 158100 25100
rect 158000 25100 158100 25200
rect 158000 25200 158100 25300
rect 158000 25300 158100 25400
rect 158000 33800 158100 33900
rect 158000 33900 158100 34000
rect 158000 34000 158100 34100
rect 158000 34100 158100 34200
rect 158000 34200 158100 34300
rect 158000 34300 158100 34400
rect 158000 34400 158100 34500
rect 158000 34500 158100 34600
rect 158000 34600 158100 34700
rect 158000 34700 158100 34800
rect 158000 34800 158100 34900
rect 158000 34900 158100 35000
rect 158000 35000 158100 35100
rect 158000 35100 158100 35200
rect 158000 35200 158100 35300
rect 158000 35300 158100 35400
rect 158000 35400 158100 35500
rect 158000 35500 158100 35600
rect 158000 35600 158100 35700
rect 158000 35700 158100 35800
rect 158000 35800 158100 35900
rect 158000 35900 158100 36000
rect 158000 36000 158100 36100
rect 158000 36100 158100 36200
rect 158000 36200 158100 36300
rect 158000 36300 158100 36400
rect 158000 36400 158100 36500
rect 158000 36500 158100 36600
rect 158000 36600 158100 36700
rect 158000 36700 158100 36800
rect 158000 36800 158100 36900
rect 158000 36900 158100 37000
rect 158000 37000 158100 37100
rect 158000 37100 158100 37200
rect 158100 22500 158200 22600
rect 158100 22600 158200 22700
rect 158100 22700 158200 22800
rect 158100 22800 158200 22900
rect 158100 22900 158200 23000
rect 158100 23000 158200 23100
rect 158100 23100 158200 23200
rect 158100 23200 158200 23300
rect 158100 23300 158200 23400
rect 158100 23400 158200 23500
rect 158100 23500 158200 23600
rect 158100 23600 158200 23700
rect 158100 23700 158200 23800
rect 158100 23800 158200 23900
rect 158100 23900 158200 24000
rect 158100 24000 158200 24100
rect 158100 24100 158200 24200
rect 158100 24200 158200 24300
rect 158100 24300 158200 24400
rect 158100 24400 158200 24500
rect 158100 24500 158200 24600
rect 158100 24600 158200 24700
rect 158100 24700 158200 24800
rect 158100 24800 158200 24900
rect 158100 24900 158200 25000
rect 158100 25000 158200 25100
rect 158100 25100 158200 25200
rect 158100 25200 158200 25300
rect 158100 33900 158200 34000
rect 158100 34000 158200 34100
rect 158100 34100 158200 34200
rect 158100 34200 158200 34300
rect 158100 34300 158200 34400
rect 158100 34400 158200 34500
rect 158100 34500 158200 34600
rect 158100 34600 158200 34700
rect 158100 34700 158200 34800
rect 158100 34800 158200 34900
rect 158100 34900 158200 35000
rect 158100 35000 158200 35100
rect 158100 35100 158200 35200
rect 158100 35200 158200 35300
rect 158100 35300 158200 35400
rect 158100 35400 158200 35500
rect 158100 35500 158200 35600
rect 158100 35600 158200 35700
rect 158100 35700 158200 35800
rect 158100 35800 158200 35900
rect 158100 35900 158200 36000
rect 158100 36000 158200 36100
rect 158100 36100 158200 36200
rect 158100 36200 158200 36300
rect 158100 36300 158200 36400
rect 158100 36400 158200 36500
rect 158100 36500 158200 36600
rect 158100 36600 158200 36700
rect 158100 36700 158200 36800
rect 158100 36800 158200 36900
rect 158100 36900 158200 37000
rect 158100 37000 158200 37100
rect 158100 37100 158200 37200
rect 158100 37200 158200 37300
rect 158200 22500 158300 22600
rect 158200 22600 158300 22700
rect 158200 22700 158300 22800
rect 158200 22800 158300 22900
rect 158200 22900 158300 23000
rect 158200 23000 158300 23100
rect 158200 23100 158300 23200
rect 158200 23200 158300 23300
rect 158200 23300 158300 23400
rect 158200 23400 158300 23500
rect 158200 23500 158300 23600
rect 158200 23600 158300 23700
rect 158200 23700 158300 23800
rect 158200 23800 158300 23900
rect 158200 23900 158300 24000
rect 158200 24000 158300 24100
rect 158200 24100 158300 24200
rect 158200 24200 158300 24300
rect 158200 24300 158300 24400
rect 158200 24400 158300 24500
rect 158200 24500 158300 24600
rect 158200 24600 158300 24700
rect 158200 24700 158300 24800
rect 158200 24800 158300 24900
rect 158200 24900 158300 25000
rect 158200 25000 158300 25100
rect 158200 25100 158300 25200
rect 158200 34000 158300 34100
rect 158200 34100 158300 34200
rect 158200 34200 158300 34300
rect 158200 34300 158300 34400
rect 158200 34400 158300 34500
rect 158200 34500 158300 34600
rect 158200 34600 158300 34700
rect 158200 34700 158300 34800
rect 158200 34800 158300 34900
rect 158200 34900 158300 35000
rect 158200 35000 158300 35100
rect 158200 35100 158300 35200
rect 158200 35200 158300 35300
rect 158200 35300 158300 35400
rect 158200 35400 158300 35500
rect 158200 35500 158300 35600
rect 158200 35600 158300 35700
rect 158200 35700 158300 35800
rect 158200 35800 158300 35900
rect 158200 35900 158300 36000
rect 158200 36000 158300 36100
rect 158200 36100 158300 36200
rect 158200 36200 158300 36300
rect 158200 36300 158300 36400
rect 158200 36400 158300 36500
rect 158200 36500 158300 36600
rect 158200 36600 158300 36700
rect 158200 36700 158300 36800
rect 158200 36800 158300 36900
rect 158200 36900 158300 37000
rect 158200 37000 158300 37100
rect 158200 37100 158300 37200
rect 158200 37200 158300 37300
rect 158200 37300 158300 37400
rect 158300 22400 158400 22500
rect 158300 22500 158400 22600
rect 158300 22600 158400 22700
rect 158300 22700 158400 22800
rect 158300 22800 158400 22900
rect 158300 22900 158400 23000
rect 158300 23000 158400 23100
rect 158300 23100 158400 23200
rect 158300 23200 158400 23300
rect 158300 23300 158400 23400
rect 158300 23400 158400 23500
rect 158300 23500 158400 23600
rect 158300 23600 158400 23700
rect 158300 23700 158400 23800
rect 158300 23800 158400 23900
rect 158300 23900 158400 24000
rect 158300 24000 158400 24100
rect 158300 24100 158400 24200
rect 158300 24200 158400 24300
rect 158300 24300 158400 24400
rect 158300 24400 158400 24500
rect 158300 24500 158400 24600
rect 158300 24600 158400 24700
rect 158300 24700 158400 24800
rect 158300 24800 158400 24900
rect 158300 24900 158400 25000
rect 158300 25000 158400 25100
rect 158300 34100 158400 34200
rect 158300 34200 158400 34300
rect 158300 34300 158400 34400
rect 158300 34400 158400 34500
rect 158300 34500 158400 34600
rect 158300 34600 158400 34700
rect 158300 34700 158400 34800
rect 158300 34800 158400 34900
rect 158300 34900 158400 35000
rect 158300 35000 158400 35100
rect 158300 35100 158400 35200
rect 158300 35200 158400 35300
rect 158300 35300 158400 35400
rect 158300 35400 158400 35500
rect 158300 35500 158400 35600
rect 158300 35600 158400 35700
rect 158300 35700 158400 35800
rect 158300 35800 158400 35900
rect 158300 35900 158400 36000
rect 158300 36000 158400 36100
rect 158300 36100 158400 36200
rect 158300 36200 158400 36300
rect 158300 36300 158400 36400
rect 158300 36400 158400 36500
rect 158300 36500 158400 36600
rect 158300 36600 158400 36700
rect 158300 36700 158400 36800
rect 158300 36800 158400 36900
rect 158300 36900 158400 37000
rect 158300 37000 158400 37100
rect 158300 37100 158400 37200
rect 158300 37200 158400 37300
rect 158300 37300 158400 37400
rect 158300 37400 158400 37500
rect 158300 37500 158400 37600
rect 158400 22400 158500 22500
rect 158400 22500 158500 22600
rect 158400 22600 158500 22700
rect 158400 22700 158500 22800
rect 158400 22800 158500 22900
rect 158400 22900 158500 23000
rect 158400 23000 158500 23100
rect 158400 23100 158500 23200
rect 158400 23200 158500 23300
rect 158400 23300 158500 23400
rect 158400 23400 158500 23500
rect 158400 23500 158500 23600
rect 158400 23600 158500 23700
rect 158400 23700 158500 23800
rect 158400 23800 158500 23900
rect 158400 23900 158500 24000
rect 158400 24000 158500 24100
rect 158400 24100 158500 24200
rect 158400 24200 158500 24300
rect 158400 24300 158500 24400
rect 158400 24400 158500 24500
rect 158400 24500 158500 24600
rect 158400 24600 158500 24700
rect 158400 24700 158500 24800
rect 158400 24800 158500 24900
rect 158400 24900 158500 25000
rect 158400 34300 158500 34400
rect 158400 34400 158500 34500
rect 158400 34500 158500 34600
rect 158400 34600 158500 34700
rect 158400 34700 158500 34800
rect 158400 34800 158500 34900
rect 158400 34900 158500 35000
rect 158400 35000 158500 35100
rect 158400 35100 158500 35200
rect 158400 35200 158500 35300
rect 158400 35300 158500 35400
rect 158400 35400 158500 35500
rect 158400 35500 158500 35600
rect 158400 35600 158500 35700
rect 158400 35700 158500 35800
rect 158400 35800 158500 35900
rect 158400 35900 158500 36000
rect 158400 36000 158500 36100
rect 158400 36100 158500 36200
rect 158400 36200 158500 36300
rect 158400 36300 158500 36400
rect 158400 36400 158500 36500
rect 158400 36500 158500 36600
rect 158400 36600 158500 36700
rect 158400 36700 158500 36800
rect 158400 36800 158500 36900
rect 158400 36900 158500 37000
rect 158400 37000 158500 37100
rect 158400 37100 158500 37200
rect 158400 37200 158500 37300
rect 158400 37300 158500 37400
rect 158400 37400 158500 37500
rect 158400 37500 158500 37600
rect 158400 37600 158500 37700
rect 158500 22300 158600 22400
rect 158500 22400 158600 22500
rect 158500 22500 158600 22600
rect 158500 22600 158600 22700
rect 158500 22700 158600 22800
rect 158500 22800 158600 22900
rect 158500 22900 158600 23000
rect 158500 23000 158600 23100
rect 158500 23100 158600 23200
rect 158500 23200 158600 23300
rect 158500 23300 158600 23400
rect 158500 23400 158600 23500
rect 158500 23500 158600 23600
rect 158500 23600 158600 23700
rect 158500 23700 158600 23800
rect 158500 23800 158600 23900
rect 158500 23900 158600 24000
rect 158500 24000 158600 24100
rect 158500 24100 158600 24200
rect 158500 24200 158600 24300
rect 158500 24300 158600 24400
rect 158500 24400 158600 24500
rect 158500 24500 158600 24600
rect 158500 24600 158600 24700
rect 158500 24700 158600 24800
rect 158500 24800 158600 24900
rect 158500 24900 158600 25000
rect 158500 34400 158600 34500
rect 158500 34500 158600 34600
rect 158500 34600 158600 34700
rect 158500 34700 158600 34800
rect 158500 34800 158600 34900
rect 158500 34900 158600 35000
rect 158500 35000 158600 35100
rect 158500 35100 158600 35200
rect 158500 35200 158600 35300
rect 158500 35300 158600 35400
rect 158500 35400 158600 35500
rect 158500 35500 158600 35600
rect 158500 35600 158600 35700
rect 158500 35700 158600 35800
rect 158500 35800 158600 35900
rect 158500 35900 158600 36000
rect 158500 36000 158600 36100
rect 158500 36100 158600 36200
rect 158500 36200 158600 36300
rect 158500 36300 158600 36400
rect 158500 36400 158600 36500
rect 158500 36500 158600 36600
rect 158500 36600 158600 36700
rect 158500 36700 158600 36800
rect 158500 36800 158600 36900
rect 158500 36900 158600 37000
rect 158500 37000 158600 37100
rect 158500 37100 158600 37200
rect 158500 37200 158600 37300
rect 158500 37300 158600 37400
rect 158500 37400 158600 37500
rect 158500 37500 158600 37600
rect 158500 37600 158600 37700
rect 158500 37700 158600 37800
rect 158600 22300 158700 22400
rect 158600 22400 158700 22500
rect 158600 22500 158700 22600
rect 158600 22600 158700 22700
rect 158600 22700 158700 22800
rect 158600 22800 158700 22900
rect 158600 22900 158700 23000
rect 158600 23000 158700 23100
rect 158600 23100 158700 23200
rect 158600 23200 158700 23300
rect 158600 23300 158700 23400
rect 158600 23400 158700 23500
rect 158600 23500 158700 23600
rect 158600 23600 158700 23700
rect 158600 23700 158700 23800
rect 158600 23800 158700 23900
rect 158600 23900 158700 24000
rect 158600 24000 158700 24100
rect 158600 24100 158700 24200
rect 158600 24200 158700 24300
rect 158600 24300 158700 24400
rect 158600 24400 158700 24500
rect 158600 24500 158700 24600
rect 158600 24600 158700 24700
rect 158600 24700 158700 24800
rect 158600 24800 158700 24900
rect 158600 34500 158700 34600
rect 158600 34600 158700 34700
rect 158600 34700 158700 34800
rect 158600 34800 158700 34900
rect 158600 34900 158700 35000
rect 158600 35000 158700 35100
rect 158600 35100 158700 35200
rect 158600 35200 158700 35300
rect 158600 35300 158700 35400
rect 158600 35400 158700 35500
rect 158600 35500 158700 35600
rect 158600 35600 158700 35700
rect 158600 35700 158700 35800
rect 158600 35800 158700 35900
rect 158600 35900 158700 36000
rect 158600 36000 158700 36100
rect 158600 36100 158700 36200
rect 158600 36200 158700 36300
rect 158600 36300 158700 36400
rect 158600 36400 158700 36500
rect 158600 36500 158700 36600
rect 158600 36600 158700 36700
rect 158600 36700 158700 36800
rect 158600 36800 158700 36900
rect 158600 36900 158700 37000
rect 158600 37000 158700 37100
rect 158600 37100 158700 37200
rect 158600 37200 158700 37300
rect 158600 37300 158700 37400
rect 158600 37400 158700 37500
rect 158600 37500 158700 37600
rect 158600 37600 158700 37700
rect 158600 37700 158700 37800
rect 158600 37800 158700 37900
rect 158700 22200 158800 22300
rect 158700 22300 158800 22400
rect 158700 22400 158800 22500
rect 158700 22500 158800 22600
rect 158700 22600 158800 22700
rect 158700 22700 158800 22800
rect 158700 22800 158800 22900
rect 158700 22900 158800 23000
rect 158700 23000 158800 23100
rect 158700 23100 158800 23200
rect 158700 23200 158800 23300
rect 158700 23300 158800 23400
rect 158700 23400 158800 23500
rect 158700 23500 158800 23600
rect 158700 23600 158800 23700
rect 158700 23700 158800 23800
rect 158700 23800 158800 23900
rect 158700 23900 158800 24000
rect 158700 24000 158800 24100
rect 158700 24100 158800 24200
rect 158700 24200 158800 24300
rect 158700 24300 158800 24400
rect 158700 24400 158800 24500
rect 158700 24500 158800 24600
rect 158700 24600 158800 24700
rect 158700 24700 158800 24800
rect 158700 34600 158800 34700
rect 158700 34700 158800 34800
rect 158700 34800 158800 34900
rect 158700 34900 158800 35000
rect 158700 35000 158800 35100
rect 158700 35100 158800 35200
rect 158700 35200 158800 35300
rect 158700 35300 158800 35400
rect 158700 35400 158800 35500
rect 158700 35500 158800 35600
rect 158700 35600 158800 35700
rect 158700 35700 158800 35800
rect 158700 35800 158800 35900
rect 158700 35900 158800 36000
rect 158700 36000 158800 36100
rect 158700 36100 158800 36200
rect 158700 36200 158800 36300
rect 158700 36300 158800 36400
rect 158700 36400 158800 36500
rect 158700 36500 158800 36600
rect 158700 36600 158800 36700
rect 158700 36700 158800 36800
rect 158700 36800 158800 36900
rect 158700 36900 158800 37000
rect 158700 37000 158800 37100
rect 158700 37100 158800 37200
rect 158700 37200 158800 37300
rect 158700 37300 158800 37400
rect 158700 37400 158800 37500
rect 158700 37500 158800 37600
rect 158700 37600 158800 37700
rect 158700 37700 158800 37800
rect 158700 37800 158800 37900
rect 158700 37900 158800 38000
rect 158800 22200 158900 22300
rect 158800 22300 158900 22400
rect 158800 22400 158900 22500
rect 158800 22500 158900 22600
rect 158800 22600 158900 22700
rect 158800 22700 158900 22800
rect 158800 22800 158900 22900
rect 158800 22900 158900 23000
rect 158800 23000 158900 23100
rect 158800 23100 158900 23200
rect 158800 23200 158900 23300
rect 158800 23300 158900 23400
rect 158800 23400 158900 23500
rect 158800 23500 158900 23600
rect 158800 23600 158900 23700
rect 158800 23700 158900 23800
rect 158800 23800 158900 23900
rect 158800 23900 158900 24000
rect 158800 24000 158900 24100
rect 158800 24100 158900 24200
rect 158800 24200 158900 24300
rect 158800 24300 158900 24400
rect 158800 24400 158900 24500
rect 158800 24500 158900 24600
rect 158800 24600 158900 24700
rect 158800 34700 158900 34800
rect 158800 34800 158900 34900
rect 158800 34900 158900 35000
rect 158800 35000 158900 35100
rect 158800 35100 158900 35200
rect 158800 35200 158900 35300
rect 158800 35300 158900 35400
rect 158800 35400 158900 35500
rect 158800 35500 158900 35600
rect 158800 35600 158900 35700
rect 158800 35700 158900 35800
rect 158800 35800 158900 35900
rect 158800 35900 158900 36000
rect 158800 36000 158900 36100
rect 158800 36100 158900 36200
rect 158800 36200 158900 36300
rect 158800 36300 158900 36400
rect 158800 36400 158900 36500
rect 158800 36500 158900 36600
rect 158800 36600 158900 36700
rect 158800 36700 158900 36800
rect 158800 36800 158900 36900
rect 158800 36900 158900 37000
rect 158800 37000 158900 37100
rect 158800 37100 158900 37200
rect 158800 37200 158900 37300
rect 158800 37300 158900 37400
rect 158800 37400 158900 37500
rect 158800 37500 158900 37600
rect 158800 37600 158900 37700
rect 158800 37700 158900 37800
rect 158800 37800 158900 37900
rect 158800 37900 158900 38000
rect 158900 22100 159000 22200
rect 158900 22200 159000 22300
rect 158900 22300 159000 22400
rect 158900 22400 159000 22500
rect 158900 22500 159000 22600
rect 158900 22600 159000 22700
rect 158900 22700 159000 22800
rect 158900 22800 159000 22900
rect 158900 22900 159000 23000
rect 158900 23000 159000 23100
rect 158900 23100 159000 23200
rect 158900 23200 159000 23300
rect 158900 23300 159000 23400
rect 158900 23400 159000 23500
rect 158900 23500 159000 23600
rect 158900 23600 159000 23700
rect 158900 23700 159000 23800
rect 158900 23800 159000 23900
rect 158900 23900 159000 24000
rect 158900 24000 159000 24100
rect 158900 24100 159000 24200
rect 158900 24200 159000 24300
rect 158900 24300 159000 24400
rect 158900 24400 159000 24500
rect 158900 24500 159000 24600
rect 158900 34800 159000 34900
rect 158900 34900 159000 35000
rect 158900 35000 159000 35100
rect 158900 35100 159000 35200
rect 158900 35200 159000 35300
rect 158900 35300 159000 35400
rect 158900 35400 159000 35500
rect 158900 35500 159000 35600
rect 158900 35600 159000 35700
rect 158900 35700 159000 35800
rect 158900 35800 159000 35900
rect 158900 35900 159000 36000
rect 158900 36000 159000 36100
rect 158900 36100 159000 36200
rect 158900 36200 159000 36300
rect 158900 36300 159000 36400
rect 158900 36400 159000 36500
rect 158900 36500 159000 36600
rect 158900 36600 159000 36700
rect 158900 36700 159000 36800
rect 158900 36800 159000 36900
rect 158900 36900 159000 37000
rect 158900 37000 159000 37100
rect 158900 37100 159000 37200
rect 158900 37200 159000 37300
rect 158900 37300 159000 37400
rect 158900 37400 159000 37500
rect 158900 37500 159000 37600
rect 158900 37600 159000 37700
rect 158900 37700 159000 37800
rect 158900 37800 159000 37900
rect 158900 37900 159000 38000
rect 158900 38000 159000 38100
rect 159000 22100 159100 22200
rect 159000 22200 159100 22300
rect 159000 22300 159100 22400
rect 159000 22400 159100 22500
rect 159000 22500 159100 22600
rect 159000 22600 159100 22700
rect 159000 22700 159100 22800
rect 159000 22800 159100 22900
rect 159000 22900 159100 23000
rect 159000 23000 159100 23100
rect 159000 23100 159100 23200
rect 159000 23200 159100 23300
rect 159000 23300 159100 23400
rect 159000 23400 159100 23500
rect 159000 23500 159100 23600
rect 159000 23600 159100 23700
rect 159000 23700 159100 23800
rect 159000 23800 159100 23900
rect 159000 23900 159100 24000
rect 159000 24000 159100 24100
rect 159000 24100 159100 24200
rect 159000 24200 159100 24300
rect 159000 24300 159100 24400
rect 159000 24400 159100 24500
rect 159000 24500 159100 24600
rect 159000 35000 159100 35100
rect 159000 35100 159100 35200
rect 159000 35200 159100 35300
rect 159000 35300 159100 35400
rect 159000 35400 159100 35500
rect 159000 35500 159100 35600
rect 159000 35600 159100 35700
rect 159000 35700 159100 35800
rect 159000 35800 159100 35900
rect 159000 35900 159100 36000
rect 159000 36000 159100 36100
rect 159000 36100 159100 36200
rect 159000 36200 159100 36300
rect 159000 36300 159100 36400
rect 159000 36400 159100 36500
rect 159000 36500 159100 36600
rect 159000 36600 159100 36700
rect 159000 36700 159100 36800
rect 159000 36800 159100 36900
rect 159000 36900 159100 37000
rect 159000 37000 159100 37100
rect 159000 37100 159100 37200
rect 159000 37200 159100 37300
rect 159000 37300 159100 37400
rect 159000 37400 159100 37500
rect 159000 37500 159100 37600
rect 159000 37600 159100 37700
rect 159000 37700 159100 37800
rect 159000 37800 159100 37900
rect 159000 37900 159100 38000
rect 159000 38000 159100 38100
rect 159100 22000 159200 22100
rect 159100 22100 159200 22200
rect 159100 22200 159200 22300
rect 159100 22300 159200 22400
rect 159100 22400 159200 22500
rect 159100 22500 159200 22600
rect 159100 22600 159200 22700
rect 159100 22700 159200 22800
rect 159100 22800 159200 22900
rect 159100 22900 159200 23000
rect 159100 23000 159200 23100
rect 159100 23100 159200 23200
rect 159100 23200 159200 23300
rect 159100 23300 159200 23400
rect 159100 23400 159200 23500
rect 159100 23500 159200 23600
rect 159100 23600 159200 23700
rect 159100 23700 159200 23800
rect 159100 23800 159200 23900
rect 159100 23900 159200 24000
rect 159100 24000 159200 24100
rect 159100 24100 159200 24200
rect 159100 24200 159200 24300
rect 159100 24300 159200 24400
rect 159100 24400 159200 24500
rect 159100 35100 159200 35200
rect 159100 35200 159200 35300
rect 159100 35300 159200 35400
rect 159100 35400 159200 35500
rect 159100 35500 159200 35600
rect 159100 35600 159200 35700
rect 159100 35700 159200 35800
rect 159100 35800 159200 35900
rect 159100 35900 159200 36000
rect 159100 36000 159200 36100
rect 159100 36100 159200 36200
rect 159100 36200 159200 36300
rect 159100 36300 159200 36400
rect 159100 36400 159200 36500
rect 159100 36500 159200 36600
rect 159100 36600 159200 36700
rect 159100 36700 159200 36800
rect 159100 36800 159200 36900
rect 159100 36900 159200 37000
rect 159100 37000 159200 37100
rect 159100 37100 159200 37200
rect 159100 37200 159200 37300
rect 159100 37300 159200 37400
rect 159100 37400 159200 37500
rect 159100 37500 159200 37600
rect 159100 37600 159200 37700
rect 159100 37700 159200 37800
rect 159100 37800 159200 37900
rect 159100 37900 159200 38000
rect 159100 38000 159200 38100
rect 159100 38100 159200 38200
rect 159200 22000 159300 22100
rect 159200 22100 159300 22200
rect 159200 22200 159300 22300
rect 159200 22300 159300 22400
rect 159200 22400 159300 22500
rect 159200 22500 159300 22600
rect 159200 22600 159300 22700
rect 159200 22700 159300 22800
rect 159200 22800 159300 22900
rect 159200 22900 159300 23000
rect 159200 23000 159300 23100
rect 159200 23100 159300 23200
rect 159200 23200 159300 23300
rect 159200 23300 159300 23400
rect 159200 23400 159300 23500
rect 159200 23500 159300 23600
rect 159200 23600 159300 23700
rect 159200 23700 159300 23800
rect 159200 23800 159300 23900
rect 159200 23900 159300 24000
rect 159200 24000 159300 24100
rect 159200 24100 159300 24200
rect 159200 24200 159300 24300
rect 159200 24300 159300 24400
rect 159200 35200 159300 35300
rect 159200 35300 159300 35400
rect 159200 35400 159300 35500
rect 159200 35500 159300 35600
rect 159200 35600 159300 35700
rect 159200 35700 159300 35800
rect 159200 35800 159300 35900
rect 159200 35900 159300 36000
rect 159200 36000 159300 36100
rect 159200 36100 159300 36200
rect 159200 36200 159300 36300
rect 159200 36300 159300 36400
rect 159200 36400 159300 36500
rect 159200 36500 159300 36600
rect 159200 36600 159300 36700
rect 159200 36700 159300 36800
rect 159200 36800 159300 36900
rect 159200 36900 159300 37000
rect 159200 37000 159300 37100
rect 159200 37100 159300 37200
rect 159200 37200 159300 37300
rect 159200 37300 159300 37400
rect 159200 37400 159300 37500
rect 159200 37500 159300 37600
rect 159200 37600 159300 37700
rect 159200 37700 159300 37800
rect 159200 37800 159300 37900
rect 159200 37900 159300 38000
rect 159200 38000 159300 38100
rect 159200 38100 159300 38200
rect 159300 22000 159400 22100
rect 159300 22100 159400 22200
rect 159300 22200 159400 22300
rect 159300 22300 159400 22400
rect 159300 22400 159400 22500
rect 159300 22500 159400 22600
rect 159300 22600 159400 22700
rect 159300 22700 159400 22800
rect 159300 22800 159400 22900
rect 159300 22900 159400 23000
rect 159300 23000 159400 23100
rect 159300 23100 159400 23200
rect 159300 23200 159400 23300
rect 159300 23300 159400 23400
rect 159300 23400 159400 23500
rect 159300 23500 159400 23600
rect 159300 23600 159400 23700
rect 159300 23700 159400 23800
rect 159300 23800 159400 23900
rect 159300 23900 159400 24000
rect 159300 24000 159400 24100
rect 159300 24100 159400 24200
rect 159300 24200 159400 24300
rect 159300 24300 159400 24400
rect 159300 35300 159400 35400
rect 159300 35400 159400 35500
rect 159300 35500 159400 35600
rect 159300 35600 159400 35700
rect 159300 35700 159400 35800
rect 159300 35800 159400 35900
rect 159300 35900 159400 36000
rect 159300 36000 159400 36100
rect 159300 36100 159400 36200
rect 159300 36200 159400 36300
rect 159300 36300 159400 36400
rect 159300 36400 159400 36500
rect 159300 36500 159400 36600
rect 159300 36600 159400 36700
rect 159300 36700 159400 36800
rect 159300 36800 159400 36900
rect 159300 36900 159400 37000
rect 159300 37000 159400 37100
rect 159300 37100 159400 37200
rect 159300 37200 159400 37300
rect 159300 37300 159400 37400
rect 159300 37400 159400 37500
rect 159300 37500 159400 37600
rect 159300 37600 159400 37700
rect 159300 37700 159400 37800
rect 159300 37800 159400 37900
rect 159300 37900 159400 38000
rect 159300 38000 159400 38100
rect 159300 38100 159400 38200
rect 159400 21900 159500 22000
rect 159400 22000 159500 22100
rect 159400 22100 159500 22200
rect 159400 22200 159500 22300
rect 159400 22300 159500 22400
rect 159400 22400 159500 22500
rect 159400 22500 159500 22600
rect 159400 22600 159500 22700
rect 159400 22700 159500 22800
rect 159400 22800 159500 22900
rect 159400 22900 159500 23000
rect 159400 23000 159500 23100
rect 159400 23100 159500 23200
rect 159400 23200 159500 23300
rect 159400 23300 159500 23400
rect 159400 23400 159500 23500
rect 159400 23500 159500 23600
rect 159400 23600 159500 23700
rect 159400 23700 159500 23800
rect 159400 23800 159500 23900
rect 159400 23900 159500 24000
rect 159400 24000 159500 24100
rect 159400 24100 159500 24200
rect 159400 24200 159500 24300
rect 159400 35500 159500 35600
rect 159400 35600 159500 35700
rect 159400 35700 159500 35800
rect 159400 35800 159500 35900
rect 159400 35900 159500 36000
rect 159400 36000 159500 36100
rect 159400 36100 159500 36200
rect 159400 36200 159500 36300
rect 159400 36300 159500 36400
rect 159400 36400 159500 36500
rect 159400 36500 159500 36600
rect 159400 36600 159500 36700
rect 159400 36700 159500 36800
rect 159400 36800 159500 36900
rect 159400 36900 159500 37000
rect 159400 37000 159500 37100
rect 159400 37100 159500 37200
rect 159400 37200 159500 37300
rect 159400 37300 159500 37400
rect 159400 37400 159500 37500
rect 159400 37500 159500 37600
rect 159400 37600 159500 37700
rect 159400 37700 159500 37800
rect 159400 37800 159500 37900
rect 159400 37900 159500 38000
rect 159400 38000 159500 38100
rect 159400 38100 159500 38200
rect 159500 21900 159600 22000
rect 159500 22000 159600 22100
rect 159500 22100 159600 22200
rect 159500 22200 159600 22300
rect 159500 22300 159600 22400
rect 159500 22400 159600 22500
rect 159500 22500 159600 22600
rect 159500 22600 159600 22700
rect 159500 22700 159600 22800
rect 159500 22800 159600 22900
rect 159500 22900 159600 23000
rect 159500 23000 159600 23100
rect 159500 23100 159600 23200
rect 159500 23200 159600 23300
rect 159500 23300 159600 23400
rect 159500 23400 159600 23500
rect 159500 23500 159600 23600
rect 159500 23600 159600 23700
rect 159500 23700 159600 23800
rect 159500 23800 159600 23900
rect 159500 23900 159600 24000
rect 159500 24000 159600 24100
rect 159500 24100 159600 24200
rect 159500 24200 159600 24300
rect 159500 35600 159600 35700
rect 159500 35700 159600 35800
rect 159500 35800 159600 35900
rect 159500 35900 159600 36000
rect 159500 36000 159600 36100
rect 159500 36100 159600 36200
rect 159500 36200 159600 36300
rect 159500 36300 159600 36400
rect 159500 36400 159600 36500
rect 159500 36500 159600 36600
rect 159500 36600 159600 36700
rect 159500 36700 159600 36800
rect 159500 36800 159600 36900
rect 159500 36900 159600 37000
rect 159500 37000 159600 37100
rect 159500 37100 159600 37200
rect 159500 37200 159600 37300
rect 159500 37300 159600 37400
rect 159500 37400 159600 37500
rect 159500 37500 159600 37600
rect 159500 37600 159600 37700
rect 159500 37700 159600 37800
rect 159500 37800 159600 37900
rect 159500 37900 159600 38000
rect 159500 38000 159600 38100
rect 159600 21900 159700 22000
rect 159600 22000 159700 22100
rect 159600 22100 159700 22200
rect 159600 22200 159700 22300
rect 159600 22300 159700 22400
rect 159600 22400 159700 22500
rect 159600 22500 159700 22600
rect 159600 22600 159700 22700
rect 159600 22700 159700 22800
rect 159600 22800 159700 22900
rect 159600 22900 159700 23000
rect 159600 23000 159700 23100
rect 159600 23100 159700 23200
rect 159600 23200 159700 23300
rect 159600 23300 159700 23400
rect 159600 23400 159700 23500
rect 159600 23500 159700 23600
rect 159600 23600 159700 23700
rect 159600 23700 159700 23800
rect 159600 23800 159700 23900
rect 159600 23900 159700 24000
rect 159600 24000 159700 24100
rect 159600 24100 159700 24200
rect 159600 35700 159700 35800
rect 159600 35800 159700 35900
rect 159600 35900 159700 36000
rect 159600 36000 159700 36100
rect 159600 36100 159700 36200
rect 159600 36200 159700 36300
rect 159600 36300 159700 36400
rect 159600 36400 159700 36500
rect 159600 36500 159700 36600
rect 159600 36600 159700 36700
rect 159600 36700 159700 36800
rect 159600 36800 159700 36900
rect 159600 36900 159700 37000
rect 159600 37000 159700 37100
rect 159600 37100 159700 37200
rect 159600 37200 159700 37300
rect 159600 37300 159700 37400
rect 159600 37400 159700 37500
rect 159600 37500 159700 37600
rect 159600 37600 159700 37700
rect 159600 37700 159700 37800
rect 159600 37800 159700 37900
rect 159600 37900 159700 38000
rect 159600 38000 159700 38100
rect 159700 21900 159800 22000
rect 159700 22000 159800 22100
rect 159700 22100 159800 22200
rect 159700 22200 159800 22300
rect 159700 22300 159800 22400
rect 159700 22400 159800 22500
rect 159700 22500 159800 22600
rect 159700 22600 159800 22700
rect 159700 22700 159800 22800
rect 159700 22800 159800 22900
rect 159700 22900 159800 23000
rect 159700 23000 159800 23100
rect 159700 23100 159800 23200
rect 159700 23200 159800 23300
rect 159700 23300 159800 23400
rect 159700 23400 159800 23500
rect 159700 23500 159800 23600
rect 159700 23600 159800 23700
rect 159700 23700 159800 23800
rect 159700 23800 159800 23900
rect 159700 23900 159800 24000
rect 159700 24000 159800 24100
rect 159700 24100 159800 24200
rect 159700 35900 159800 36000
rect 159700 36000 159800 36100
rect 159700 36100 159800 36200
rect 159700 36200 159800 36300
rect 159700 36300 159800 36400
rect 159700 36400 159800 36500
rect 159700 36500 159800 36600
rect 159700 36600 159800 36700
rect 159700 36700 159800 36800
rect 159700 36800 159800 36900
rect 159700 36900 159800 37000
rect 159700 37000 159800 37100
rect 159700 37100 159800 37200
rect 159700 37200 159800 37300
rect 159700 37300 159800 37400
rect 159700 37400 159800 37500
rect 159700 37500 159800 37600
rect 159700 37600 159800 37700
rect 159700 37700 159800 37800
rect 159700 37800 159800 37900
rect 159700 37900 159800 38000
rect 159700 38000 159800 38100
rect 159800 21900 159900 22000
rect 159800 22000 159900 22100
rect 159800 22100 159900 22200
rect 159800 22200 159900 22300
rect 159800 22300 159900 22400
rect 159800 22400 159900 22500
rect 159800 22500 159900 22600
rect 159800 22600 159900 22700
rect 159800 22700 159900 22800
rect 159800 22800 159900 22900
rect 159800 22900 159900 23000
rect 159800 23000 159900 23100
rect 159800 23100 159900 23200
rect 159800 23200 159900 23300
rect 159800 23300 159900 23400
rect 159800 23400 159900 23500
rect 159800 23500 159900 23600
rect 159800 23600 159900 23700
rect 159800 23700 159900 23800
rect 159800 23800 159900 23900
rect 159800 23900 159900 24000
rect 159800 24000 159900 24100
rect 159800 36000 159900 36100
rect 159800 36100 159900 36200
rect 159800 36200 159900 36300
rect 159800 36300 159900 36400
rect 159800 36400 159900 36500
rect 159800 36500 159900 36600
rect 159800 36600 159900 36700
rect 159800 36700 159900 36800
rect 159800 36800 159900 36900
rect 159800 36900 159900 37000
rect 159800 37000 159900 37100
rect 159800 37100 159900 37200
rect 159800 37200 159900 37300
rect 159800 37300 159900 37400
rect 159800 37400 159900 37500
rect 159800 37500 159900 37600
rect 159800 37600 159900 37700
rect 159800 37700 159900 37800
rect 159800 37800 159900 37900
rect 159800 37900 159900 38000
rect 159900 21900 160000 22000
rect 159900 22000 160000 22100
rect 159900 22100 160000 22200
rect 159900 22200 160000 22300
rect 159900 22300 160000 22400
rect 159900 22400 160000 22500
rect 159900 22500 160000 22600
rect 159900 22600 160000 22700
rect 159900 22700 160000 22800
rect 159900 22800 160000 22900
rect 159900 22900 160000 23000
rect 159900 23000 160000 23100
rect 159900 23100 160000 23200
rect 159900 23200 160000 23300
rect 159900 23300 160000 23400
rect 159900 23400 160000 23500
rect 159900 23500 160000 23600
rect 159900 23600 160000 23700
rect 159900 23700 160000 23800
rect 159900 23800 160000 23900
rect 159900 23900 160000 24000
rect 159900 24000 160000 24100
rect 159900 36100 160000 36200
rect 159900 36200 160000 36300
rect 159900 36300 160000 36400
rect 159900 36400 160000 36500
rect 159900 36500 160000 36600
rect 159900 36600 160000 36700
rect 159900 36700 160000 36800
rect 159900 36800 160000 36900
rect 159900 36900 160000 37000
rect 159900 37000 160000 37100
rect 159900 37100 160000 37200
rect 159900 37200 160000 37300
rect 159900 37300 160000 37400
rect 159900 37400 160000 37500
rect 159900 37500 160000 37600
rect 159900 37600 160000 37700
rect 159900 37700 160000 37800
rect 159900 37800 160000 37900
rect 159900 37900 160000 38000
rect 160000 21900 160100 22000
rect 160000 22000 160100 22100
rect 160000 22100 160100 22200
rect 160000 22200 160100 22300
rect 160000 22300 160100 22400
rect 160000 22400 160100 22500
rect 160000 22500 160100 22600
rect 160000 22600 160100 22700
rect 160000 22700 160100 22800
rect 160000 22800 160100 22900
rect 160000 22900 160100 23000
rect 160000 23000 160100 23100
rect 160000 23100 160100 23200
rect 160000 23200 160100 23300
rect 160000 23300 160100 23400
rect 160000 23400 160100 23500
rect 160000 23500 160100 23600
rect 160000 23600 160100 23700
rect 160000 23700 160100 23800
rect 160000 23800 160100 23900
rect 160000 23900 160100 24000
rect 160000 36300 160100 36400
rect 160000 36400 160100 36500
rect 160000 36500 160100 36600
rect 160000 36600 160100 36700
rect 160000 36700 160100 36800
rect 160000 36800 160100 36900
rect 160000 36900 160100 37000
rect 160000 37000 160100 37100
rect 160000 37100 160100 37200
rect 160000 37200 160100 37300
rect 160000 37300 160100 37400
rect 160000 37400 160100 37500
rect 160000 37500 160100 37600
rect 160000 37600 160100 37700
rect 160000 37700 160100 37800
rect 160000 37800 160100 37900
rect 160100 21900 160200 22000
rect 160100 22000 160200 22100
rect 160100 22100 160200 22200
rect 160100 22200 160200 22300
rect 160100 22300 160200 22400
rect 160100 22400 160200 22500
rect 160100 22500 160200 22600
rect 160100 22600 160200 22700
rect 160100 22700 160200 22800
rect 160100 22800 160200 22900
rect 160100 22900 160200 23000
rect 160100 23000 160200 23100
rect 160100 23100 160200 23200
rect 160100 23200 160200 23300
rect 160100 23300 160200 23400
rect 160100 23400 160200 23500
rect 160100 23500 160200 23600
rect 160100 23600 160200 23700
rect 160100 23700 160200 23800
rect 160100 23800 160200 23900
rect 160100 23900 160200 24000
rect 160100 36500 160200 36600
rect 160100 36600 160200 36700
rect 160100 36700 160200 36800
rect 160100 36800 160200 36900
rect 160100 36900 160200 37000
rect 160100 37000 160200 37100
rect 160100 37100 160200 37200
rect 160100 37200 160200 37300
rect 160100 37300 160200 37400
rect 160100 37400 160200 37500
rect 160100 37500 160200 37600
rect 160100 37600 160200 37700
rect 160100 37700 160200 37800
rect 160200 21900 160300 22000
rect 160200 22000 160300 22100
rect 160200 22100 160300 22200
rect 160200 22200 160300 22300
rect 160200 22300 160300 22400
rect 160200 22400 160300 22500
rect 160200 22500 160300 22600
rect 160200 22600 160300 22700
rect 160200 22700 160300 22800
rect 160200 22800 160300 22900
rect 160200 22900 160300 23000
rect 160200 23000 160300 23100
rect 160200 23100 160300 23200
rect 160200 23200 160300 23300
rect 160200 23300 160300 23400
rect 160200 23400 160300 23500
rect 160200 23500 160300 23600
rect 160200 23600 160300 23700
rect 160200 23700 160300 23800
rect 160200 23800 160300 23900
rect 160200 23900 160300 24000
rect 160200 36600 160300 36700
rect 160200 36700 160300 36800
rect 160200 36800 160300 36900
rect 160200 36900 160300 37000
rect 160200 37000 160300 37100
rect 160200 37100 160300 37200
rect 160200 37200 160300 37300
rect 160200 37300 160300 37400
rect 160200 37400 160300 37500
rect 160200 37500 160300 37600
rect 160300 21900 160400 22000
rect 160300 22000 160400 22100
rect 160300 22100 160400 22200
rect 160300 22200 160400 22300
rect 160300 22300 160400 22400
rect 160300 22400 160400 22500
rect 160300 22500 160400 22600
rect 160300 22600 160400 22700
rect 160300 22700 160400 22800
rect 160300 22800 160400 22900
rect 160300 22900 160400 23000
rect 160300 23000 160400 23100
rect 160300 23100 160400 23200
rect 160300 23200 160400 23300
rect 160300 23300 160400 23400
rect 160300 23400 160400 23500
rect 160300 23500 160400 23600
rect 160300 23600 160400 23700
rect 160300 23700 160400 23800
rect 160300 23800 160400 23900
rect 160300 36900 160400 37000
rect 160300 37000 160400 37100
rect 160300 37100 160400 37200
rect 160300 37200 160400 37300
rect 160300 37300 160400 37400
rect 160400 22000 160500 22100
rect 160400 22100 160500 22200
rect 160400 22200 160500 22300
rect 160400 22300 160500 22400
rect 160400 22400 160500 22500
rect 160400 22500 160500 22600
rect 160400 22600 160500 22700
rect 160400 22700 160500 22800
rect 160400 22800 160500 22900
rect 160400 22900 160500 23000
rect 160400 23000 160500 23100
rect 160400 23100 160500 23200
rect 160400 23200 160500 23300
rect 160400 23300 160500 23400
rect 160400 23400 160500 23500
rect 160400 23500 160500 23600
rect 160400 23600 160500 23700
rect 160400 23700 160500 23800
rect 160400 23800 160500 23900
rect 160500 22000 160600 22100
rect 160500 22100 160600 22200
rect 160500 22200 160600 22300
rect 160500 22300 160600 22400
rect 160500 22400 160600 22500
rect 160500 22500 160600 22600
rect 160500 22600 160600 22700
rect 160500 22700 160600 22800
rect 160500 22800 160600 22900
rect 160500 22900 160600 23000
rect 160500 23000 160600 23100
rect 160500 23100 160600 23200
rect 160500 23200 160600 23300
rect 160500 23300 160600 23400
rect 160500 23400 160600 23500
rect 160500 23500 160600 23600
rect 160500 23600 160600 23700
rect 160500 23700 160600 23800
rect 160600 22100 160700 22200
rect 160600 22200 160700 22300
rect 160600 22300 160700 22400
rect 160600 22400 160700 22500
rect 160600 22500 160700 22600
rect 160600 22600 160700 22700
rect 160600 22700 160700 22800
rect 160600 22800 160700 22900
rect 160600 22900 160700 23000
rect 160600 23000 160700 23100
rect 160600 23100 160700 23200
rect 160600 23200 160700 23300
rect 160600 23300 160700 23400
rect 160600 23400 160700 23500
rect 160600 23500 160700 23600
rect 160600 23600 160700 23700
rect 160700 22200 160800 22300
rect 160700 22300 160800 22400
rect 160700 22400 160800 22500
rect 160700 22500 160800 22600
rect 160700 22600 160800 22700
rect 160700 22700 160800 22800
rect 160700 22800 160800 22900
rect 160700 22900 160800 23000
rect 160700 23000 160800 23100
rect 160700 23100 160800 23200
rect 160700 23200 160800 23300
rect 160700 23300 160800 23400
rect 160700 23400 160800 23500
rect 160700 23500 160800 23600
rect 160800 22400 160900 22500
rect 160800 22500 160900 22600
rect 160800 22600 160900 22700
rect 160800 22700 160900 22800
rect 160800 22800 160900 22900
rect 160800 22900 160900 23000
rect 160800 23000 160900 23100
rect 160800 23100 160900 23200
rect 160800 23200 160900 23300
rect 160800 23300 160900 23400
rect 160800 23400 160900 23500
rect 160900 22600 161000 22700
rect 160900 22700 161000 22800
rect 160900 22800 161000 22900
rect 160900 22900 161000 23000
rect 160900 23000 161000 23100
rect 160900 23100 161000 23200
rect 160900 23200 161000 23300
rect 162500 37200 162600 37300
rect 162500 37400 162600 37500
rect 162600 36800 162700 36900
rect 162600 36900 162700 37000
rect 162600 37000 162700 37100
rect 162600 37100 162700 37200
rect 162600 37200 162700 37300
rect 162600 37300 162700 37400
rect 162600 37400 162700 37500
rect 162600 37500 162700 37600
rect 162600 37600 162700 37700
rect 162600 37700 162700 37800
rect 162700 36500 162800 36600
rect 162700 36600 162800 36700
rect 162700 36700 162800 36800
rect 162700 36800 162800 36900
rect 162700 36900 162800 37000
rect 162700 37000 162800 37100
rect 162700 37100 162800 37200
rect 162700 37200 162800 37300
rect 162700 37300 162800 37400
rect 162700 37400 162800 37500
rect 162700 37500 162800 37600
rect 162700 37600 162800 37700
rect 162700 37700 162800 37800
rect 162700 37800 162800 37900
rect 162700 37900 162800 38000
rect 162800 36200 162900 36300
rect 162800 36300 162900 36400
rect 162800 36400 162900 36500
rect 162800 36500 162900 36600
rect 162800 36600 162900 36700
rect 162800 36700 162900 36800
rect 162800 36800 162900 36900
rect 162800 36900 162900 37000
rect 162800 37000 162900 37100
rect 162800 37100 162900 37200
rect 162800 37200 162900 37300
rect 162800 37300 162900 37400
rect 162800 37400 162900 37500
rect 162800 37500 162900 37600
rect 162800 37600 162900 37700
rect 162800 37700 162900 37800
rect 162800 37800 162900 37900
rect 162800 37900 162900 38000
rect 162800 38000 162900 38100
rect 162900 35900 163000 36000
rect 162900 36000 163000 36100
rect 162900 36100 163000 36200
rect 162900 36200 163000 36300
rect 162900 36300 163000 36400
rect 162900 36400 163000 36500
rect 162900 36500 163000 36600
rect 162900 36600 163000 36700
rect 162900 36700 163000 36800
rect 162900 36800 163000 36900
rect 162900 36900 163000 37000
rect 162900 37000 163000 37100
rect 162900 37100 163000 37200
rect 162900 37200 163000 37300
rect 162900 37300 163000 37400
rect 162900 37400 163000 37500
rect 162900 37500 163000 37600
rect 162900 37600 163000 37700
rect 162900 37700 163000 37800
rect 162900 37800 163000 37900
rect 162900 37900 163000 38000
rect 162900 38000 163000 38100
rect 163000 35600 163100 35700
rect 163000 35700 163100 35800
rect 163000 35800 163100 35900
rect 163000 35900 163100 36000
rect 163000 36000 163100 36100
rect 163000 36100 163100 36200
rect 163000 36200 163100 36300
rect 163000 36300 163100 36400
rect 163000 36400 163100 36500
rect 163000 36500 163100 36600
rect 163000 36600 163100 36700
rect 163000 36700 163100 36800
rect 163000 36800 163100 36900
rect 163000 36900 163100 37000
rect 163000 37000 163100 37100
rect 163000 37100 163100 37200
rect 163000 37200 163100 37300
rect 163000 37300 163100 37400
rect 163000 37400 163100 37500
rect 163000 37500 163100 37600
rect 163000 37600 163100 37700
rect 163000 37700 163100 37800
rect 163000 37800 163100 37900
rect 163000 37900 163100 38000
rect 163000 38000 163100 38100
rect 163000 38100 163100 38200
rect 163100 35300 163200 35400
rect 163100 35400 163200 35500
rect 163100 35500 163200 35600
rect 163100 35600 163200 35700
rect 163100 35700 163200 35800
rect 163100 35800 163200 35900
rect 163100 35900 163200 36000
rect 163100 36000 163200 36100
rect 163100 36100 163200 36200
rect 163100 36200 163200 36300
rect 163100 36300 163200 36400
rect 163100 36400 163200 36500
rect 163100 36500 163200 36600
rect 163100 36600 163200 36700
rect 163100 36700 163200 36800
rect 163100 36800 163200 36900
rect 163100 36900 163200 37000
rect 163100 37000 163200 37100
rect 163100 37100 163200 37200
rect 163100 37200 163200 37300
rect 163100 37300 163200 37400
rect 163100 37400 163200 37500
rect 163100 37500 163200 37600
rect 163100 37600 163200 37700
rect 163100 37700 163200 37800
rect 163100 37800 163200 37900
rect 163100 37900 163200 38000
rect 163100 38000 163200 38100
rect 163100 38100 163200 38200
rect 163200 35000 163300 35100
rect 163200 35100 163300 35200
rect 163200 35200 163300 35300
rect 163200 35300 163300 35400
rect 163200 35400 163300 35500
rect 163200 35500 163300 35600
rect 163200 35600 163300 35700
rect 163200 35700 163300 35800
rect 163200 35800 163300 35900
rect 163200 35900 163300 36000
rect 163200 36000 163300 36100
rect 163200 36100 163300 36200
rect 163200 36200 163300 36300
rect 163200 36300 163300 36400
rect 163200 36400 163300 36500
rect 163200 36500 163300 36600
rect 163200 36600 163300 36700
rect 163200 36700 163300 36800
rect 163200 36800 163300 36900
rect 163200 36900 163300 37000
rect 163200 37000 163300 37100
rect 163200 37100 163300 37200
rect 163200 37200 163300 37300
rect 163200 37300 163300 37400
rect 163200 37400 163300 37500
rect 163200 37500 163300 37600
rect 163200 37600 163300 37700
rect 163200 37700 163300 37800
rect 163200 37800 163300 37900
rect 163200 37900 163300 38000
rect 163200 38000 163300 38100
rect 163200 38100 163300 38200
rect 163200 38200 163300 38300
rect 163300 34700 163400 34800
rect 163300 34800 163400 34900
rect 163300 34900 163400 35000
rect 163300 35000 163400 35100
rect 163300 35100 163400 35200
rect 163300 35200 163400 35300
rect 163300 35300 163400 35400
rect 163300 35400 163400 35500
rect 163300 35500 163400 35600
rect 163300 35600 163400 35700
rect 163300 35700 163400 35800
rect 163300 35800 163400 35900
rect 163300 35900 163400 36000
rect 163300 36000 163400 36100
rect 163300 36100 163400 36200
rect 163300 36200 163400 36300
rect 163300 36300 163400 36400
rect 163300 36400 163400 36500
rect 163300 36500 163400 36600
rect 163300 36600 163400 36700
rect 163300 36700 163400 36800
rect 163300 36800 163400 36900
rect 163300 36900 163400 37000
rect 163300 37000 163400 37100
rect 163300 37100 163400 37200
rect 163300 37200 163400 37300
rect 163300 37300 163400 37400
rect 163300 37400 163400 37500
rect 163300 37500 163400 37600
rect 163300 37600 163400 37700
rect 163300 37700 163400 37800
rect 163300 37800 163400 37900
rect 163300 37900 163400 38000
rect 163300 38000 163400 38100
rect 163300 38100 163400 38200
rect 163300 38200 163400 38300
rect 163400 34400 163500 34500
rect 163400 34500 163500 34600
rect 163400 34600 163500 34700
rect 163400 34700 163500 34800
rect 163400 34800 163500 34900
rect 163400 34900 163500 35000
rect 163400 35000 163500 35100
rect 163400 35100 163500 35200
rect 163400 35200 163500 35300
rect 163400 35300 163500 35400
rect 163400 35400 163500 35500
rect 163400 35500 163500 35600
rect 163400 35600 163500 35700
rect 163400 35700 163500 35800
rect 163400 35800 163500 35900
rect 163400 35900 163500 36000
rect 163400 36000 163500 36100
rect 163400 36100 163500 36200
rect 163400 36200 163500 36300
rect 163400 36300 163500 36400
rect 163400 36400 163500 36500
rect 163400 36500 163500 36600
rect 163400 36600 163500 36700
rect 163400 36700 163500 36800
rect 163400 36800 163500 36900
rect 163400 36900 163500 37000
rect 163400 37000 163500 37100
rect 163400 37100 163500 37200
rect 163400 37200 163500 37300
rect 163400 37300 163500 37400
rect 163400 37400 163500 37500
rect 163400 37500 163500 37600
rect 163400 37600 163500 37700
rect 163400 37700 163500 37800
rect 163400 37800 163500 37900
rect 163400 37900 163500 38000
rect 163400 38000 163500 38100
rect 163400 38100 163500 38200
rect 163400 38200 163500 38300
rect 163500 34100 163600 34200
rect 163500 34200 163600 34300
rect 163500 34300 163600 34400
rect 163500 34400 163600 34500
rect 163500 34500 163600 34600
rect 163500 34600 163600 34700
rect 163500 34700 163600 34800
rect 163500 34800 163600 34900
rect 163500 34900 163600 35000
rect 163500 35000 163600 35100
rect 163500 35100 163600 35200
rect 163500 35200 163600 35300
rect 163500 35300 163600 35400
rect 163500 35400 163600 35500
rect 163500 35500 163600 35600
rect 163500 35600 163600 35700
rect 163500 35700 163600 35800
rect 163500 35800 163600 35900
rect 163500 35900 163600 36000
rect 163500 36000 163600 36100
rect 163500 36100 163600 36200
rect 163500 36200 163600 36300
rect 163500 36300 163600 36400
rect 163500 36400 163600 36500
rect 163500 36500 163600 36600
rect 163500 36600 163600 36700
rect 163500 36700 163600 36800
rect 163500 36800 163600 36900
rect 163500 36900 163600 37000
rect 163500 37000 163600 37100
rect 163500 37100 163600 37200
rect 163500 37200 163600 37300
rect 163500 37300 163600 37400
rect 163500 37400 163600 37500
rect 163500 37500 163600 37600
rect 163500 37600 163600 37700
rect 163500 37700 163600 37800
rect 163500 37800 163600 37900
rect 163500 37900 163600 38000
rect 163500 38000 163600 38100
rect 163500 38100 163600 38200
rect 163500 38200 163600 38300
rect 163600 33800 163700 33900
rect 163600 33900 163700 34000
rect 163600 34000 163700 34100
rect 163600 34100 163700 34200
rect 163600 34200 163700 34300
rect 163600 34300 163700 34400
rect 163600 34400 163700 34500
rect 163600 34500 163700 34600
rect 163600 34600 163700 34700
rect 163600 34700 163700 34800
rect 163600 34800 163700 34900
rect 163600 34900 163700 35000
rect 163600 35000 163700 35100
rect 163600 35100 163700 35200
rect 163600 35200 163700 35300
rect 163600 35300 163700 35400
rect 163600 35400 163700 35500
rect 163600 35500 163700 35600
rect 163600 35600 163700 35700
rect 163600 35700 163700 35800
rect 163600 35800 163700 35900
rect 163600 35900 163700 36000
rect 163600 36000 163700 36100
rect 163600 36100 163700 36200
rect 163600 36200 163700 36300
rect 163600 36300 163700 36400
rect 163600 36400 163700 36500
rect 163600 36500 163700 36600
rect 163600 36600 163700 36700
rect 163600 36700 163700 36800
rect 163600 36800 163700 36900
rect 163600 36900 163700 37000
rect 163600 37000 163700 37100
rect 163600 37100 163700 37200
rect 163600 37200 163700 37300
rect 163600 37300 163700 37400
rect 163600 37400 163700 37500
rect 163600 37500 163700 37600
rect 163600 37600 163700 37700
rect 163600 37700 163700 37800
rect 163600 37800 163700 37900
rect 163600 37900 163700 38000
rect 163600 38000 163700 38100
rect 163600 38100 163700 38200
rect 163600 38200 163700 38300
rect 163700 33500 163800 33600
rect 163700 33600 163800 33700
rect 163700 33700 163800 33800
rect 163700 33800 163800 33900
rect 163700 33900 163800 34000
rect 163700 34000 163800 34100
rect 163700 34100 163800 34200
rect 163700 34200 163800 34300
rect 163700 34300 163800 34400
rect 163700 34400 163800 34500
rect 163700 34500 163800 34600
rect 163700 34600 163800 34700
rect 163700 34700 163800 34800
rect 163700 34800 163800 34900
rect 163700 34900 163800 35000
rect 163700 35000 163800 35100
rect 163700 35100 163800 35200
rect 163700 35200 163800 35300
rect 163700 35300 163800 35400
rect 163700 35400 163800 35500
rect 163700 35500 163800 35600
rect 163700 35600 163800 35700
rect 163700 35700 163800 35800
rect 163700 35800 163800 35900
rect 163700 35900 163800 36000
rect 163700 36000 163800 36100
rect 163700 36100 163800 36200
rect 163700 36200 163800 36300
rect 163700 36300 163800 36400
rect 163700 36400 163800 36500
rect 163700 36500 163800 36600
rect 163700 36600 163800 36700
rect 163700 36700 163800 36800
rect 163700 36800 163800 36900
rect 163700 36900 163800 37000
rect 163700 37000 163800 37100
rect 163700 37100 163800 37200
rect 163700 37200 163800 37300
rect 163700 37300 163800 37400
rect 163700 37400 163800 37500
rect 163700 37500 163800 37600
rect 163700 37600 163800 37700
rect 163700 37700 163800 37800
rect 163700 37800 163800 37900
rect 163700 37900 163800 38000
rect 163700 38000 163800 38100
rect 163700 38100 163800 38200
rect 163700 38200 163800 38300
rect 163800 33100 163900 33200
rect 163800 33200 163900 33300
rect 163800 33300 163900 33400
rect 163800 33400 163900 33500
rect 163800 33500 163900 33600
rect 163800 33600 163900 33700
rect 163800 33700 163900 33800
rect 163800 33800 163900 33900
rect 163800 33900 163900 34000
rect 163800 34000 163900 34100
rect 163800 34100 163900 34200
rect 163800 34200 163900 34300
rect 163800 34300 163900 34400
rect 163800 34400 163900 34500
rect 163800 34500 163900 34600
rect 163800 34600 163900 34700
rect 163800 34700 163900 34800
rect 163800 34800 163900 34900
rect 163800 34900 163900 35000
rect 163800 35000 163900 35100
rect 163800 35100 163900 35200
rect 163800 35200 163900 35300
rect 163800 35300 163900 35400
rect 163800 35400 163900 35500
rect 163800 35500 163900 35600
rect 163800 35600 163900 35700
rect 163800 35700 163900 35800
rect 163800 35800 163900 35900
rect 163800 35900 163900 36000
rect 163800 36000 163900 36100
rect 163800 36100 163900 36200
rect 163800 36200 163900 36300
rect 163800 36300 163900 36400
rect 163800 36400 163900 36500
rect 163800 36500 163900 36600
rect 163800 36600 163900 36700
rect 163800 36700 163900 36800
rect 163800 36800 163900 36900
rect 163800 36900 163900 37000
rect 163800 37000 163900 37100
rect 163800 37100 163900 37200
rect 163800 37200 163900 37300
rect 163800 37300 163900 37400
rect 163800 37400 163900 37500
rect 163800 37500 163900 37600
rect 163800 37600 163900 37700
rect 163800 37700 163900 37800
rect 163800 37800 163900 37900
rect 163800 37900 163900 38000
rect 163800 38000 163900 38100
rect 163800 38100 163900 38200
rect 163800 38200 163900 38300
rect 163900 32800 164000 32900
rect 163900 32900 164000 33000
rect 163900 33000 164000 33100
rect 163900 33100 164000 33200
rect 163900 33200 164000 33300
rect 163900 33300 164000 33400
rect 163900 33400 164000 33500
rect 163900 33500 164000 33600
rect 163900 33600 164000 33700
rect 163900 33700 164000 33800
rect 163900 33800 164000 33900
rect 163900 33900 164000 34000
rect 163900 34000 164000 34100
rect 163900 34100 164000 34200
rect 163900 34200 164000 34300
rect 163900 34300 164000 34400
rect 163900 34400 164000 34500
rect 163900 34500 164000 34600
rect 163900 34600 164000 34700
rect 163900 34700 164000 34800
rect 163900 34800 164000 34900
rect 163900 34900 164000 35000
rect 163900 35000 164000 35100
rect 163900 35100 164000 35200
rect 163900 35200 164000 35300
rect 163900 35300 164000 35400
rect 163900 35400 164000 35500
rect 163900 35500 164000 35600
rect 163900 35600 164000 35700
rect 163900 35700 164000 35800
rect 163900 35800 164000 35900
rect 163900 35900 164000 36000
rect 163900 36000 164000 36100
rect 163900 36100 164000 36200
rect 163900 36200 164000 36300
rect 163900 36300 164000 36400
rect 163900 36400 164000 36500
rect 163900 36500 164000 36600
rect 163900 36600 164000 36700
rect 163900 36700 164000 36800
rect 163900 36800 164000 36900
rect 163900 36900 164000 37000
rect 163900 37000 164000 37100
rect 163900 37100 164000 37200
rect 163900 37200 164000 37300
rect 163900 37300 164000 37400
rect 163900 37400 164000 37500
rect 163900 37500 164000 37600
rect 163900 37600 164000 37700
rect 163900 37700 164000 37800
rect 163900 37800 164000 37900
rect 163900 37900 164000 38000
rect 163900 38000 164000 38100
rect 163900 38100 164000 38200
rect 163900 38200 164000 38300
rect 164000 32500 164100 32600
rect 164000 32600 164100 32700
rect 164000 32700 164100 32800
rect 164000 32800 164100 32900
rect 164000 32900 164100 33000
rect 164000 33000 164100 33100
rect 164000 33100 164100 33200
rect 164000 33200 164100 33300
rect 164000 33300 164100 33400
rect 164000 33400 164100 33500
rect 164000 33500 164100 33600
rect 164000 33600 164100 33700
rect 164000 33700 164100 33800
rect 164000 33800 164100 33900
rect 164000 33900 164100 34000
rect 164000 34000 164100 34100
rect 164000 34100 164100 34200
rect 164000 34200 164100 34300
rect 164000 34300 164100 34400
rect 164000 34400 164100 34500
rect 164000 34500 164100 34600
rect 164000 34600 164100 34700
rect 164000 34700 164100 34800
rect 164000 34800 164100 34900
rect 164000 34900 164100 35000
rect 164000 35000 164100 35100
rect 164000 35100 164100 35200
rect 164000 35200 164100 35300
rect 164000 35300 164100 35400
rect 164000 35400 164100 35500
rect 164000 35500 164100 35600
rect 164000 35600 164100 35700
rect 164000 35700 164100 35800
rect 164000 35800 164100 35900
rect 164000 35900 164100 36000
rect 164000 36000 164100 36100
rect 164000 36100 164100 36200
rect 164000 36200 164100 36300
rect 164000 36300 164100 36400
rect 164000 36400 164100 36500
rect 164000 36500 164100 36600
rect 164000 36600 164100 36700
rect 164000 36700 164100 36800
rect 164000 36800 164100 36900
rect 164000 36900 164100 37000
rect 164000 37000 164100 37100
rect 164000 37100 164100 37200
rect 164000 37200 164100 37300
rect 164000 37300 164100 37400
rect 164000 37400 164100 37500
rect 164000 37500 164100 37600
rect 164000 37600 164100 37700
rect 164000 37700 164100 37800
rect 164000 37800 164100 37900
rect 164000 37900 164100 38000
rect 164000 38000 164100 38100
rect 164000 38100 164100 38200
rect 164100 32200 164200 32300
rect 164100 32300 164200 32400
rect 164100 32400 164200 32500
rect 164100 32500 164200 32600
rect 164100 32600 164200 32700
rect 164100 32700 164200 32800
rect 164100 32800 164200 32900
rect 164100 32900 164200 33000
rect 164100 33000 164200 33100
rect 164100 33100 164200 33200
rect 164100 33200 164200 33300
rect 164100 33300 164200 33400
rect 164100 33400 164200 33500
rect 164100 33500 164200 33600
rect 164100 33600 164200 33700
rect 164100 33700 164200 33800
rect 164100 33800 164200 33900
rect 164100 33900 164200 34000
rect 164100 34000 164200 34100
rect 164100 34100 164200 34200
rect 164100 34200 164200 34300
rect 164100 34300 164200 34400
rect 164100 34400 164200 34500
rect 164100 34500 164200 34600
rect 164100 34600 164200 34700
rect 164100 34700 164200 34800
rect 164100 34800 164200 34900
rect 164100 34900 164200 35000
rect 164100 35000 164200 35100
rect 164100 35100 164200 35200
rect 164100 35200 164200 35300
rect 164100 35300 164200 35400
rect 164100 35400 164200 35500
rect 164100 35500 164200 35600
rect 164100 35600 164200 35700
rect 164100 35700 164200 35800
rect 164100 35800 164200 35900
rect 164100 35900 164200 36000
rect 164100 36000 164200 36100
rect 164100 36100 164200 36200
rect 164100 36200 164200 36300
rect 164100 36300 164200 36400
rect 164100 36400 164200 36500
rect 164100 36500 164200 36600
rect 164100 36600 164200 36700
rect 164100 36700 164200 36800
rect 164100 36800 164200 36900
rect 164100 36900 164200 37000
rect 164100 37000 164200 37100
rect 164100 37100 164200 37200
rect 164100 37200 164200 37300
rect 164100 37300 164200 37400
rect 164100 37400 164200 37500
rect 164100 37500 164200 37600
rect 164100 37600 164200 37700
rect 164100 37700 164200 37800
rect 164100 37800 164200 37900
rect 164100 37900 164200 38000
rect 164100 38000 164200 38100
rect 164100 38100 164200 38200
rect 164200 31900 164300 32000
rect 164200 32000 164300 32100
rect 164200 32100 164300 32200
rect 164200 32200 164300 32300
rect 164200 32300 164300 32400
rect 164200 32400 164300 32500
rect 164200 32500 164300 32600
rect 164200 32600 164300 32700
rect 164200 32700 164300 32800
rect 164200 32800 164300 32900
rect 164200 32900 164300 33000
rect 164200 33000 164300 33100
rect 164200 33100 164300 33200
rect 164200 33200 164300 33300
rect 164200 33300 164300 33400
rect 164200 33400 164300 33500
rect 164200 33500 164300 33600
rect 164200 33600 164300 33700
rect 164200 33700 164300 33800
rect 164200 33800 164300 33900
rect 164200 33900 164300 34000
rect 164200 34000 164300 34100
rect 164200 34100 164300 34200
rect 164200 34200 164300 34300
rect 164200 34300 164300 34400
rect 164200 34400 164300 34500
rect 164200 34500 164300 34600
rect 164200 34600 164300 34700
rect 164200 34700 164300 34800
rect 164200 34800 164300 34900
rect 164200 34900 164300 35000
rect 164200 35000 164300 35100
rect 164200 35100 164300 35200
rect 164200 35200 164300 35300
rect 164200 35300 164300 35400
rect 164200 35400 164300 35500
rect 164200 35500 164300 35600
rect 164200 35600 164300 35700
rect 164200 35700 164300 35800
rect 164200 35800 164300 35900
rect 164200 35900 164300 36000
rect 164200 36000 164300 36100
rect 164200 36100 164300 36200
rect 164200 36200 164300 36300
rect 164200 36300 164300 36400
rect 164200 36400 164300 36500
rect 164200 36500 164300 36600
rect 164200 36600 164300 36700
rect 164200 36700 164300 36800
rect 164200 36800 164300 36900
rect 164200 36900 164300 37000
rect 164200 37000 164300 37100
rect 164200 37100 164300 37200
rect 164200 37200 164300 37300
rect 164200 37300 164300 37400
rect 164200 37400 164300 37500
rect 164200 37500 164300 37600
rect 164200 37600 164300 37700
rect 164200 37700 164300 37800
rect 164200 37800 164300 37900
rect 164200 37900 164300 38000
rect 164200 38000 164300 38100
rect 164300 31500 164400 31600
rect 164300 31600 164400 31700
rect 164300 31700 164400 31800
rect 164300 31800 164400 31900
rect 164300 31900 164400 32000
rect 164300 32000 164400 32100
rect 164300 32100 164400 32200
rect 164300 32200 164400 32300
rect 164300 32300 164400 32400
rect 164300 32400 164400 32500
rect 164300 32500 164400 32600
rect 164300 32600 164400 32700
rect 164300 32700 164400 32800
rect 164300 32800 164400 32900
rect 164300 32900 164400 33000
rect 164300 33000 164400 33100
rect 164300 33100 164400 33200
rect 164300 33200 164400 33300
rect 164300 33300 164400 33400
rect 164300 33400 164400 33500
rect 164300 33500 164400 33600
rect 164300 33600 164400 33700
rect 164300 33700 164400 33800
rect 164300 33800 164400 33900
rect 164300 33900 164400 34000
rect 164300 34000 164400 34100
rect 164300 34100 164400 34200
rect 164300 34200 164400 34300
rect 164300 34300 164400 34400
rect 164300 34400 164400 34500
rect 164300 34500 164400 34600
rect 164300 34600 164400 34700
rect 164300 34700 164400 34800
rect 164300 34800 164400 34900
rect 164300 34900 164400 35000
rect 164300 35000 164400 35100
rect 164300 35100 164400 35200
rect 164300 35200 164400 35300
rect 164300 35300 164400 35400
rect 164300 35400 164400 35500
rect 164300 35500 164400 35600
rect 164300 35600 164400 35700
rect 164300 35700 164400 35800
rect 164300 35800 164400 35900
rect 164300 35900 164400 36000
rect 164300 36000 164400 36100
rect 164300 36100 164400 36200
rect 164300 36200 164400 36300
rect 164300 36300 164400 36400
rect 164300 36400 164400 36500
rect 164300 36500 164400 36600
rect 164300 36600 164400 36700
rect 164300 36700 164400 36800
rect 164300 36800 164400 36900
rect 164300 36900 164400 37000
rect 164300 37000 164400 37100
rect 164300 37100 164400 37200
rect 164300 37200 164400 37300
rect 164300 37300 164400 37400
rect 164300 37400 164400 37500
rect 164300 37500 164400 37600
rect 164300 37600 164400 37700
rect 164300 37700 164400 37800
rect 164300 37800 164400 37900
rect 164300 37900 164400 38000
rect 164400 31200 164500 31300
rect 164400 31300 164500 31400
rect 164400 31400 164500 31500
rect 164400 31500 164500 31600
rect 164400 31600 164500 31700
rect 164400 31700 164500 31800
rect 164400 31800 164500 31900
rect 164400 31900 164500 32000
rect 164400 32000 164500 32100
rect 164400 32100 164500 32200
rect 164400 32200 164500 32300
rect 164400 32300 164500 32400
rect 164400 32400 164500 32500
rect 164400 32500 164500 32600
rect 164400 32600 164500 32700
rect 164400 32700 164500 32800
rect 164400 32800 164500 32900
rect 164400 32900 164500 33000
rect 164400 33000 164500 33100
rect 164400 33100 164500 33200
rect 164400 33200 164500 33300
rect 164400 33300 164500 33400
rect 164400 33400 164500 33500
rect 164400 33500 164500 33600
rect 164400 33600 164500 33700
rect 164400 33700 164500 33800
rect 164400 33800 164500 33900
rect 164400 33900 164500 34000
rect 164400 34000 164500 34100
rect 164400 34100 164500 34200
rect 164400 34200 164500 34300
rect 164400 34300 164500 34400
rect 164400 34400 164500 34500
rect 164400 34500 164500 34600
rect 164400 34600 164500 34700
rect 164400 34700 164500 34800
rect 164400 34800 164500 34900
rect 164400 34900 164500 35000
rect 164400 35000 164500 35100
rect 164400 35100 164500 35200
rect 164400 35200 164500 35300
rect 164400 35300 164500 35400
rect 164400 35400 164500 35500
rect 164400 35500 164500 35600
rect 164400 35600 164500 35700
rect 164400 35700 164500 35800
rect 164400 35800 164500 35900
rect 164400 35900 164500 36000
rect 164400 36000 164500 36100
rect 164400 36100 164500 36200
rect 164400 36200 164500 36300
rect 164400 36300 164500 36400
rect 164400 36400 164500 36500
rect 164400 36500 164500 36600
rect 164400 36600 164500 36700
rect 164400 36700 164500 36800
rect 164400 36800 164500 36900
rect 164400 36900 164500 37000
rect 164400 37000 164500 37100
rect 164400 37100 164500 37200
rect 164400 37200 164500 37300
rect 164400 37300 164500 37400
rect 164400 37400 164500 37500
rect 164400 37500 164500 37600
rect 164400 37600 164500 37700
rect 164400 37700 164500 37800
rect 164400 37800 164500 37900
rect 164500 30900 164600 31000
rect 164500 31000 164600 31100
rect 164500 31100 164600 31200
rect 164500 31200 164600 31300
rect 164500 31300 164600 31400
rect 164500 31400 164600 31500
rect 164500 31500 164600 31600
rect 164500 31600 164600 31700
rect 164500 31700 164600 31800
rect 164500 31800 164600 31900
rect 164500 31900 164600 32000
rect 164500 32000 164600 32100
rect 164500 32100 164600 32200
rect 164500 32200 164600 32300
rect 164500 32300 164600 32400
rect 164500 32400 164600 32500
rect 164500 32500 164600 32600
rect 164500 32600 164600 32700
rect 164500 32700 164600 32800
rect 164500 32800 164600 32900
rect 164500 32900 164600 33000
rect 164500 33000 164600 33100
rect 164500 33100 164600 33200
rect 164500 33200 164600 33300
rect 164500 33300 164600 33400
rect 164500 33400 164600 33500
rect 164500 33500 164600 33600
rect 164500 33600 164600 33700
rect 164500 33700 164600 33800
rect 164500 33800 164600 33900
rect 164500 33900 164600 34000
rect 164500 34000 164600 34100
rect 164500 34100 164600 34200
rect 164500 34200 164600 34300
rect 164500 34300 164600 34400
rect 164500 34400 164600 34500
rect 164500 34500 164600 34600
rect 164500 34600 164600 34700
rect 164500 34700 164600 34800
rect 164500 34800 164600 34900
rect 164500 34900 164600 35000
rect 164500 35000 164600 35100
rect 164500 35100 164600 35200
rect 164500 35200 164600 35300
rect 164500 35300 164600 35400
rect 164500 35400 164600 35500
rect 164500 35500 164600 35600
rect 164500 35600 164600 35700
rect 164500 35700 164600 35800
rect 164500 35800 164600 35900
rect 164500 35900 164600 36000
rect 164500 36000 164600 36100
rect 164500 36100 164600 36200
rect 164500 36200 164600 36300
rect 164500 36300 164600 36400
rect 164500 36400 164600 36500
rect 164500 36500 164600 36600
rect 164500 36600 164600 36700
rect 164500 36700 164600 36800
rect 164500 36800 164600 36900
rect 164500 36900 164600 37000
rect 164500 37000 164600 37100
rect 164500 37100 164600 37200
rect 164500 37200 164600 37300
rect 164500 37300 164600 37400
rect 164500 37400 164600 37500
rect 164500 37500 164600 37600
rect 164500 37600 164600 37700
rect 164500 37700 164600 37800
rect 164600 30500 164700 30600
rect 164600 30600 164700 30700
rect 164600 30700 164700 30800
rect 164600 30800 164700 30900
rect 164600 30900 164700 31000
rect 164600 31000 164700 31100
rect 164600 31100 164700 31200
rect 164600 31200 164700 31300
rect 164600 31300 164700 31400
rect 164600 31400 164700 31500
rect 164600 31500 164700 31600
rect 164600 31600 164700 31700
rect 164600 31700 164700 31800
rect 164600 31800 164700 31900
rect 164600 31900 164700 32000
rect 164600 32000 164700 32100
rect 164600 32100 164700 32200
rect 164600 32200 164700 32300
rect 164600 32300 164700 32400
rect 164600 32400 164700 32500
rect 164600 32500 164700 32600
rect 164600 32600 164700 32700
rect 164600 32700 164700 32800
rect 164600 32800 164700 32900
rect 164600 32900 164700 33000
rect 164600 33000 164700 33100
rect 164600 33100 164700 33200
rect 164600 33200 164700 33300
rect 164600 33300 164700 33400
rect 164600 33400 164700 33500
rect 164600 33500 164700 33600
rect 164600 33600 164700 33700
rect 164600 33700 164700 33800
rect 164600 33800 164700 33900
rect 164600 33900 164700 34000
rect 164600 34000 164700 34100
rect 164600 34100 164700 34200
rect 164600 34200 164700 34300
rect 164600 34300 164700 34400
rect 164600 34400 164700 34500
rect 164600 34500 164700 34600
rect 164600 34600 164700 34700
rect 164600 34700 164700 34800
rect 164600 34800 164700 34900
rect 164600 34900 164700 35000
rect 164600 35000 164700 35100
rect 164600 35100 164700 35200
rect 164600 35200 164700 35300
rect 164600 35300 164700 35400
rect 164600 35400 164700 35500
rect 164600 35500 164700 35600
rect 164600 35600 164700 35700
rect 164600 35700 164700 35800
rect 164600 35800 164700 35900
rect 164600 35900 164700 36000
rect 164600 36000 164700 36100
rect 164600 36100 164700 36200
rect 164600 36200 164700 36300
rect 164600 36300 164700 36400
rect 164600 36400 164700 36500
rect 164600 36500 164700 36600
rect 164600 36600 164700 36700
rect 164600 36700 164700 36800
rect 164600 36800 164700 36900
rect 164600 36900 164700 37000
rect 164600 37000 164700 37100
rect 164600 37100 164700 37200
rect 164600 37200 164700 37300
rect 164600 37300 164700 37400
rect 164600 37400 164700 37500
rect 164600 37500 164700 37600
rect 164600 37600 164700 37700
rect 164700 30100 164800 30200
rect 164700 30200 164800 30300
rect 164700 30300 164800 30400
rect 164700 30400 164800 30500
rect 164700 30500 164800 30600
rect 164700 30600 164800 30700
rect 164700 30700 164800 30800
rect 164700 30800 164800 30900
rect 164700 30900 164800 31000
rect 164700 31000 164800 31100
rect 164700 31100 164800 31200
rect 164700 31200 164800 31300
rect 164700 31300 164800 31400
rect 164700 31400 164800 31500
rect 164700 31500 164800 31600
rect 164700 31600 164800 31700
rect 164700 31700 164800 31800
rect 164700 31800 164800 31900
rect 164700 31900 164800 32000
rect 164700 32000 164800 32100
rect 164700 32100 164800 32200
rect 164700 32200 164800 32300
rect 164700 32300 164800 32400
rect 164700 32400 164800 32500
rect 164700 32500 164800 32600
rect 164700 32600 164800 32700
rect 164700 32700 164800 32800
rect 164700 32800 164800 32900
rect 164700 32900 164800 33000
rect 164700 33000 164800 33100
rect 164700 33100 164800 33200
rect 164700 33200 164800 33300
rect 164700 33300 164800 33400
rect 164700 33400 164800 33500
rect 164700 33500 164800 33600
rect 164700 33600 164800 33700
rect 164700 33700 164800 33800
rect 164700 33800 164800 33900
rect 164700 33900 164800 34000
rect 164700 34000 164800 34100
rect 164700 34100 164800 34200
rect 164700 34200 164800 34300
rect 164700 34300 164800 34400
rect 164700 34400 164800 34500
rect 164700 34500 164800 34600
rect 164700 34600 164800 34700
rect 164700 34700 164800 34800
rect 164700 34800 164800 34900
rect 164700 34900 164800 35000
rect 164700 35000 164800 35100
rect 164700 35100 164800 35200
rect 164700 35200 164800 35300
rect 164700 35300 164800 35400
rect 164700 35400 164800 35500
rect 164700 35500 164800 35600
rect 164700 35600 164800 35700
rect 164700 35700 164800 35800
rect 164700 35800 164800 35900
rect 164700 35900 164800 36000
rect 164700 36000 164800 36100
rect 164700 36100 164800 36200
rect 164700 36200 164800 36300
rect 164700 36300 164800 36400
rect 164700 36400 164800 36500
rect 164700 36500 164800 36600
rect 164700 36600 164800 36700
rect 164700 36700 164800 36800
rect 164700 36800 164800 36900
rect 164700 36900 164800 37000
rect 164700 37000 164800 37100
rect 164700 37100 164800 37200
rect 164700 37200 164800 37300
rect 164700 37300 164800 37400
rect 164800 29800 164900 29900
rect 164800 29900 164900 30000
rect 164800 30000 164900 30100
rect 164800 30100 164900 30200
rect 164800 30200 164900 30300
rect 164800 30300 164900 30400
rect 164800 30400 164900 30500
rect 164800 30500 164900 30600
rect 164800 30600 164900 30700
rect 164800 30700 164900 30800
rect 164800 30800 164900 30900
rect 164800 30900 164900 31000
rect 164800 31000 164900 31100
rect 164800 31100 164900 31200
rect 164800 31200 164900 31300
rect 164800 31300 164900 31400
rect 164800 31400 164900 31500
rect 164800 31500 164900 31600
rect 164800 31600 164900 31700
rect 164800 31700 164900 31800
rect 164800 31800 164900 31900
rect 164800 31900 164900 32000
rect 164800 32000 164900 32100
rect 164800 32100 164900 32200
rect 164800 32200 164900 32300
rect 164800 32300 164900 32400
rect 164800 32400 164900 32500
rect 164800 32500 164900 32600
rect 164800 32600 164900 32700
rect 164800 32700 164900 32800
rect 164800 32800 164900 32900
rect 164800 32900 164900 33000
rect 164800 33000 164900 33100
rect 164800 33100 164900 33200
rect 164800 33200 164900 33300
rect 164800 33300 164900 33400
rect 164800 33400 164900 33500
rect 164800 33500 164900 33600
rect 164800 33600 164900 33700
rect 164800 33700 164900 33800
rect 164800 33800 164900 33900
rect 164800 33900 164900 34000
rect 164800 34000 164900 34100
rect 164800 34100 164900 34200
rect 164800 34200 164900 34300
rect 164800 34300 164900 34400
rect 164800 34400 164900 34500
rect 164800 34500 164900 34600
rect 164800 34600 164900 34700
rect 164800 34700 164900 34800
rect 164800 34800 164900 34900
rect 164800 34900 164900 35000
rect 164800 35000 164900 35100
rect 164800 35100 164900 35200
rect 164800 35200 164900 35300
rect 164800 35300 164900 35400
rect 164800 35400 164900 35500
rect 164800 35500 164900 35600
rect 164800 35600 164900 35700
rect 164800 35700 164900 35800
rect 164800 35800 164900 35900
rect 164800 35900 164900 36000
rect 164800 36000 164900 36100
rect 164800 36100 164900 36200
rect 164800 36200 164900 36300
rect 164800 36300 164900 36400
rect 164800 36400 164900 36500
rect 164800 36500 164900 36600
rect 164800 36600 164900 36700
rect 164800 36700 164900 36800
rect 164800 36800 164900 36900
rect 164800 36900 164900 37000
rect 164800 37000 164900 37100
rect 164800 37100 164900 37200
rect 164900 29400 165000 29500
rect 164900 29500 165000 29600
rect 164900 29600 165000 29700
rect 164900 29700 165000 29800
rect 164900 29800 165000 29900
rect 164900 29900 165000 30000
rect 164900 30000 165000 30100
rect 164900 30100 165000 30200
rect 164900 30200 165000 30300
rect 164900 30300 165000 30400
rect 164900 30400 165000 30500
rect 164900 30500 165000 30600
rect 164900 30600 165000 30700
rect 164900 30700 165000 30800
rect 164900 30800 165000 30900
rect 164900 30900 165000 31000
rect 164900 31000 165000 31100
rect 164900 31100 165000 31200
rect 164900 31200 165000 31300
rect 164900 31300 165000 31400
rect 164900 31400 165000 31500
rect 164900 31500 165000 31600
rect 164900 31600 165000 31700
rect 164900 31700 165000 31800
rect 164900 31800 165000 31900
rect 164900 31900 165000 32000
rect 164900 32000 165000 32100
rect 164900 32100 165000 32200
rect 164900 32200 165000 32300
rect 164900 32300 165000 32400
rect 164900 32400 165000 32500
rect 164900 32500 165000 32600
rect 164900 32600 165000 32700
rect 164900 32700 165000 32800
rect 164900 32800 165000 32900
rect 164900 32900 165000 33000
rect 164900 33000 165000 33100
rect 164900 33100 165000 33200
rect 164900 33200 165000 33300
rect 164900 33300 165000 33400
rect 164900 33400 165000 33500
rect 164900 33500 165000 33600
rect 164900 33600 165000 33700
rect 164900 33700 165000 33800
rect 164900 33800 165000 33900
rect 164900 33900 165000 34000
rect 164900 34000 165000 34100
rect 164900 34100 165000 34200
rect 164900 34200 165000 34300
rect 164900 34300 165000 34400
rect 164900 34400 165000 34500
rect 164900 34500 165000 34600
rect 164900 34600 165000 34700
rect 164900 34700 165000 34800
rect 164900 34800 165000 34900
rect 164900 34900 165000 35000
rect 164900 35000 165000 35100
rect 164900 35100 165000 35200
rect 164900 35200 165000 35300
rect 164900 35300 165000 35400
rect 164900 35400 165000 35500
rect 164900 35500 165000 35600
rect 164900 35600 165000 35700
rect 164900 35700 165000 35800
rect 164900 35800 165000 35900
rect 164900 35900 165000 36000
rect 164900 36000 165000 36100
rect 164900 36100 165000 36200
rect 164900 36200 165000 36300
rect 164900 36300 165000 36400
rect 164900 36400 165000 36500
rect 164900 36500 165000 36600
rect 164900 36600 165000 36700
rect 164900 36700 165000 36800
rect 164900 36800 165000 36900
rect 165000 29000 165100 29100
rect 165000 29100 165100 29200
rect 165000 29200 165100 29300
rect 165000 29300 165100 29400
rect 165000 29400 165100 29500
rect 165000 29500 165100 29600
rect 165000 29600 165100 29700
rect 165000 29700 165100 29800
rect 165000 29800 165100 29900
rect 165000 29900 165100 30000
rect 165000 30000 165100 30100
rect 165000 30100 165100 30200
rect 165000 30200 165100 30300
rect 165000 30300 165100 30400
rect 165000 30400 165100 30500
rect 165000 30500 165100 30600
rect 165000 30600 165100 30700
rect 165000 30700 165100 30800
rect 165000 30800 165100 30900
rect 165000 30900 165100 31000
rect 165000 31000 165100 31100
rect 165000 31100 165100 31200
rect 165000 31200 165100 31300
rect 165000 31300 165100 31400
rect 165000 31400 165100 31500
rect 165000 31500 165100 31600
rect 165000 31600 165100 31700
rect 165000 31700 165100 31800
rect 165000 31800 165100 31900
rect 165000 31900 165100 32000
rect 165000 32000 165100 32100
rect 165000 32100 165100 32200
rect 165000 32200 165100 32300
rect 165000 32300 165100 32400
rect 165000 32400 165100 32500
rect 165000 32500 165100 32600
rect 165000 32600 165100 32700
rect 165000 32700 165100 32800
rect 165000 32800 165100 32900
rect 165000 32900 165100 33000
rect 165000 33000 165100 33100
rect 165000 33100 165100 33200
rect 165000 33200 165100 33300
rect 165000 33300 165100 33400
rect 165000 33400 165100 33500
rect 165000 33500 165100 33600
rect 165000 33600 165100 33700
rect 165000 33700 165100 33800
rect 165000 33800 165100 33900
rect 165000 33900 165100 34000
rect 165000 34000 165100 34100
rect 165000 34100 165100 34200
rect 165000 34200 165100 34300
rect 165000 34300 165100 34400
rect 165000 34400 165100 34500
rect 165000 34500 165100 34600
rect 165000 34600 165100 34700
rect 165000 34700 165100 34800
rect 165000 34800 165100 34900
rect 165000 34900 165100 35000
rect 165000 35000 165100 35100
rect 165000 35100 165100 35200
rect 165000 35200 165100 35300
rect 165000 35300 165100 35400
rect 165000 35400 165100 35500
rect 165000 35500 165100 35600
rect 165000 35600 165100 35700
rect 165000 35700 165100 35800
rect 165000 35800 165100 35900
rect 165000 35900 165100 36000
rect 165000 36000 165100 36100
rect 165000 36100 165100 36200
rect 165000 36200 165100 36300
rect 165000 36300 165100 36400
rect 165000 36400 165100 36500
rect 165000 36500 165100 36600
rect 165100 28500 165200 28600
rect 165100 28600 165200 28700
rect 165100 28700 165200 28800
rect 165100 28800 165200 28900
rect 165100 28900 165200 29000
rect 165100 29000 165200 29100
rect 165100 29100 165200 29200
rect 165100 29200 165200 29300
rect 165100 29300 165200 29400
rect 165100 29400 165200 29500
rect 165100 29500 165200 29600
rect 165100 29600 165200 29700
rect 165100 29700 165200 29800
rect 165100 29800 165200 29900
rect 165100 29900 165200 30000
rect 165100 30000 165200 30100
rect 165100 30100 165200 30200
rect 165100 30200 165200 30300
rect 165100 30300 165200 30400
rect 165100 30400 165200 30500
rect 165100 30500 165200 30600
rect 165100 30600 165200 30700
rect 165100 30700 165200 30800
rect 165100 30800 165200 30900
rect 165100 30900 165200 31000
rect 165100 31000 165200 31100
rect 165100 31100 165200 31200
rect 165100 31200 165200 31300
rect 165100 31300 165200 31400
rect 165100 31400 165200 31500
rect 165100 31500 165200 31600
rect 165100 31600 165200 31700
rect 165100 31700 165200 31800
rect 165100 31800 165200 31900
rect 165100 31900 165200 32000
rect 165100 32000 165200 32100
rect 165100 32100 165200 32200
rect 165100 32200 165200 32300
rect 165100 32300 165200 32400
rect 165100 32400 165200 32500
rect 165100 32500 165200 32600
rect 165100 32600 165200 32700
rect 165100 32700 165200 32800
rect 165100 32800 165200 32900
rect 165100 32900 165200 33000
rect 165100 33000 165200 33100
rect 165100 33100 165200 33200
rect 165100 33200 165200 33300
rect 165100 33300 165200 33400
rect 165100 33400 165200 33500
rect 165100 33500 165200 33600
rect 165100 33600 165200 33700
rect 165100 33700 165200 33800
rect 165100 33800 165200 33900
rect 165100 33900 165200 34000
rect 165100 34000 165200 34100
rect 165100 34100 165200 34200
rect 165100 34200 165200 34300
rect 165100 34300 165200 34400
rect 165100 34400 165200 34500
rect 165100 34500 165200 34600
rect 165100 34600 165200 34700
rect 165100 34700 165200 34800
rect 165100 34800 165200 34900
rect 165100 34900 165200 35000
rect 165100 35000 165200 35100
rect 165100 35100 165200 35200
rect 165100 35200 165200 35300
rect 165100 35300 165200 35400
rect 165100 35400 165200 35500
rect 165100 35500 165200 35600
rect 165100 35600 165200 35700
rect 165100 35700 165200 35800
rect 165100 35800 165200 35900
rect 165100 35900 165200 36000
rect 165100 36000 165200 36100
rect 165100 36100 165200 36200
rect 165100 36200 165200 36300
rect 165200 28100 165300 28200
rect 165200 28200 165300 28300
rect 165200 28300 165300 28400
rect 165200 28400 165300 28500
rect 165200 28500 165300 28600
rect 165200 28600 165300 28700
rect 165200 28700 165300 28800
rect 165200 28800 165300 28900
rect 165200 28900 165300 29000
rect 165200 29000 165300 29100
rect 165200 29100 165300 29200
rect 165200 29200 165300 29300
rect 165200 29300 165300 29400
rect 165200 29400 165300 29500
rect 165200 29500 165300 29600
rect 165200 29600 165300 29700
rect 165200 29700 165300 29800
rect 165200 29800 165300 29900
rect 165200 29900 165300 30000
rect 165200 30000 165300 30100
rect 165200 30100 165300 30200
rect 165200 30200 165300 30300
rect 165200 30300 165300 30400
rect 165200 30400 165300 30500
rect 165200 30500 165300 30600
rect 165200 30600 165300 30700
rect 165200 30700 165300 30800
rect 165200 30800 165300 30900
rect 165200 30900 165300 31000
rect 165200 31000 165300 31100
rect 165200 31100 165300 31200
rect 165200 31200 165300 31300
rect 165200 31300 165300 31400
rect 165200 31400 165300 31500
rect 165200 31500 165300 31600
rect 165200 31600 165300 31700
rect 165200 31700 165300 31800
rect 165200 31800 165300 31900
rect 165200 31900 165300 32000
rect 165200 32000 165300 32100
rect 165200 32100 165300 32200
rect 165200 32200 165300 32300
rect 165200 32300 165300 32400
rect 165200 32400 165300 32500
rect 165200 32500 165300 32600
rect 165200 32600 165300 32700
rect 165200 32700 165300 32800
rect 165200 32800 165300 32900
rect 165200 32900 165300 33000
rect 165200 33000 165300 33100
rect 165200 33100 165300 33200
rect 165200 33200 165300 33300
rect 165200 33300 165300 33400
rect 165200 33400 165300 33500
rect 165200 33500 165300 33600
rect 165200 33600 165300 33700
rect 165200 33700 165300 33800
rect 165200 33800 165300 33900
rect 165200 33900 165300 34000
rect 165200 34000 165300 34100
rect 165200 34100 165300 34200
rect 165200 34200 165300 34300
rect 165200 34300 165300 34400
rect 165200 34400 165300 34500
rect 165200 34500 165300 34600
rect 165200 34600 165300 34700
rect 165200 34700 165300 34800
rect 165200 34800 165300 34900
rect 165200 34900 165300 35000
rect 165200 35000 165300 35100
rect 165200 35100 165300 35200
rect 165200 35200 165300 35300
rect 165200 35300 165300 35400
rect 165200 35400 165300 35500
rect 165200 35500 165300 35600
rect 165200 35600 165300 35700
rect 165200 35700 165300 35800
rect 165200 35800 165300 35900
rect 165200 35900 165300 36000
rect 165300 27600 165400 27700
rect 165300 27700 165400 27800
rect 165300 27800 165400 27900
rect 165300 27900 165400 28000
rect 165300 28000 165400 28100
rect 165300 28100 165400 28200
rect 165300 28200 165400 28300
rect 165300 28300 165400 28400
rect 165300 28400 165400 28500
rect 165300 28500 165400 28600
rect 165300 28600 165400 28700
rect 165300 28700 165400 28800
rect 165300 28800 165400 28900
rect 165300 28900 165400 29000
rect 165300 29000 165400 29100
rect 165300 29100 165400 29200
rect 165300 29200 165400 29300
rect 165300 29300 165400 29400
rect 165300 29400 165400 29500
rect 165300 29500 165400 29600
rect 165300 29600 165400 29700
rect 165300 29700 165400 29800
rect 165300 29800 165400 29900
rect 165300 29900 165400 30000
rect 165300 30000 165400 30100
rect 165300 30100 165400 30200
rect 165300 30200 165400 30300
rect 165300 30300 165400 30400
rect 165300 30400 165400 30500
rect 165300 30500 165400 30600
rect 165300 30600 165400 30700
rect 165300 30700 165400 30800
rect 165300 30800 165400 30900
rect 165300 30900 165400 31000
rect 165300 31000 165400 31100
rect 165300 31100 165400 31200
rect 165300 31200 165400 31300
rect 165300 31300 165400 31400
rect 165300 31400 165400 31500
rect 165300 31500 165400 31600
rect 165300 31600 165400 31700
rect 165300 31700 165400 31800
rect 165300 31800 165400 31900
rect 165300 31900 165400 32000
rect 165300 32000 165400 32100
rect 165300 32100 165400 32200
rect 165300 32200 165400 32300
rect 165300 32300 165400 32400
rect 165300 32400 165400 32500
rect 165300 32500 165400 32600
rect 165300 32600 165400 32700
rect 165300 32700 165400 32800
rect 165300 32800 165400 32900
rect 165300 32900 165400 33000
rect 165300 33000 165400 33100
rect 165300 33100 165400 33200
rect 165300 33200 165400 33300
rect 165300 33300 165400 33400
rect 165300 33400 165400 33500
rect 165300 33500 165400 33600
rect 165300 33600 165400 33700
rect 165300 33700 165400 33800
rect 165300 33800 165400 33900
rect 165300 33900 165400 34000
rect 165300 34000 165400 34100
rect 165300 34100 165400 34200
rect 165300 34200 165400 34300
rect 165300 34300 165400 34400
rect 165300 34400 165400 34500
rect 165300 34500 165400 34600
rect 165300 34600 165400 34700
rect 165300 34700 165400 34800
rect 165300 34800 165400 34900
rect 165300 34900 165400 35000
rect 165300 35000 165400 35100
rect 165300 35100 165400 35200
rect 165300 35200 165400 35300
rect 165300 35300 165400 35400
rect 165300 35400 165400 35500
rect 165300 35500 165400 35600
rect 165300 35600 165400 35700
rect 165400 27200 165500 27300
rect 165400 27300 165500 27400
rect 165400 27400 165500 27500
rect 165400 27500 165500 27600
rect 165400 27600 165500 27700
rect 165400 27700 165500 27800
rect 165400 27800 165500 27900
rect 165400 27900 165500 28000
rect 165400 28000 165500 28100
rect 165400 28100 165500 28200
rect 165400 28200 165500 28300
rect 165400 28300 165500 28400
rect 165400 28400 165500 28500
rect 165400 28500 165500 28600
rect 165400 28600 165500 28700
rect 165400 28700 165500 28800
rect 165400 28800 165500 28900
rect 165400 28900 165500 29000
rect 165400 29000 165500 29100
rect 165400 29100 165500 29200
rect 165400 29200 165500 29300
rect 165400 29300 165500 29400
rect 165400 29400 165500 29500
rect 165400 29500 165500 29600
rect 165400 29600 165500 29700
rect 165400 29700 165500 29800
rect 165400 29800 165500 29900
rect 165400 29900 165500 30000
rect 165400 30000 165500 30100
rect 165400 30100 165500 30200
rect 165400 30200 165500 30300
rect 165400 30300 165500 30400
rect 165400 30400 165500 30500
rect 165400 30500 165500 30600
rect 165400 30600 165500 30700
rect 165400 30700 165500 30800
rect 165400 30800 165500 30900
rect 165400 30900 165500 31000
rect 165400 31000 165500 31100
rect 165400 31100 165500 31200
rect 165400 31200 165500 31300
rect 165400 31300 165500 31400
rect 165400 31400 165500 31500
rect 165400 31500 165500 31600
rect 165400 31600 165500 31700
rect 165400 31700 165500 31800
rect 165400 31800 165500 31900
rect 165400 31900 165500 32000
rect 165400 32000 165500 32100
rect 165400 32100 165500 32200
rect 165400 32200 165500 32300
rect 165400 32300 165500 32400
rect 165400 32400 165500 32500
rect 165400 32500 165500 32600
rect 165400 32600 165500 32700
rect 165400 32700 165500 32800
rect 165400 32800 165500 32900
rect 165400 32900 165500 33000
rect 165400 33000 165500 33100
rect 165400 33100 165500 33200
rect 165400 33200 165500 33300
rect 165400 33300 165500 33400
rect 165400 33400 165500 33500
rect 165400 33500 165500 33600
rect 165400 33600 165500 33700
rect 165400 33700 165500 33800
rect 165400 33800 165500 33900
rect 165400 33900 165500 34000
rect 165400 34000 165500 34100
rect 165400 34100 165500 34200
rect 165400 34200 165500 34300
rect 165400 34300 165500 34400
rect 165400 34400 165500 34500
rect 165400 34500 165500 34600
rect 165400 34600 165500 34700
rect 165400 34700 165500 34800
rect 165400 34800 165500 34900
rect 165400 34900 165500 35000
rect 165400 35000 165500 35100
rect 165400 35100 165500 35200
rect 165400 35200 165500 35300
rect 165400 35300 165500 35400
rect 165500 26700 165600 26800
rect 165500 26800 165600 26900
rect 165500 26900 165600 27000
rect 165500 27000 165600 27100
rect 165500 27100 165600 27200
rect 165500 27200 165600 27300
rect 165500 27300 165600 27400
rect 165500 27400 165600 27500
rect 165500 27500 165600 27600
rect 165500 27600 165600 27700
rect 165500 27700 165600 27800
rect 165500 27800 165600 27900
rect 165500 27900 165600 28000
rect 165500 28000 165600 28100
rect 165500 28100 165600 28200
rect 165500 28200 165600 28300
rect 165500 28300 165600 28400
rect 165500 28400 165600 28500
rect 165500 28500 165600 28600
rect 165500 28600 165600 28700
rect 165500 28700 165600 28800
rect 165500 28800 165600 28900
rect 165500 28900 165600 29000
rect 165500 29000 165600 29100
rect 165500 29100 165600 29200
rect 165500 29200 165600 29300
rect 165500 29300 165600 29400
rect 165500 29400 165600 29500
rect 165500 29500 165600 29600
rect 165500 29600 165600 29700
rect 165500 29700 165600 29800
rect 165500 29800 165600 29900
rect 165500 29900 165600 30000
rect 165500 30000 165600 30100
rect 165500 30100 165600 30200
rect 165500 30200 165600 30300
rect 165500 30300 165600 30400
rect 165500 30400 165600 30500
rect 165500 30500 165600 30600
rect 165500 30600 165600 30700
rect 165500 30700 165600 30800
rect 165500 30800 165600 30900
rect 165500 30900 165600 31000
rect 165500 31000 165600 31100
rect 165500 31100 165600 31200
rect 165500 31200 165600 31300
rect 165500 31300 165600 31400
rect 165500 31400 165600 31500
rect 165500 31500 165600 31600
rect 165500 31600 165600 31700
rect 165500 31700 165600 31800
rect 165500 31800 165600 31900
rect 165500 31900 165600 32000
rect 165500 32000 165600 32100
rect 165500 32100 165600 32200
rect 165500 32200 165600 32300
rect 165500 32300 165600 32400
rect 165500 32400 165600 32500
rect 165500 32500 165600 32600
rect 165500 32600 165600 32700
rect 165500 32700 165600 32800
rect 165500 32800 165600 32900
rect 165500 32900 165600 33000
rect 165500 33000 165600 33100
rect 165500 33100 165600 33200
rect 165500 33200 165600 33300
rect 165500 33300 165600 33400
rect 165500 33400 165600 33500
rect 165500 33500 165600 33600
rect 165500 33600 165600 33700
rect 165500 33700 165600 33800
rect 165500 33800 165600 33900
rect 165500 33900 165600 34000
rect 165500 34000 165600 34100
rect 165500 34100 165600 34200
rect 165500 34200 165600 34300
rect 165500 34300 165600 34400
rect 165500 34400 165600 34500
rect 165500 34500 165600 34600
rect 165500 34600 165600 34700
rect 165500 34700 165600 34800
rect 165500 34800 165600 34900
rect 165500 34900 165600 35000
rect 165500 35000 165600 35100
rect 165600 26300 165700 26400
rect 165600 26400 165700 26500
rect 165600 26500 165700 26600
rect 165600 26600 165700 26700
rect 165600 26700 165700 26800
rect 165600 26800 165700 26900
rect 165600 26900 165700 27000
rect 165600 27000 165700 27100
rect 165600 27100 165700 27200
rect 165600 27200 165700 27300
rect 165600 27300 165700 27400
rect 165600 27400 165700 27500
rect 165600 27500 165700 27600
rect 165600 27600 165700 27700
rect 165600 27700 165700 27800
rect 165600 27800 165700 27900
rect 165600 27900 165700 28000
rect 165600 28000 165700 28100
rect 165600 28100 165700 28200
rect 165600 28200 165700 28300
rect 165600 28300 165700 28400
rect 165600 28400 165700 28500
rect 165600 28500 165700 28600
rect 165600 28600 165700 28700
rect 165600 28700 165700 28800
rect 165600 28800 165700 28900
rect 165600 28900 165700 29000
rect 165600 29000 165700 29100
rect 165600 29100 165700 29200
rect 165600 29200 165700 29300
rect 165600 29300 165700 29400
rect 165600 29400 165700 29500
rect 165600 29500 165700 29600
rect 165600 29600 165700 29700
rect 165600 29700 165700 29800
rect 165600 29800 165700 29900
rect 165600 29900 165700 30000
rect 165600 30000 165700 30100
rect 165600 30100 165700 30200
rect 165600 30200 165700 30300
rect 165600 30300 165700 30400
rect 165600 30400 165700 30500
rect 165600 30500 165700 30600
rect 165600 30600 165700 30700
rect 165600 30700 165700 30800
rect 165600 30800 165700 30900
rect 165600 30900 165700 31000
rect 165600 31000 165700 31100
rect 165600 31100 165700 31200
rect 165600 31200 165700 31300
rect 165600 31300 165700 31400
rect 165600 31400 165700 31500
rect 165600 31500 165700 31600
rect 165600 31600 165700 31700
rect 165600 31700 165700 31800
rect 165600 31800 165700 31900
rect 165600 31900 165700 32000
rect 165600 32000 165700 32100
rect 165600 32100 165700 32200
rect 165600 32200 165700 32300
rect 165600 32300 165700 32400
rect 165600 32400 165700 32500
rect 165600 32500 165700 32600
rect 165600 32600 165700 32700
rect 165600 32700 165700 32800
rect 165600 32800 165700 32900
rect 165600 32900 165700 33000
rect 165600 33000 165700 33100
rect 165600 33100 165700 33200
rect 165600 33200 165700 33300
rect 165600 33300 165700 33400
rect 165600 33400 165700 33500
rect 165600 33500 165700 33600
rect 165600 33600 165700 33700
rect 165600 33700 165700 33800
rect 165600 33800 165700 33900
rect 165600 33900 165700 34000
rect 165600 34000 165700 34100
rect 165600 34100 165700 34200
rect 165600 34200 165700 34300
rect 165600 34300 165700 34400
rect 165600 34400 165700 34500
rect 165600 34500 165700 34600
rect 165600 34600 165700 34700
rect 165600 34700 165700 34800
rect 165700 25800 165800 25900
rect 165700 25900 165800 26000
rect 165700 26000 165800 26100
rect 165700 26100 165800 26200
rect 165700 26200 165800 26300
rect 165700 26300 165800 26400
rect 165700 26400 165800 26500
rect 165700 26500 165800 26600
rect 165700 26600 165800 26700
rect 165700 26700 165800 26800
rect 165700 26800 165800 26900
rect 165700 26900 165800 27000
rect 165700 27000 165800 27100
rect 165700 27100 165800 27200
rect 165700 27200 165800 27300
rect 165700 27300 165800 27400
rect 165700 27400 165800 27500
rect 165700 27500 165800 27600
rect 165700 27600 165800 27700
rect 165700 27700 165800 27800
rect 165700 27800 165800 27900
rect 165700 27900 165800 28000
rect 165700 28000 165800 28100
rect 165700 28100 165800 28200
rect 165700 28200 165800 28300
rect 165700 28300 165800 28400
rect 165700 28400 165800 28500
rect 165700 28500 165800 28600
rect 165700 28600 165800 28700
rect 165700 28700 165800 28800
rect 165700 28800 165800 28900
rect 165700 28900 165800 29000
rect 165700 29000 165800 29100
rect 165700 29100 165800 29200
rect 165700 29200 165800 29300
rect 165700 29300 165800 29400
rect 165700 29400 165800 29500
rect 165700 29500 165800 29600
rect 165700 29600 165800 29700
rect 165700 29700 165800 29800
rect 165700 29800 165800 29900
rect 165700 29900 165800 30000
rect 165700 30000 165800 30100
rect 165700 30100 165800 30200
rect 165700 30200 165800 30300
rect 165700 30300 165800 30400
rect 165700 30400 165800 30500
rect 165700 30500 165800 30600
rect 165700 30600 165800 30700
rect 165700 30700 165800 30800
rect 165700 30800 165800 30900
rect 165700 30900 165800 31000
rect 165700 31000 165800 31100
rect 165700 31100 165800 31200
rect 165700 31200 165800 31300
rect 165700 31300 165800 31400
rect 165700 31400 165800 31500
rect 165700 31500 165800 31600
rect 165700 31600 165800 31700
rect 165700 31700 165800 31800
rect 165700 31800 165800 31900
rect 165700 31900 165800 32000
rect 165700 32000 165800 32100
rect 165700 32100 165800 32200
rect 165700 32200 165800 32300
rect 165700 32300 165800 32400
rect 165700 32400 165800 32500
rect 165700 32500 165800 32600
rect 165700 32600 165800 32700
rect 165700 32700 165800 32800
rect 165700 32800 165800 32900
rect 165700 32900 165800 33000
rect 165700 33000 165800 33100
rect 165700 33100 165800 33200
rect 165700 33200 165800 33300
rect 165700 33300 165800 33400
rect 165700 33400 165800 33500
rect 165700 33500 165800 33600
rect 165700 33600 165800 33700
rect 165700 33700 165800 33800
rect 165700 33800 165800 33900
rect 165700 33900 165800 34000
rect 165700 34000 165800 34100
rect 165700 34100 165800 34200
rect 165700 34200 165800 34300
rect 165700 34300 165800 34400
rect 165700 34400 165800 34500
rect 165800 25400 165900 25500
rect 165800 25500 165900 25600
rect 165800 25600 165900 25700
rect 165800 25700 165900 25800
rect 165800 25800 165900 25900
rect 165800 25900 165900 26000
rect 165800 26000 165900 26100
rect 165800 26100 165900 26200
rect 165800 26200 165900 26300
rect 165800 26300 165900 26400
rect 165800 26400 165900 26500
rect 165800 26500 165900 26600
rect 165800 26600 165900 26700
rect 165800 26700 165900 26800
rect 165800 26800 165900 26900
rect 165800 26900 165900 27000
rect 165800 27000 165900 27100
rect 165800 27100 165900 27200
rect 165800 27200 165900 27300
rect 165800 27300 165900 27400
rect 165800 27400 165900 27500
rect 165800 27500 165900 27600
rect 165800 27600 165900 27700
rect 165800 27700 165900 27800
rect 165800 27800 165900 27900
rect 165800 27900 165900 28000
rect 165800 28000 165900 28100
rect 165800 28100 165900 28200
rect 165800 28200 165900 28300
rect 165800 28300 165900 28400
rect 165800 28400 165900 28500
rect 165800 28500 165900 28600
rect 165800 28600 165900 28700
rect 165800 28700 165900 28800
rect 165800 28800 165900 28900
rect 165800 28900 165900 29000
rect 165800 29000 165900 29100
rect 165800 29100 165900 29200
rect 165800 29200 165900 29300
rect 165800 29300 165900 29400
rect 165800 29400 165900 29500
rect 165800 29500 165900 29600
rect 165800 29600 165900 29700
rect 165800 29700 165900 29800
rect 165800 29800 165900 29900
rect 165800 29900 165900 30000
rect 165800 30000 165900 30100
rect 165800 30100 165900 30200
rect 165800 30200 165900 30300
rect 165800 30300 165900 30400
rect 165800 30400 165900 30500
rect 165800 30500 165900 30600
rect 165800 30600 165900 30700
rect 165800 30700 165900 30800
rect 165800 30800 165900 30900
rect 165800 30900 165900 31000
rect 165800 31000 165900 31100
rect 165800 31100 165900 31200
rect 165800 31200 165900 31300
rect 165800 31300 165900 31400
rect 165800 31400 165900 31500
rect 165800 31500 165900 31600
rect 165800 31600 165900 31700
rect 165800 31700 165900 31800
rect 165800 31800 165900 31900
rect 165800 31900 165900 32000
rect 165800 32000 165900 32100
rect 165800 32100 165900 32200
rect 165800 32200 165900 32300
rect 165800 32300 165900 32400
rect 165800 32400 165900 32500
rect 165800 32500 165900 32600
rect 165800 32600 165900 32700
rect 165800 32700 165900 32800
rect 165800 32800 165900 32900
rect 165800 32900 165900 33000
rect 165800 33000 165900 33100
rect 165800 33100 165900 33200
rect 165800 33200 165900 33300
rect 165800 33300 165900 33400
rect 165800 33400 165900 33500
rect 165800 33500 165900 33600
rect 165800 33600 165900 33700
rect 165800 33700 165900 33800
rect 165800 33800 165900 33900
rect 165800 33900 165900 34000
rect 165800 34000 165900 34100
rect 165900 24900 166000 25000
rect 165900 25000 166000 25100
rect 165900 25100 166000 25200
rect 165900 25200 166000 25300
rect 165900 25300 166000 25400
rect 165900 25400 166000 25500
rect 165900 25500 166000 25600
rect 165900 25600 166000 25700
rect 165900 25700 166000 25800
rect 165900 25800 166000 25900
rect 165900 25900 166000 26000
rect 165900 26000 166000 26100
rect 165900 26100 166000 26200
rect 165900 26200 166000 26300
rect 165900 26300 166000 26400
rect 165900 26400 166000 26500
rect 165900 26500 166000 26600
rect 165900 26600 166000 26700
rect 165900 26700 166000 26800
rect 165900 26800 166000 26900
rect 165900 26900 166000 27000
rect 165900 27000 166000 27100
rect 165900 27100 166000 27200
rect 165900 27200 166000 27300
rect 165900 27300 166000 27400
rect 165900 27400 166000 27500
rect 165900 27500 166000 27600
rect 165900 27600 166000 27700
rect 165900 27700 166000 27800
rect 165900 27800 166000 27900
rect 165900 27900 166000 28000
rect 165900 28000 166000 28100
rect 165900 28100 166000 28200
rect 165900 28200 166000 28300
rect 165900 28300 166000 28400
rect 165900 28400 166000 28500
rect 165900 28500 166000 28600
rect 165900 28600 166000 28700
rect 165900 28700 166000 28800
rect 165900 28800 166000 28900
rect 165900 28900 166000 29000
rect 165900 29000 166000 29100
rect 165900 29100 166000 29200
rect 165900 29200 166000 29300
rect 165900 29300 166000 29400
rect 165900 29400 166000 29500
rect 165900 29500 166000 29600
rect 165900 29600 166000 29700
rect 165900 29700 166000 29800
rect 165900 29800 166000 29900
rect 165900 29900 166000 30000
rect 165900 30000 166000 30100
rect 165900 30100 166000 30200
rect 165900 30200 166000 30300
rect 165900 30300 166000 30400
rect 165900 30400 166000 30500
rect 165900 30500 166000 30600
rect 165900 30600 166000 30700
rect 165900 30700 166000 30800
rect 165900 30800 166000 30900
rect 165900 30900 166000 31000
rect 165900 31000 166000 31100
rect 165900 31100 166000 31200
rect 165900 31200 166000 31300
rect 165900 31300 166000 31400
rect 165900 31400 166000 31500
rect 165900 31500 166000 31600
rect 165900 31600 166000 31700
rect 165900 31700 166000 31800
rect 165900 31800 166000 31900
rect 165900 31900 166000 32000
rect 165900 32000 166000 32100
rect 165900 32100 166000 32200
rect 165900 32200 166000 32300
rect 165900 32300 166000 32400
rect 165900 32400 166000 32500
rect 165900 32500 166000 32600
rect 165900 32600 166000 32700
rect 165900 32700 166000 32800
rect 165900 32800 166000 32900
rect 165900 32900 166000 33000
rect 165900 33000 166000 33100
rect 165900 33100 166000 33200
rect 165900 33200 166000 33300
rect 165900 33300 166000 33400
rect 165900 33400 166000 33500
rect 165900 33500 166000 33600
rect 165900 33600 166000 33700
rect 165900 33700 166000 33800
rect 166000 24500 166100 24600
rect 166000 24600 166100 24700
rect 166000 24700 166100 24800
rect 166000 24800 166100 24900
rect 166000 24900 166100 25000
rect 166000 25000 166100 25100
rect 166000 25100 166100 25200
rect 166000 25200 166100 25300
rect 166000 25300 166100 25400
rect 166000 25400 166100 25500
rect 166000 25500 166100 25600
rect 166000 25600 166100 25700
rect 166000 25700 166100 25800
rect 166000 25800 166100 25900
rect 166000 25900 166100 26000
rect 166000 26000 166100 26100
rect 166000 26100 166100 26200
rect 166000 26200 166100 26300
rect 166000 26300 166100 26400
rect 166000 26400 166100 26500
rect 166000 26500 166100 26600
rect 166000 26600 166100 26700
rect 166000 26700 166100 26800
rect 166000 26800 166100 26900
rect 166000 26900 166100 27000
rect 166000 27000 166100 27100
rect 166000 27100 166100 27200
rect 166000 27200 166100 27300
rect 166000 27300 166100 27400
rect 166000 27400 166100 27500
rect 166000 27500 166100 27600
rect 166000 27600 166100 27700
rect 166000 27700 166100 27800
rect 166000 27800 166100 27900
rect 166000 27900 166100 28000
rect 166000 28000 166100 28100
rect 166000 28100 166100 28200
rect 166000 28200 166100 28300
rect 166000 28300 166100 28400
rect 166000 28400 166100 28500
rect 166000 28500 166100 28600
rect 166000 28600 166100 28700
rect 166000 28700 166100 28800
rect 166000 28800 166100 28900
rect 166000 28900 166100 29000
rect 166000 29000 166100 29100
rect 166000 29100 166100 29200
rect 166000 29200 166100 29300
rect 166000 29300 166100 29400
rect 166000 29400 166100 29500
rect 166000 29500 166100 29600
rect 166000 29600 166100 29700
rect 166000 29700 166100 29800
rect 166000 29800 166100 29900
rect 166000 29900 166100 30000
rect 166000 30000 166100 30100
rect 166000 30100 166100 30200
rect 166000 30200 166100 30300
rect 166000 30300 166100 30400
rect 166000 30400 166100 30500
rect 166000 30500 166100 30600
rect 166000 30600 166100 30700
rect 166000 30700 166100 30800
rect 166000 30800 166100 30900
rect 166000 30900 166100 31000
rect 166000 31000 166100 31100
rect 166000 31100 166100 31200
rect 166000 31200 166100 31300
rect 166000 31300 166100 31400
rect 166000 31400 166100 31500
rect 166000 31500 166100 31600
rect 166000 31600 166100 31700
rect 166000 31700 166100 31800
rect 166000 31800 166100 31900
rect 166000 31900 166100 32000
rect 166000 32000 166100 32100
rect 166000 32100 166100 32200
rect 166000 32200 166100 32300
rect 166000 32300 166100 32400
rect 166000 32400 166100 32500
rect 166000 32500 166100 32600
rect 166000 32600 166100 32700
rect 166000 32700 166100 32800
rect 166000 32800 166100 32900
rect 166000 32900 166100 33000
rect 166000 33000 166100 33100
rect 166000 33100 166100 33200
rect 166000 33200 166100 33300
rect 166000 33300 166100 33400
rect 166100 24100 166200 24200
rect 166100 24200 166200 24300
rect 166100 24300 166200 24400
rect 166100 24400 166200 24500
rect 166100 24500 166200 24600
rect 166100 24600 166200 24700
rect 166100 24700 166200 24800
rect 166100 24800 166200 24900
rect 166100 24900 166200 25000
rect 166100 25000 166200 25100
rect 166100 25100 166200 25200
rect 166100 25200 166200 25300
rect 166100 25300 166200 25400
rect 166100 25400 166200 25500
rect 166100 25500 166200 25600
rect 166100 25600 166200 25700
rect 166100 25700 166200 25800
rect 166100 25800 166200 25900
rect 166100 25900 166200 26000
rect 166100 26000 166200 26100
rect 166100 26100 166200 26200
rect 166100 26200 166200 26300
rect 166100 26300 166200 26400
rect 166100 26400 166200 26500
rect 166100 26500 166200 26600
rect 166100 26600 166200 26700
rect 166100 26700 166200 26800
rect 166100 26800 166200 26900
rect 166100 26900 166200 27000
rect 166100 27000 166200 27100
rect 166100 27100 166200 27200
rect 166100 27200 166200 27300
rect 166100 27300 166200 27400
rect 166100 27400 166200 27500
rect 166100 27500 166200 27600
rect 166100 27600 166200 27700
rect 166100 27700 166200 27800
rect 166100 27800 166200 27900
rect 166100 27900 166200 28000
rect 166100 28000 166200 28100
rect 166100 28100 166200 28200
rect 166100 28200 166200 28300
rect 166100 28300 166200 28400
rect 166100 28400 166200 28500
rect 166100 28500 166200 28600
rect 166100 28600 166200 28700
rect 166100 28700 166200 28800
rect 166100 28800 166200 28900
rect 166100 28900 166200 29000
rect 166100 29000 166200 29100
rect 166100 29100 166200 29200
rect 166100 29200 166200 29300
rect 166100 29300 166200 29400
rect 166100 29400 166200 29500
rect 166100 29500 166200 29600
rect 166100 29600 166200 29700
rect 166100 29700 166200 29800
rect 166100 29800 166200 29900
rect 166100 29900 166200 30000
rect 166100 30000 166200 30100
rect 166100 30100 166200 30200
rect 166100 30200 166200 30300
rect 166100 30300 166200 30400
rect 166100 30400 166200 30500
rect 166100 30500 166200 30600
rect 166100 30600 166200 30700
rect 166100 30700 166200 30800
rect 166100 30800 166200 30900
rect 166100 30900 166200 31000
rect 166100 31000 166200 31100
rect 166100 31100 166200 31200
rect 166100 31200 166200 31300
rect 166100 31300 166200 31400
rect 166100 31400 166200 31500
rect 166100 31500 166200 31600
rect 166100 31600 166200 31700
rect 166100 31700 166200 31800
rect 166100 31800 166200 31900
rect 166100 31900 166200 32000
rect 166100 32000 166200 32100
rect 166100 32100 166200 32200
rect 166100 32200 166200 32300
rect 166100 32300 166200 32400
rect 166100 32400 166200 32500
rect 166100 32500 166200 32600
rect 166100 32600 166200 32700
rect 166100 32700 166200 32800
rect 166100 32800 166200 32900
rect 166100 32900 166200 33000
rect 166100 33000 166200 33100
rect 166200 23600 166300 23700
rect 166200 23700 166300 23800
rect 166200 23800 166300 23900
rect 166200 23900 166300 24000
rect 166200 24000 166300 24100
rect 166200 24100 166300 24200
rect 166200 24200 166300 24300
rect 166200 24300 166300 24400
rect 166200 24400 166300 24500
rect 166200 24500 166300 24600
rect 166200 24600 166300 24700
rect 166200 24700 166300 24800
rect 166200 24800 166300 24900
rect 166200 24900 166300 25000
rect 166200 25000 166300 25100
rect 166200 25100 166300 25200
rect 166200 25200 166300 25300
rect 166200 25300 166300 25400
rect 166200 25400 166300 25500
rect 166200 25500 166300 25600
rect 166200 25600 166300 25700
rect 166200 25700 166300 25800
rect 166200 25800 166300 25900
rect 166200 25900 166300 26000
rect 166200 26000 166300 26100
rect 166200 26100 166300 26200
rect 166200 26200 166300 26300
rect 166200 26300 166300 26400
rect 166200 26400 166300 26500
rect 166200 26500 166300 26600
rect 166200 26600 166300 26700
rect 166200 26700 166300 26800
rect 166200 26800 166300 26900
rect 166200 26900 166300 27000
rect 166200 27000 166300 27100
rect 166200 27100 166300 27200
rect 166200 27200 166300 27300
rect 166200 27300 166300 27400
rect 166200 27400 166300 27500
rect 166200 27500 166300 27600
rect 166200 27600 166300 27700
rect 166200 27700 166300 27800
rect 166200 27800 166300 27900
rect 166200 27900 166300 28000
rect 166200 28000 166300 28100
rect 166200 28100 166300 28200
rect 166200 28200 166300 28300
rect 166200 28300 166300 28400
rect 166200 28400 166300 28500
rect 166200 28500 166300 28600
rect 166200 28600 166300 28700
rect 166200 28700 166300 28800
rect 166200 28800 166300 28900
rect 166200 28900 166300 29000
rect 166200 29000 166300 29100
rect 166200 29100 166300 29200
rect 166200 29200 166300 29300
rect 166200 29300 166300 29400
rect 166200 29400 166300 29500
rect 166200 29500 166300 29600
rect 166200 29600 166300 29700
rect 166200 29700 166300 29800
rect 166200 29800 166300 29900
rect 166200 29900 166300 30000
rect 166200 30000 166300 30100
rect 166200 30100 166300 30200
rect 166200 30200 166300 30300
rect 166200 30300 166300 30400
rect 166200 30400 166300 30500
rect 166200 30500 166300 30600
rect 166200 30600 166300 30700
rect 166200 30700 166300 30800
rect 166200 30800 166300 30900
rect 166200 30900 166300 31000
rect 166200 31000 166300 31100
rect 166200 31100 166300 31200
rect 166200 31200 166300 31300
rect 166200 31300 166300 31400
rect 166200 31400 166300 31500
rect 166200 31500 166300 31600
rect 166200 31600 166300 31700
rect 166200 31700 166300 31800
rect 166200 31800 166300 31900
rect 166200 31900 166300 32000
rect 166200 32000 166300 32100
rect 166200 32100 166300 32200
rect 166200 32200 166300 32300
rect 166200 32300 166300 32400
rect 166200 32400 166300 32500
rect 166200 32500 166300 32600
rect 166200 32600 166300 32700
rect 166300 23200 166400 23300
rect 166300 23300 166400 23400
rect 166300 23400 166400 23500
rect 166300 23500 166400 23600
rect 166300 23600 166400 23700
rect 166300 23700 166400 23800
rect 166300 23800 166400 23900
rect 166300 23900 166400 24000
rect 166300 24000 166400 24100
rect 166300 24100 166400 24200
rect 166300 24200 166400 24300
rect 166300 24300 166400 24400
rect 166300 24400 166400 24500
rect 166300 24500 166400 24600
rect 166300 24600 166400 24700
rect 166300 24700 166400 24800
rect 166300 24800 166400 24900
rect 166300 24900 166400 25000
rect 166300 25000 166400 25100
rect 166300 25100 166400 25200
rect 166300 25200 166400 25300
rect 166300 25300 166400 25400
rect 166300 25400 166400 25500
rect 166300 25500 166400 25600
rect 166300 25600 166400 25700
rect 166300 25700 166400 25800
rect 166300 25800 166400 25900
rect 166300 25900 166400 26000
rect 166300 26000 166400 26100
rect 166300 26100 166400 26200
rect 166300 26200 166400 26300
rect 166300 26300 166400 26400
rect 166300 26400 166400 26500
rect 166300 26500 166400 26600
rect 166300 26600 166400 26700
rect 166300 26700 166400 26800
rect 166300 26800 166400 26900
rect 166300 26900 166400 27000
rect 166300 27000 166400 27100
rect 166300 27100 166400 27200
rect 166300 27200 166400 27300
rect 166300 27300 166400 27400
rect 166300 27400 166400 27500
rect 166300 27500 166400 27600
rect 166300 27600 166400 27700
rect 166300 27700 166400 27800
rect 166300 27800 166400 27900
rect 166300 27900 166400 28000
rect 166300 28000 166400 28100
rect 166300 28100 166400 28200
rect 166300 28200 166400 28300
rect 166300 28300 166400 28400
rect 166300 28400 166400 28500
rect 166300 28500 166400 28600
rect 166300 28600 166400 28700
rect 166300 28700 166400 28800
rect 166300 28800 166400 28900
rect 166300 28900 166400 29000
rect 166300 29000 166400 29100
rect 166300 29100 166400 29200
rect 166300 29200 166400 29300
rect 166300 29300 166400 29400
rect 166300 29400 166400 29500
rect 166300 29500 166400 29600
rect 166300 29600 166400 29700
rect 166300 29700 166400 29800
rect 166300 29800 166400 29900
rect 166300 29900 166400 30000
rect 166300 30000 166400 30100
rect 166300 30100 166400 30200
rect 166300 30200 166400 30300
rect 166300 30300 166400 30400
rect 166300 30400 166400 30500
rect 166300 30500 166400 30600
rect 166300 30600 166400 30700
rect 166300 30700 166400 30800
rect 166300 30800 166400 30900
rect 166300 30900 166400 31000
rect 166300 31000 166400 31100
rect 166300 31100 166400 31200
rect 166300 31200 166400 31300
rect 166300 31300 166400 31400
rect 166300 31400 166400 31500
rect 166300 31500 166400 31600
rect 166300 31600 166400 31700
rect 166300 31700 166400 31800
rect 166300 31800 166400 31900
rect 166300 31900 166400 32000
rect 166300 32000 166400 32100
rect 166300 32100 166400 32200
rect 166300 32200 166400 32300
rect 166400 22600 166500 22700
rect 166400 22700 166500 22800
rect 166400 22800 166500 22900
rect 166400 22900 166500 23000
rect 166400 23000 166500 23100
rect 166400 23100 166500 23200
rect 166400 23200 166500 23300
rect 166400 23300 166500 23400
rect 166400 23400 166500 23500
rect 166400 23500 166500 23600
rect 166400 23600 166500 23700
rect 166400 23700 166500 23800
rect 166400 23800 166500 23900
rect 166400 23900 166500 24000
rect 166400 24000 166500 24100
rect 166400 24100 166500 24200
rect 166400 24200 166500 24300
rect 166400 24300 166500 24400
rect 166400 24400 166500 24500
rect 166400 24500 166500 24600
rect 166400 24600 166500 24700
rect 166400 24700 166500 24800
rect 166400 24800 166500 24900
rect 166400 24900 166500 25000
rect 166400 25000 166500 25100
rect 166400 25100 166500 25200
rect 166400 25200 166500 25300
rect 166400 25300 166500 25400
rect 166400 25400 166500 25500
rect 166400 25500 166500 25600
rect 166400 25600 166500 25700
rect 166400 25700 166500 25800
rect 166400 25800 166500 25900
rect 166400 25900 166500 26000
rect 166400 26000 166500 26100
rect 166400 26100 166500 26200
rect 166400 26200 166500 26300
rect 166400 26300 166500 26400
rect 166400 26400 166500 26500
rect 166400 26500 166500 26600
rect 166400 26600 166500 26700
rect 166400 26700 166500 26800
rect 166400 26800 166500 26900
rect 166400 26900 166500 27000
rect 166400 27000 166500 27100
rect 166400 27100 166500 27200
rect 166400 27200 166500 27300
rect 166400 27300 166500 27400
rect 166400 27400 166500 27500
rect 166400 27500 166500 27600
rect 166400 27600 166500 27700
rect 166400 27700 166500 27800
rect 166400 27800 166500 27900
rect 166400 27900 166500 28000
rect 166400 28000 166500 28100
rect 166400 28100 166500 28200
rect 166400 28200 166500 28300
rect 166400 28300 166500 28400
rect 166400 28400 166500 28500
rect 166400 28500 166500 28600
rect 166400 28600 166500 28700
rect 166400 28700 166500 28800
rect 166400 28800 166500 28900
rect 166400 28900 166500 29000
rect 166400 29000 166500 29100
rect 166400 29100 166500 29200
rect 166400 29200 166500 29300
rect 166400 29300 166500 29400
rect 166400 29400 166500 29500
rect 166400 29500 166500 29600
rect 166400 29600 166500 29700
rect 166400 29700 166500 29800
rect 166400 29800 166500 29900
rect 166400 29900 166500 30000
rect 166400 30000 166500 30100
rect 166400 30100 166500 30200
rect 166400 30200 166500 30300
rect 166400 30300 166500 30400
rect 166400 30400 166500 30500
rect 166400 30500 166500 30600
rect 166400 30600 166500 30700
rect 166400 30700 166500 30800
rect 166400 30800 166500 30900
rect 166400 30900 166500 31000
rect 166400 31000 166500 31100
rect 166400 31100 166500 31200
rect 166400 31200 166500 31300
rect 166400 31300 166500 31400
rect 166400 31400 166500 31500
rect 166400 31500 166500 31600
rect 166400 31600 166500 31700
rect 166400 31700 166500 31800
rect 166400 31800 166500 31900
rect 166500 22300 166600 22400
rect 166500 22400 166600 22500
rect 166500 22500 166600 22600
rect 166500 22600 166600 22700
rect 166500 22700 166600 22800
rect 166500 22800 166600 22900
rect 166500 22900 166600 23000
rect 166500 23000 166600 23100
rect 166500 23100 166600 23200
rect 166500 23200 166600 23300
rect 166500 23300 166600 23400
rect 166500 23400 166600 23500
rect 166500 23500 166600 23600
rect 166500 23600 166600 23700
rect 166500 23700 166600 23800
rect 166500 23800 166600 23900
rect 166500 23900 166600 24000
rect 166500 24000 166600 24100
rect 166500 24100 166600 24200
rect 166500 24200 166600 24300
rect 166500 24300 166600 24400
rect 166500 24400 166600 24500
rect 166500 24500 166600 24600
rect 166500 24600 166600 24700
rect 166500 24700 166600 24800
rect 166500 24800 166600 24900
rect 166500 24900 166600 25000
rect 166500 25000 166600 25100
rect 166500 25100 166600 25200
rect 166500 25200 166600 25300
rect 166500 25300 166600 25400
rect 166500 25400 166600 25500
rect 166500 25500 166600 25600
rect 166500 25600 166600 25700
rect 166500 25700 166600 25800
rect 166500 25800 166600 25900
rect 166500 25900 166600 26000
rect 166500 26000 166600 26100
rect 166500 26100 166600 26200
rect 166500 26200 166600 26300
rect 166500 26300 166600 26400
rect 166500 26400 166600 26500
rect 166500 26500 166600 26600
rect 166500 26600 166600 26700
rect 166500 26700 166600 26800
rect 166500 26800 166600 26900
rect 166500 26900 166600 27000
rect 166500 27000 166600 27100
rect 166500 27100 166600 27200
rect 166500 27200 166600 27300
rect 166500 27300 166600 27400
rect 166500 27400 166600 27500
rect 166500 27500 166600 27600
rect 166500 27600 166600 27700
rect 166500 27700 166600 27800
rect 166500 27800 166600 27900
rect 166500 27900 166600 28000
rect 166500 28000 166600 28100
rect 166500 28100 166600 28200
rect 166500 28200 166600 28300
rect 166500 28300 166600 28400
rect 166500 28400 166600 28500
rect 166500 28500 166600 28600
rect 166500 28600 166600 28700
rect 166500 28700 166600 28800
rect 166500 28800 166600 28900
rect 166500 28900 166600 29000
rect 166500 29000 166600 29100
rect 166500 29100 166600 29200
rect 166500 29200 166600 29300
rect 166500 29300 166600 29400
rect 166500 29400 166600 29500
rect 166500 29500 166600 29600
rect 166500 29600 166600 29700
rect 166500 29700 166600 29800
rect 166500 29800 166600 29900
rect 166500 29900 166600 30000
rect 166500 30000 166600 30100
rect 166500 30100 166600 30200
rect 166500 30200 166600 30300
rect 166500 30300 166600 30400
rect 166500 30400 166600 30500
rect 166500 30500 166600 30600
rect 166500 30600 166600 30700
rect 166500 30700 166600 30800
rect 166500 30800 166600 30900
rect 166500 30900 166600 31000
rect 166500 31000 166600 31100
rect 166500 31100 166600 31200
rect 166500 31200 166600 31300
rect 166500 31300 166600 31400
rect 166500 31400 166600 31500
rect 166600 22200 166700 22300
rect 166600 22300 166700 22400
rect 166600 22400 166700 22500
rect 166600 22500 166700 22600
rect 166600 22600 166700 22700
rect 166600 22700 166700 22800
rect 166600 22800 166700 22900
rect 166600 22900 166700 23000
rect 166600 23000 166700 23100
rect 166600 23100 166700 23200
rect 166600 23200 166700 23300
rect 166600 23300 166700 23400
rect 166600 23400 166700 23500
rect 166600 23500 166700 23600
rect 166600 23600 166700 23700
rect 166600 23700 166700 23800
rect 166600 23800 166700 23900
rect 166600 23900 166700 24000
rect 166600 24000 166700 24100
rect 166600 24100 166700 24200
rect 166600 24200 166700 24300
rect 166600 24300 166700 24400
rect 166600 24400 166700 24500
rect 166600 24500 166700 24600
rect 166600 24600 166700 24700
rect 166600 24700 166700 24800
rect 166600 24800 166700 24900
rect 166600 24900 166700 25000
rect 166600 25000 166700 25100
rect 166600 25100 166700 25200
rect 166600 25200 166700 25300
rect 166600 25300 166700 25400
rect 166600 25400 166700 25500
rect 166600 25500 166700 25600
rect 166600 25600 166700 25700
rect 166600 25700 166700 25800
rect 166600 25800 166700 25900
rect 166600 25900 166700 26000
rect 166600 26000 166700 26100
rect 166600 26100 166700 26200
rect 166600 26200 166700 26300
rect 166600 26300 166700 26400
rect 166600 26400 166700 26500
rect 166600 26500 166700 26600
rect 166600 26600 166700 26700
rect 166600 26700 166700 26800
rect 166600 26800 166700 26900
rect 166600 26900 166700 27000
rect 166600 27000 166700 27100
rect 166600 27100 166700 27200
rect 166600 27200 166700 27300
rect 166600 27300 166700 27400
rect 166600 27400 166700 27500
rect 166600 27500 166700 27600
rect 166600 27600 166700 27700
rect 166600 27700 166700 27800
rect 166600 27800 166700 27900
rect 166600 27900 166700 28000
rect 166600 28000 166700 28100
rect 166600 28100 166700 28200
rect 166600 28200 166700 28300
rect 166600 28300 166700 28400
rect 166600 28400 166700 28500
rect 166600 28500 166700 28600
rect 166600 28600 166700 28700
rect 166600 28700 166700 28800
rect 166600 28800 166700 28900
rect 166600 28900 166700 29000
rect 166600 29000 166700 29100
rect 166600 29100 166700 29200
rect 166600 29200 166700 29300
rect 166600 29300 166700 29400
rect 166600 29400 166700 29500
rect 166600 29500 166700 29600
rect 166600 29600 166700 29700
rect 166600 29700 166700 29800
rect 166600 29800 166700 29900
rect 166600 29900 166700 30000
rect 166600 30000 166700 30100
rect 166600 30100 166700 30200
rect 166600 30200 166700 30300
rect 166600 30300 166700 30400
rect 166600 30400 166700 30500
rect 166600 30500 166700 30600
rect 166600 30600 166700 30700
rect 166600 30700 166700 30800
rect 166600 30800 166700 30900
rect 166600 30900 166700 31000
rect 166700 22000 166800 22100
rect 166700 22100 166800 22200
rect 166700 22200 166800 22300
rect 166700 22300 166800 22400
rect 166700 22400 166800 22500
rect 166700 22500 166800 22600
rect 166700 22600 166800 22700
rect 166700 22700 166800 22800
rect 166700 22800 166800 22900
rect 166700 22900 166800 23000
rect 166700 23000 166800 23100
rect 166700 23100 166800 23200
rect 166700 23200 166800 23300
rect 166700 23300 166800 23400
rect 166700 23400 166800 23500
rect 166700 23500 166800 23600
rect 166700 23600 166800 23700
rect 166700 23700 166800 23800
rect 166700 23800 166800 23900
rect 166700 23900 166800 24000
rect 166700 24000 166800 24100
rect 166700 24100 166800 24200
rect 166700 24200 166800 24300
rect 166700 24300 166800 24400
rect 166700 24400 166800 24500
rect 166700 24500 166800 24600
rect 166700 24600 166800 24700
rect 166700 24700 166800 24800
rect 166700 24800 166800 24900
rect 166700 24900 166800 25000
rect 166700 25000 166800 25100
rect 166700 25100 166800 25200
rect 166700 25200 166800 25300
rect 166700 25300 166800 25400
rect 166700 25400 166800 25500
rect 166700 25500 166800 25600
rect 166700 25600 166800 25700
rect 166700 25700 166800 25800
rect 166700 25800 166800 25900
rect 166700 25900 166800 26000
rect 166700 26000 166800 26100
rect 166700 26100 166800 26200
rect 166700 26200 166800 26300
rect 166700 26300 166800 26400
rect 166700 26400 166800 26500
rect 166700 26500 166800 26600
rect 166700 26600 166800 26700
rect 166700 26700 166800 26800
rect 166700 26800 166800 26900
rect 166700 26900 166800 27000
rect 166700 27000 166800 27100
rect 166700 27100 166800 27200
rect 166700 27200 166800 27300
rect 166700 27300 166800 27400
rect 166700 27400 166800 27500
rect 166700 27500 166800 27600
rect 166700 27600 166800 27700
rect 166700 27700 166800 27800
rect 166700 27800 166800 27900
rect 166700 27900 166800 28000
rect 166700 28000 166800 28100
rect 166700 28100 166800 28200
rect 166700 28200 166800 28300
rect 166700 28300 166800 28400
rect 166700 28400 166800 28500
rect 166700 28500 166800 28600
rect 166700 28600 166800 28700
rect 166700 28700 166800 28800
rect 166700 28800 166800 28900
rect 166700 28900 166800 29000
rect 166700 29000 166800 29100
rect 166700 29100 166800 29200
rect 166700 29200 166800 29300
rect 166700 29300 166800 29400
rect 166700 29400 166800 29500
rect 166700 29500 166800 29600
rect 166700 29600 166800 29700
rect 166700 29700 166800 29800
rect 166700 29800 166800 29900
rect 166700 29900 166800 30000
rect 166700 30000 166800 30100
rect 166700 30100 166800 30200
rect 166700 30200 166800 30300
rect 166700 30300 166800 30400
rect 166700 30400 166800 30500
rect 166700 30500 166800 30600
rect 166800 22000 166900 22100
rect 166800 22100 166900 22200
rect 166800 22200 166900 22300
rect 166800 22300 166900 22400
rect 166800 22400 166900 22500
rect 166800 22500 166900 22600
rect 166800 22600 166900 22700
rect 166800 22700 166900 22800
rect 166800 22800 166900 22900
rect 166800 22900 166900 23000
rect 166800 23000 166900 23100
rect 166800 23100 166900 23200
rect 166800 23200 166900 23300
rect 166800 23300 166900 23400
rect 166800 23400 166900 23500
rect 166800 23500 166900 23600
rect 166800 23600 166900 23700
rect 166800 23700 166900 23800
rect 166800 23800 166900 23900
rect 166800 23900 166900 24000
rect 166800 24000 166900 24100
rect 166800 24100 166900 24200
rect 166800 24200 166900 24300
rect 166800 24300 166900 24400
rect 166800 24400 166900 24500
rect 166800 24500 166900 24600
rect 166800 24600 166900 24700
rect 166800 24700 166900 24800
rect 166800 24800 166900 24900
rect 166800 24900 166900 25000
rect 166800 25000 166900 25100
rect 166800 25100 166900 25200
rect 166800 25200 166900 25300
rect 166800 25300 166900 25400
rect 166800 25400 166900 25500
rect 166800 25500 166900 25600
rect 166800 25600 166900 25700
rect 166800 25700 166900 25800
rect 166800 25800 166900 25900
rect 166800 25900 166900 26000
rect 166800 26000 166900 26100
rect 166800 26100 166900 26200
rect 166800 26200 166900 26300
rect 166800 26300 166900 26400
rect 166800 26400 166900 26500
rect 166800 26500 166900 26600
rect 166800 26600 166900 26700
rect 166800 26700 166900 26800
rect 166800 26800 166900 26900
rect 166800 26900 166900 27000
rect 166800 27000 166900 27100
rect 166800 27100 166900 27200
rect 166800 27200 166900 27300
rect 166800 27300 166900 27400
rect 166800 27400 166900 27500
rect 166800 27500 166900 27600
rect 166800 27600 166900 27700
rect 166800 27700 166900 27800
rect 166800 27800 166900 27900
rect 166800 27900 166900 28000
rect 166800 28000 166900 28100
rect 166800 28100 166900 28200
rect 166800 28200 166900 28300
rect 166800 28300 166900 28400
rect 166800 28400 166900 28500
rect 166800 28500 166900 28600
rect 166800 28600 166900 28700
rect 166800 28700 166900 28800
rect 166800 28800 166900 28900
rect 166800 28900 166900 29000
rect 166800 29000 166900 29100
rect 166800 29100 166900 29200
rect 166800 29200 166900 29300
rect 166800 29300 166900 29400
rect 166800 29400 166900 29500
rect 166800 29500 166900 29600
rect 166800 29600 166900 29700
rect 166800 29700 166900 29800
rect 166800 29800 166900 29900
rect 166800 29900 166900 30000
rect 166800 30000 166900 30100
rect 166800 30100 166900 30200
rect 166900 21900 167000 22000
rect 166900 22000 167000 22100
rect 166900 22100 167000 22200
rect 166900 22200 167000 22300
rect 166900 22300 167000 22400
rect 166900 22400 167000 22500
rect 166900 22500 167000 22600
rect 166900 22600 167000 22700
rect 166900 22700 167000 22800
rect 166900 22800 167000 22900
rect 166900 22900 167000 23000
rect 166900 23000 167000 23100
rect 166900 23100 167000 23200
rect 166900 23200 167000 23300
rect 166900 23300 167000 23400
rect 166900 23400 167000 23500
rect 166900 23500 167000 23600
rect 166900 23600 167000 23700
rect 166900 23700 167000 23800
rect 166900 23800 167000 23900
rect 166900 23900 167000 24000
rect 166900 24000 167000 24100
rect 166900 24100 167000 24200
rect 166900 24200 167000 24300
rect 166900 24300 167000 24400
rect 166900 24400 167000 24500
rect 166900 24500 167000 24600
rect 166900 24600 167000 24700
rect 166900 24700 167000 24800
rect 166900 24800 167000 24900
rect 166900 24900 167000 25000
rect 166900 25000 167000 25100
rect 166900 25100 167000 25200
rect 166900 25200 167000 25300
rect 166900 25300 167000 25400
rect 166900 25400 167000 25500
rect 166900 25500 167000 25600
rect 166900 25600 167000 25700
rect 166900 25700 167000 25800
rect 166900 25800 167000 25900
rect 166900 25900 167000 26000
rect 166900 26000 167000 26100
rect 166900 26100 167000 26200
rect 166900 26200 167000 26300
rect 166900 26300 167000 26400
rect 166900 26400 167000 26500
rect 166900 26500 167000 26600
rect 166900 26600 167000 26700
rect 166900 26700 167000 26800
rect 166900 26800 167000 26900
rect 166900 26900 167000 27000
rect 166900 27000 167000 27100
rect 166900 27100 167000 27200
rect 166900 27200 167000 27300
rect 166900 27300 167000 27400
rect 166900 27400 167000 27500
rect 166900 27500 167000 27600
rect 166900 27600 167000 27700
rect 166900 27700 167000 27800
rect 166900 27800 167000 27900
rect 166900 27900 167000 28000
rect 166900 28000 167000 28100
rect 166900 28100 167000 28200
rect 166900 28200 167000 28300
rect 166900 28300 167000 28400
rect 166900 28400 167000 28500
rect 166900 28500 167000 28600
rect 166900 28600 167000 28700
rect 166900 28700 167000 28800
rect 166900 28800 167000 28900
rect 166900 28900 167000 29000
rect 166900 29000 167000 29100
rect 166900 29100 167000 29200
rect 166900 29200 167000 29300
rect 166900 29300 167000 29400
rect 166900 29400 167000 29500
rect 166900 29500 167000 29600
rect 166900 29600 167000 29700
rect 167000 21800 167100 21900
rect 167000 21900 167100 22000
rect 167000 22000 167100 22100
rect 167000 22100 167100 22200
rect 167000 22200 167100 22300
rect 167000 22300 167100 22400
rect 167000 22400 167100 22500
rect 167000 22500 167100 22600
rect 167000 22600 167100 22700
rect 167000 22700 167100 22800
rect 167000 22800 167100 22900
rect 167000 22900 167100 23000
rect 167000 23000 167100 23100
rect 167000 23100 167100 23200
rect 167000 23200 167100 23300
rect 167000 23300 167100 23400
rect 167000 23400 167100 23500
rect 167000 23500 167100 23600
rect 167000 23600 167100 23700
rect 167000 23700 167100 23800
rect 167000 23800 167100 23900
rect 167000 23900 167100 24000
rect 167000 24000 167100 24100
rect 167000 24100 167100 24200
rect 167000 24200 167100 24300
rect 167000 24300 167100 24400
rect 167000 24400 167100 24500
rect 167000 24500 167100 24600
rect 167000 24600 167100 24700
rect 167000 24700 167100 24800
rect 167000 24800 167100 24900
rect 167000 24900 167100 25000
rect 167000 25000 167100 25100
rect 167000 25100 167100 25200
rect 167000 25200 167100 25300
rect 167000 25300 167100 25400
rect 167000 25400 167100 25500
rect 167000 25500 167100 25600
rect 167000 25600 167100 25700
rect 167000 25700 167100 25800
rect 167000 25800 167100 25900
rect 167000 25900 167100 26000
rect 167000 26000 167100 26100
rect 167000 26100 167100 26200
rect 167000 26200 167100 26300
rect 167000 26300 167100 26400
rect 167000 26400 167100 26500
rect 167000 26500 167100 26600
rect 167000 26600 167100 26700
rect 167000 26700 167100 26800
rect 167000 26800 167100 26900
rect 167000 26900 167100 27000
rect 167000 27000 167100 27100
rect 167000 27100 167100 27200
rect 167000 27200 167100 27300
rect 167000 27300 167100 27400
rect 167000 27400 167100 27500
rect 167000 27500 167100 27600
rect 167000 27600 167100 27700
rect 167000 27700 167100 27800
rect 167000 27800 167100 27900
rect 167000 27900 167100 28000
rect 167000 28000 167100 28100
rect 167000 28100 167100 28200
rect 167000 28200 167100 28300
rect 167000 28300 167100 28400
rect 167000 28400 167100 28500
rect 167000 28500 167100 28600
rect 167000 28600 167100 28700
rect 167000 28700 167100 28800
rect 167000 28800 167100 28900
rect 167000 28900 167100 29000
rect 167000 29000 167100 29100
rect 167000 29100 167100 29200
rect 167100 21800 167200 21900
rect 167100 21900 167200 22000
rect 167100 22000 167200 22100
rect 167100 22100 167200 22200
rect 167100 22200 167200 22300
rect 167100 22300 167200 22400
rect 167100 22400 167200 22500
rect 167100 22500 167200 22600
rect 167100 22600 167200 22700
rect 167100 22700 167200 22800
rect 167100 22800 167200 22900
rect 167100 22900 167200 23000
rect 167100 23000 167200 23100
rect 167100 23100 167200 23200
rect 167100 23200 167200 23300
rect 167100 23300 167200 23400
rect 167100 23400 167200 23500
rect 167100 23500 167200 23600
rect 167100 23600 167200 23700
rect 167100 23700 167200 23800
rect 167100 23800 167200 23900
rect 167100 23900 167200 24000
rect 167100 24000 167200 24100
rect 167100 24100 167200 24200
rect 167100 24200 167200 24300
rect 167100 24300 167200 24400
rect 167100 24400 167200 24500
rect 167100 24500 167200 24600
rect 167100 24600 167200 24700
rect 167100 24700 167200 24800
rect 167100 24800 167200 24900
rect 167100 24900 167200 25000
rect 167100 25000 167200 25100
rect 167100 25100 167200 25200
rect 167100 25200 167200 25300
rect 167100 25300 167200 25400
rect 167100 25400 167200 25500
rect 167100 25500 167200 25600
rect 167100 25600 167200 25700
rect 167100 25700 167200 25800
rect 167100 25800 167200 25900
rect 167100 25900 167200 26000
rect 167100 26000 167200 26100
rect 167100 26100 167200 26200
rect 167100 26200 167200 26300
rect 167100 26300 167200 26400
rect 167100 26400 167200 26500
rect 167100 26500 167200 26600
rect 167100 26600 167200 26700
rect 167100 26700 167200 26800
rect 167100 26800 167200 26900
rect 167100 26900 167200 27000
rect 167100 27000 167200 27100
rect 167100 27100 167200 27200
rect 167100 27200 167200 27300
rect 167100 27300 167200 27400
rect 167100 27400 167200 27500
rect 167100 27500 167200 27600
rect 167100 27600 167200 27700
rect 167100 27700 167200 27800
rect 167100 27800 167200 27900
rect 167100 27900 167200 28000
rect 167100 28000 167200 28100
rect 167100 28100 167200 28200
rect 167100 28200 167200 28300
rect 167100 28300 167200 28400
rect 167100 28400 167200 28500
rect 167100 28500 167200 28600
rect 167100 28600 167200 28700
rect 167100 28700 167200 28800
rect 167200 21800 167300 21900
rect 167200 21900 167300 22000
rect 167200 22000 167300 22100
rect 167200 22100 167300 22200
rect 167200 22200 167300 22300
rect 167200 22300 167300 22400
rect 167200 22400 167300 22500
rect 167200 22500 167300 22600
rect 167200 22600 167300 22700
rect 167200 22700 167300 22800
rect 167200 22800 167300 22900
rect 167200 22900 167300 23000
rect 167200 23000 167300 23100
rect 167200 23100 167300 23200
rect 167200 23200 167300 23300
rect 167200 23300 167300 23400
rect 167200 23400 167300 23500
rect 167200 23500 167300 23600
rect 167200 23600 167300 23700
rect 167200 23700 167300 23800
rect 167200 23800 167300 23900
rect 167200 23900 167300 24000
rect 167200 24000 167300 24100
rect 167200 24100 167300 24200
rect 167200 24200 167300 24300
rect 167200 24300 167300 24400
rect 167200 24400 167300 24500
rect 167200 24500 167300 24600
rect 167200 24600 167300 24700
rect 167200 24700 167300 24800
rect 167200 24800 167300 24900
rect 167200 24900 167300 25000
rect 167200 25000 167300 25100
rect 167200 25100 167300 25200
rect 167200 25200 167300 25300
rect 167200 25300 167300 25400
rect 167200 25400 167300 25500
rect 167200 25500 167300 25600
rect 167200 25600 167300 25700
rect 167200 25700 167300 25800
rect 167200 25800 167300 25900
rect 167200 25900 167300 26000
rect 167200 26000 167300 26100
rect 167200 26100 167300 26200
rect 167200 26200 167300 26300
rect 167200 26300 167300 26400
rect 167200 26400 167300 26500
rect 167200 26500 167300 26600
rect 167200 26600 167300 26700
rect 167200 26700 167300 26800
rect 167200 26800 167300 26900
rect 167200 26900 167300 27000
rect 167200 27000 167300 27100
rect 167200 27100 167300 27200
rect 167200 27200 167300 27300
rect 167200 27300 167300 27400
rect 167200 27400 167300 27500
rect 167200 27500 167300 27600
rect 167200 27600 167300 27700
rect 167200 27700 167300 27800
rect 167200 27800 167300 27900
rect 167200 27900 167300 28000
rect 167200 28000 167300 28100
rect 167200 28100 167300 28200
rect 167200 28200 167300 28300
rect 167300 21800 167400 21900
rect 167300 21900 167400 22000
rect 167300 22000 167400 22100
rect 167300 22100 167400 22200
rect 167300 22200 167400 22300
rect 167300 22300 167400 22400
rect 167300 22400 167400 22500
rect 167300 22500 167400 22600
rect 167300 22600 167400 22700
rect 167300 22700 167400 22800
rect 167300 22800 167400 22900
rect 167300 22900 167400 23000
rect 167300 23000 167400 23100
rect 167300 23100 167400 23200
rect 167300 23200 167400 23300
rect 167300 23300 167400 23400
rect 167300 23400 167400 23500
rect 167300 23500 167400 23600
rect 167300 23600 167400 23700
rect 167300 23700 167400 23800
rect 167300 23800 167400 23900
rect 167300 23900 167400 24000
rect 167300 24000 167400 24100
rect 167300 24100 167400 24200
rect 167300 24200 167400 24300
rect 167300 24300 167400 24400
rect 167300 24400 167400 24500
rect 167300 24500 167400 24600
rect 167300 24600 167400 24700
rect 167300 24700 167400 24800
rect 167300 24800 167400 24900
rect 167300 24900 167400 25000
rect 167300 25000 167400 25100
rect 167300 25100 167400 25200
rect 167300 25200 167400 25300
rect 167300 25300 167400 25400
rect 167300 25400 167400 25500
rect 167300 25500 167400 25600
rect 167300 25600 167400 25700
rect 167300 25700 167400 25800
rect 167300 25800 167400 25900
rect 167300 25900 167400 26000
rect 167300 26000 167400 26100
rect 167300 26100 167400 26200
rect 167300 26200 167400 26300
rect 167300 26300 167400 26400
rect 167300 26400 167400 26500
rect 167300 26500 167400 26600
rect 167300 26600 167400 26700
rect 167300 26700 167400 26800
rect 167300 26800 167400 26900
rect 167300 26900 167400 27000
rect 167300 27000 167400 27100
rect 167300 27100 167400 27200
rect 167300 27200 167400 27300
rect 167300 27300 167400 27400
rect 167300 27400 167400 27500
rect 167300 27500 167400 27600
rect 167300 27600 167400 27700
rect 167300 27700 167400 27800
rect 167300 27800 167400 27900
rect 167400 21700 167500 21800
rect 167400 21800 167500 21900
rect 167400 21900 167500 22000
rect 167400 22000 167500 22100
rect 167400 22100 167500 22200
rect 167400 22200 167500 22300
rect 167400 22300 167500 22400
rect 167400 22400 167500 22500
rect 167400 22500 167500 22600
rect 167400 22600 167500 22700
rect 167400 22700 167500 22800
rect 167400 22800 167500 22900
rect 167400 22900 167500 23000
rect 167400 23000 167500 23100
rect 167400 23100 167500 23200
rect 167400 23200 167500 23300
rect 167400 23300 167500 23400
rect 167400 23400 167500 23500
rect 167400 23500 167500 23600
rect 167400 23600 167500 23700
rect 167400 23700 167500 23800
rect 167400 23800 167500 23900
rect 167400 23900 167500 24000
rect 167400 24000 167500 24100
rect 167400 24100 167500 24200
rect 167400 24200 167500 24300
rect 167400 24300 167500 24400
rect 167400 24400 167500 24500
rect 167400 24500 167500 24600
rect 167400 24600 167500 24700
rect 167400 24700 167500 24800
rect 167400 24800 167500 24900
rect 167400 24900 167500 25000
rect 167400 25000 167500 25100
rect 167400 25100 167500 25200
rect 167400 25200 167500 25300
rect 167400 25300 167500 25400
rect 167400 25400 167500 25500
rect 167400 25500 167500 25600
rect 167400 25600 167500 25700
rect 167400 25700 167500 25800
rect 167400 25800 167500 25900
rect 167400 25900 167500 26000
rect 167400 26000 167500 26100
rect 167400 26100 167500 26200
rect 167400 26200 167500 26300
rect 167400 26300 167500 26400
rect 167400 26400 167500 26500
rect 167400 26500 167500 26600
rect 167400 26600 167500 26700
rect 167400 26700 167500 26800
rect 167400 26800 167500 26900
rect 167400 26900 167500 27000
rect 167400 27000 167500 27100
rect 167400 27100 167500 27200
rect 167400 27200 167500 27300
rect 167400 27300 167500 27400
rect 167500 21700 167600 21800
rect 167500 21800 167600 21900
rect 167500 21900 167600 22000
rect 167500 22000 167600 22100
rect 167500 22100 167600 22200
rect 167500 22200 167600 22300
rect 167500 22300 167600 22400
rect 167500 22400 167600 22500
rect 167500 22500 167600 22600
rect 167500 22600 167600 22700
rect 167500 22700 167600 22800
rect 167500 22800 167600 22900
rect 167500 22900 167600 23000
rect 167500 23000 167600 23100
rect 167500 23100 167600 23200
rect 167500 23200 167600 23300
rect 167500 23300 167600 23400
rect 167500 23400 167600 23500
rect 167500 23500 167600 23600
rect 167500 23600 167600 23700
rect 167500 23700 167600 23800
rect 167500 23800 167600 23900
rect 167500 23900 167600 24000
rect 167500 24000 167600 24100
rect 167500 24100 167600 24200
rect 167500 24200 167600 24300
rect 167500 24300 167600 24400
rect 167500 24400 167600 24500
rect 167500 24500 167600 24600
rect 167500 24600 167600 24700
rect 167500 24700 167600 24800
rect 167500 24800 167600 24900
rect 167500 24900 167600 25000
rect 167500 25000 167600 25100
rect 167500 25100 167600 25200
rect 167500 25200 167600 25300
rect 167500 25300 167600 25400
rect 167500 25400 167600 25500
rect 167500 25500 167600 25600
rect 167500 25600 167600 25700
rect 167500 25700 167600 25800
rect 167500 25800 167600 25900
rect 167500 25900 167600 26000
rect 167500 26000 167600 26100
rect 167500 26100 167600 26200
rect 167500 26200 167600 26300
rect 167500 26300 167600 26400
rect 167500 26400 167600 26500
rect 167500 26500 167600 26600
rect 167500 26600 167600 26700
rect 167500 26700 167600 26800
rect 167500 26800 167600 26900
rect 167500 26900 167600 27000
rect 167600 21700 167700 21800
rect 167600 21800 167700 21900
rect 167600 21900 167700 22000
rect 167600 22000 167700 22100
rect 167600 22100 167700 22200
rect 167600 22200 167700 22300
rect 167600 22300 167700 22400
rect 167600 22400 167700 22500
rect 167600 22500 167700 22600
rect 167600 22600 167700 22700
rect 167600 22700 167700 22800
rect 167600 22800 167700 22900
rect 167600 22900 167700 23000
rect 167600 23000 167700 23100
rect 167600 23100 167700 23200
rect 167600 23200 167700 23300
rect 167600 23300 167700 23400
rect 167600 23400 167700 23500
rect 167600 23500 167700 23600
rect 167600 23600 167700 23700
rect 167600 23700 167700 23800
rect 167600 23800 167700 23900
rect 167600 23900 167700 24000
rect 167600 24000 167700 24100
rect 167600 24100 167700 24200
rect 167600 24200 167700 24300
rect 167600 24300 167700 24400
rect 167600 24400 167700 24500
rect 167600 24500 167700 24600
rect 167600 24600 167700 24700
rect 167600 24700 167700 24800
rect 167600 24800 167700 24900
rect 167600 24900 167700 25000
rect 167600 25000 167700 25100
rect 167600 25100 167700 25200
rect 167600 25200 167700 25300
rect 167600 25300 167700 25400
rect 167600 25400 167700 25500
rect 167600 25500 167700 25600
rect 167600 25600 167700 25700
rect 167600 25700 167700 25800
rect 167600 25800 167700 25900
rect 167600 25900 167700 26000
rect 167600 26000 167700 26100
rect 167600 26100 167700 26200
rect 167600 26200 167700 26300
rect 167600 26300 167700 26400
rect 167600 26400 167700 26500
rect 167700 21700 167800 21800
rect 167700 21800 167800 21900
rect 167700 21900 167800 22000
rect 167700 22000 167800 22100
rect 167700 22100 167800 22200
rect 167700 22200 167800 22300
rect 167700 22300 167800 22400
rect 167700 22400 167800 22500
rect 167700 22500 167800 22600
rect 167700 22600 167800 22700
rect 167700 22700 167800 22800
rect 167700 22800 167800 22900
rect 167700 22900 167800 23000
rect 167700 23000 167800 23100
rect 167700 23100 167800 23200
rect 167700 23200 167800 23300
rect 167700 23300 167800 23400
rect 167700 23400 167800 23500
rect 167700 23500 167800 23600
rect 167700 23600 167800 23700
rect 167700 23700 167800 23800
rect 167700 23800 167800 23900
rect 167700 23900 167800 24000
rect 167700 24000 167800 24100
rect 167700 24100 167800 24200
rect 167700 24200 167800 24300
rect 167700 24300 167800 24400
rect 167700 24400 167800 24500
rect 167700 24500 167800 24600
rect 167700 24600 167800 24700
rect 167700 24700 167800 24800
rect 167700 24800 167800 24900
rect 167700 24900 167800 25000
rect 167700 25000 167800 25100
rect 167700 25100 167800 25200
rect 167700 25200 167800 25300
rect 167700 25300 167800 25400
rect 167700 25400 167800 25500
rect 167700 25500 167800 25600
rect 167700 25600 167800 25700
rect 167700 25700 167800 25800
rect 167700 25800 167800 25900
rect 167700 25900 167800 26000
rect 167700 26000 167800 26100
rect 167700 26100 167800 26200
rect 167700 26200 167800 26300
rect 167800 21700 167900 21800
rect 167800 21800 167900 21900
rect 167800 21900 167900 22000
rect 167800 22000 167900 22100
rect 167800 22100 167900 22200
rect 167800 22200 167900 22300
rect 167800 22300 167900 22400
rect 167800 22400 167900 22500
rect 167800 22500 167900 22600
rect 167800 22600 167900 22700
rect 167800 22700 167900 22800
rect 167800 22800 167900 22900
rect 167800 22900 167900 23000
rect 167800 23000 167900 23100
rect 167800 23100 167900 23200
rect 167800 23200 167900 23300
rect 167800 23300 167900 23400
rect 167800 23400 167900 23500
rect 167800 23500 167900 23600
rect 167800 23600 167900 23700
rect 167800 23700 167900 23800
rect 167800 23800 167900 23900
rect 167800 23900 167900 24000
rect 167800 24000 167900 24100
rect 167800 24100 167900 24200
rect 167800 24200 167900 24300
rect 167800 24300 167900 24400
rect 167800 24400 167900 24500
rect 167800 24500 167900 24600
rect 167800 24600 167900 24700
rect 167800 24700 167900 24800
rect 167800 24800 167900 24900
rect 167800 24900 167900 25000
rect 167800 25000 167900 25100
rect 167800 25100 167900 25200
rect 167800 25200 167900 25300
rect 167800 25300 167900 25400
rect 167800 25400 167900 25500
rect 167800 25500 167900 25600
rect 167800 25600 167900 25700
rect 167800 25700 167900 25800
rect 167800 25800 167900 25900
rect 167800 25900 167900 26000
rect 167800 26000 167900 26100
rect 167800 26100 167900 26200
rect 167800 26200 167900 26300
rect 167800 26300 167900 26400
rect 167800 26400 167900 26500
rect 167900 21700 168000 21800
rect 167900 21800 168000 21900
rect 167900 21900 168000 22000
rect 167900 22000 168000 22100
rect 167900 22100 168000 22200
rect 167900 22200 168000 22300
rect 167900 22300 168000 22400
rect 167900 22400 168000 22500
rect 167900 22500 168000 22600
rect 167900 22600 168000 22700
rect 167900 22700 168000 22800
rect 167900 22800 168000 22900
rect 167900 22900 168000 23000
rect 167900 23000 168000 23100
rect 167900 23100 168000 23200
rect 167900 23200 168000 23300
rect 167900 23300 168000 23400
rect 167900 23400 168000 23500
rect 167900 23500 168000 23600
rect 167900 23600 168000 23700
rect 167900 23700 168000 23800
rect 167900 23800 168000 23900
rect 167900 23900 168000 24000
rect 167900 24000 168000 24100
rect 167900 24100 168000 24200
rect 167900 24200 168000 24300
rect 167900 24300 168000 24400
rect 167900 24400 168000 24500
rect 167900 24500 168000 24600
rect 167900 24600 168000 24700
rect 167900 24700 168000 24800
rect 167900 24800 168000 24900
rect 167900 24900 168000 25000
rect 167900 25000 168000 25100
rect 167900 25100 168000 25200
rect 167900 25200 168000 25300
rect 167900 25300 168000 25400
rect 167900 25400 168000 25500
rect 167900 25500 168000 25600
rect 167900 25600 168000 25700
rect 167900 25700 168000 25800
rect 167900 25800 168000 25900
rect 167900 25900 168000 26000
rect 167900 26000 168000 26100
rect 167900 26100 168000 26200
rect 167900 26200 168000 26300
rect 167900 26300 168000 26400
rect 167900 26400 168000 26500
rect 167900 26500 168000 26600
rect 167900 26600 168000 26700
rect 167900 26700 168000 26800
rect 168000 21700 168100 21800
rect 168000 21800 168100 21900
rect 168000 21900 168100 22000
rect 168000 22000 168100 22100
rect 168000 22100 168100 22200
rect 168000 22200 168100 22300
rect 168000 22300 168100 22400
rect 168000 22400 168100 22500
rect 168000 22500 168100 22600
rect 168000 22600 168100 22700
rect 168000 22700 168100 22800
rect 168000 22800 168100 22900
rect 168000 22900 168100 23000
rect 168000 23000 168100 23100
rect 168000 23100 168100 23200
rect 168000 23200 168100 23300
rect 168000 23300 168100 23400
rect 168000 23400 168100 23500
rect 168000 23500 168100 23600
rect 168000 23600 168100 23700
rect 168000 23700 168100 23800
rect 168000 23800 168100 23900
rect 168000 23900 168100 24000
rect 168000 24000 168100 24100
rect 168000 24100 168100 24200
rect 168000 24200 168100 24300
rect 168000 24300 168100 24400
rect 168000 24400 168100 24500
rect 168000 24500 168100 24600
rect 168000 24600 168100 24700
rect 168000 24700 168100 24800
rect 168000 24800 168100 24900
rect 168000 24900 168100 25000
rect 168000 25000 168100 25100
rect 168000 25100 168100 25200
rect 168000 25200 168100 25300
rect 168000 25300 168100 25400
rect 168000 25400 168100 25500
rect 168000 25500 168100 25600
rect 168000 25600 168100 25700
rect 168000 25700 168100 25800
rect 168000 25800 168100 25900
rect 168000 25900 168100 26000
rect 168000 26000 168100 26100
rect 168000 26100 168100 26200
rect 168000 26200 168100 26300
rect 168000 26300 168100 26400
rect 168000 26400 168100 26500
rect 168000 26500 168100 26600
rect 168000 26600 168100 26700
rect 168000 26700 168100 26800
rect 168000 26800 168100 26900
rect 168000 26900 168100 27000
rect 168100 21700 168200 21800
rect 168100 21800 168200 21900
rect 168100 21900 168200 22000
rect 168100 22000 168200 22100
rect 168100 22100 168200 22200
rect 168100 22200 168200 22300
rect 168100 22300 168200 22400
rect 168100 22400 168200 22500
rect 168100 22500 168200 22600
rect 168100 22600 168200 22700
rect 168100 22700 168200 22800
rect 168100 22800 168200 22900
rect 168100 22900 168200 23000
rect 168100 23000 168200 23100
rect 168100 23100 168200 23200
rect 168100 23200 168200 23300
rect 168100 23300 168200 23400
rect 168100 23400 168200 23500
rect 168100 23500 168200 23600
rect 168100 23600 168200 23700
rect 168100 23700 168200 23800
rect 168100 23800 168200 23900
rect 168100 23900 168200 24000
rect 168100 24000 168200 24100
rect 168100 24100 168200 24200
rect 168100 24200 168200 24300
rect 168100 24300 168200 24400
rect 168100 24400 168200 24500
rect 168100 24500 168200 24600
rect 168100 24600 168200 24700
rect 168100 24700 168200 24800
rect 168100 24800 168200 24900
rect 168100 24900 168200 25000
rect 168100 25000 168200 25100
rect 168100 25100 168200 25200
rect 168100 25200 168200 25300
rect 168100 25300 168200 25400
rect 168100 25400 168200 25500
rect 168100 25500 168200 25600
rect 168100 25600 168200 25700
rect 168100 25700 168200 25800
rect 168100 25800 168200 25900
rect 168100 25900 168200 26000
rect 168100 26000 168200 26100
rect 168100 26100 168200 26200
rect 168100 26200 168200 26300
rect 168100 26300 168200 26400
rect 168100 26400 168200 26500
rect 168100 26500 168200 26600
rect 168100 26600 168200 26700
rect 168100 26700 168200 26800
rect 168100 26800 168200 26900
rect 168100 26900 168200 27000
rect 168100 27000 168200 27100
rect 168100 27100 168200 27200
rect 168200 21800 168300 21900
rect 168200 21900 168300 22000
rect 168200 22000 168300 22100
rect 168200 22100 168300 22200
rect 168200 22200 168300 22300
rect 168200 22300 168300 22400
rect 168200 22400 168300 22500
rect 168200 22500 168300 22600
rect 168200 22600 168300 22700
rect 168200 22700 168300 22800
rect 168200 22800 168300 22900
rect 168200 22900 168300 23000
rect 168200 23000 168300 23100
rect 168200 23100 168300 23200
rect 168200 23200 168300 23300
rect 168200 23300 168300 23400
rect 168200 23400 168300 23500
rect 168200 23500 168300 23600
rect 168200 23600 168300 23700
rect 168200 23700 168300 23800
rect 168200 23800 168300 23900
rect 168200 23900 168300 24000
rect 168200 24000 168300 24100
rect 168200 24100 168300 24200
rect 168200 24200 168300 24300
rect 168200 24300 168300 24400
rect 168200 24400 168300 24500
rect 168200 24500 168300 24600
rect 168200 24600 168300 24700
rect 168200 24700 168300 24800
rect 168200 24800 168300 24900
rect 168200 24900 168300 25000
rect 168200 25000 168300 25100
rect 168200 25100 168300 25200
rect 168200 25200 168300 25300
rect 168200 25300 168300 25400
rect 168200 25400 168300 25500
rect 168200 25500 168300 25600
rect 168200 25600 168300 25700
rect 168200 25700 168300 25800
rect 168200 25800 168300 25900
rect 168200 25900 168300 26000
rect 168200 26000 168300 26100
rect 168200 26100 168300 26200
rect 168200 26200 168300 26300
rect 168200 26300 168300 26400
rect 168200 26400 168300 26500
rect 168200 26500 168300 26600
rect 168200 26600 168300 26700
rect 168200 26700 168300 26800
rect 168200 26800 168300 26900
rect 168200 26900 168300 27000
rect 168200 27000 168300 27100
rect 168200 27100 168300 27200
rect 168200 27200 168300 27300
rect 168200 27300 168300 27400
rect 168200 27400 168300 27500
rect 168300 21800 168400 21900
rect 168300 21900 168400 22000
rect 168300 22000 168400 22100
rect 168300 22100 168400 22200
rect 168300 22200 168400 22300
rect 168300 22300 168400 22400
rect 168300 22400 168400 22500
rect 168300 22500 168400 22600
rect 168300 22600 168400 22700
rect 168300 22700 168400 22800
rect 168300 22800 168400 22900
rect 168300 22900 168400 23000
rect 168300 23000 168400 23100
rect 168300 23100 168400 23200
rect 168300 23200 168400 23300
rect 168300 23300 168400 23400
rect 168300 23400 168400 23500
rect 168300 23500 168400 23600
rect 168300 23600 168400 23700
rect 168300 23700 168400 23800
rect 168300 23800 168400 23900
rect 168300 23900 168400 24000
rect 168300 24000 168400 24100
rect 168300 24100 168400 24200
rect 168300 24200 168400 24300
rect 168300 24300 168400 24400
rect 168300 24400 168400 24500
rect 168300 24500 168400 24600
rect 168300 24600 168400 24700
rect 168300 24700 168400 24800
rect 168300 24800 168400 24900
rect 168300 24900 168400 25000
rect 168300 25000 168400 25100
rect 168300 25100 168400 25200
rect 168300 25200 168400 25300
rect 168300 25300 168400 25400
rect 168300 25400 168400 25500
rect 168300 25500 168400 25600
rect 168300 25600 168400 25700
rect 168300 25700 168400 25800
rect 168300 25800 168400 25900
rect 168300 25900 168400 26000
rect 168300 26000 168400 26100
rect 168300 26100 168400 26200
rect 168300 26200 168400 26300
rect 168300 26300 168400 26400
rect 168300 26400 168400 26500
rect 168300 26500 168400 26600
rect 168300 26600 168400 26700
rect 168300 26700 168400 26800
rect 168300 26800 168400 26900
rect 168300 26900 168400 27000
rect 168300 27000 168400 27100
rect 168300 27100 168400 27200
rect 168300 27200 168400 27300
rect 168300 27300 168400 27400
rect 168300 27400 168400 27500
rect 168300 27500 168400 27600
rect 168300 27600 168400 27700
rect 168300 27700 168400 27800
rect 168400 21800 168500 21900
rect 168400 21900 168500 22000
rect 168400 22000 168500 22100
rect 168400 22100 168500 22200
rect 168400 22200 168500 22300
rect 168400 22300 168500 22400
rect 168400 22400 168500 22500
rect 168400 22500 168500 22600
rect 168400 22600 168500 22700
rect 168400 22700 168500 22800
rect 168400 22800 168500 22900
rect 168400 22900 168500 23000
rect 168400 23000 168500 23100
rect 168400 23100 168500 23200
rect 168400 23200 168500 23300
rect 168400 23300 168500 23400
rect 168400 23400 168500 23500
rect 168400 23500 168500 23600
rect 168400 23600 168500 23700
rect 168400 23700 168500 23800
rect 168400 23800 168500 23900
rect 168400 23900 168500 24000
rect 168400 24000 168500 24100
rect 168400 24100 168500 24200
rect 168400 24200 168500 24300
rect 168400 24300 168500 24400
rect 168400 24400 168500 24500
rect 168400 24500 168500 24600
rect 168400 24600 168500 24700
rect 168400 24700 168500 24800
rect 168400 24800 168500 24900
rect 168400 24900 168500 25000
rect 168400 25000 168500 25100
rect 168400 25100 168500 25200
rect 168400 25200 168500 25300
rect 168400 25300 168500 25400
rect 168400 25400 168500 25500
rect 168400 25500 168500 25600
rect 168400 25600 168500 25700
rect 168400 25700 168500 25800
rect 168400 25800 168500 25900
rect 168400 25900 168500 26000
rect 168400 26000 168500 26100
rect 168400 26100 168500 26200
rect 168400 26200 168500 26300
rect 168400 26300 168500 26400
rect 168400 26400 168500 26500
rect 168400 26500 168500 26600
rect 168400 26600 168500 26700
rect 168400 26700 168500 26800
rect 168400 26800 168500 26900
rect 168400 26900 168500 27000
rect 168400 27000 168500 27100
rect 168400 27100 168500 27200
rect 168400 27200 168500 27300
rect 168400 27300 168500 27400
rect 168400 27400 168500 27500
rect 168400 27500 168500 27600
rect 168400 27600 168500 27700
rect 168400 27700 168500 27800
rect 168400 27800 168500 27900
rect 168400 27900 168500 28000
rect 168500 21900 168600 22000
rect 168500 22000 168600 22100
rect 168500 22100 168600 22200
rect 168500 22200 168600 22300
rect 168500 22300 168600 22400
rect 168500 22400 168600 22500
rect 168500 22500 168600 22600
rect 168500 22600 168600 22700
rect 168500 22700 168600 22800
rect 168500 22800 168600 22900
rect 168500 22900 168600 23000
rect 168500 23000 168600 23100
rect 168500 23100 168600 23200
rect 168500 23200 168600 23300
rect 168500 23300 168600 23400
rect 168500 23400 168600 23500
rect 168500 23500 168600 23600
rect 168500 23600 168600 23700
rect 168500 23700 168600 23800
rect 168500 23800 168600 23900
rect 168500 23900 168600 24000
rect 168500 24000 168600 24100
rect 168500 24100 168600 24200
rect 168500 24200 168600 24300
rect 168500 24300 168600 24400
rect 168500 24400 168600 24500
rect 168500 24500 168600 24600
rect 168500 24600 168600 24700
rect 168500 24700 168600 24800
rect 168500 24800 168600 24900
rect 168500 24900 168600 25000
rect 168500 25000 168600 25100
rect 168500 25100 168600 25200
rect 168500 25200 168600 25300
rect 168500 25300 168600 25400
rect 168500 25400 168600 25500
rect 168500 25500 168600 25600
rect 168500 25600 168600 25700
rect 168500 25700 168600 25800
rect 168500 25800 168600 25900
rect 168500 25900 168600 26000
rect 168500 26000 168600 26100
rect 168500 26100 168600 26200
rect 168500 26200 168600 26300
rect 168500 26300 168600 26400
rect 168500 26400 168600 26500
rect 168500 26500 168600 26600
rect 168500 26600 168600 26700
rect 168500 26700 168600 26800
rect 168500 26800 168600 26900
rect 168500 26900 168600 27000
rect 168500 27000 168600 27100
rect 168500 27100 168600 27200
rect 168500 27200 168600 27300
rect 168500 27300 168600 27400
rect 168500 27400 168600 27500
rect 168500 27500 168600 27600
rect 168500 27600 168600 27700
rect 168500 27700 168600 27800
rect 168500 27800 168600 27900
rect 168500 27900 168600 28000
rect 168500 28000 168600 28100
rect 168500 28100 168600 28200
rect 168500 28200 168600 28300
rect 168600 22000 168700 22100
rect 168600 22100 168700 22200
rect 168600 22200 168700 22300
rect 168600 22300 168700 22400
rect 168600 22400 168700 22500
rect 168600 22500 168700 22600
rect 168600 22600 168700 22700
rect 168600 22700 168700 22800
rect 168600 22800 168700 22900
rect 168600 22900 168700 23000
rect 168600 23000 168700 23100
rect 168600 23100 168700 23200
rect 168600 23200 168700 23300
rect 168600 23300 168700 23400
rect 168600 23400 168700 23500
rect 168600 23500 168700 23600
rect 168600 23600 168700 23700
rect 168600 23700 168700 23800
rect 168600 23800 168700 23900
rect 168600 23900 168700 24000
rect 168600 24000 168700 24100
rect 168600 24100 168700 24200
rect 168600 24200 168700 24300
rect 168600 24300 168700 24400
rect 168600 24400 168700 24500
rect 168600 24500 168700 24600
rect 168600 24600 168700 24700
rect 168600 24700 168700 24800
rect 168600 24800 168700 24900
rect 168600 24900 168700 25000
rect 168600 25000 168700 25100
rect 168600 25100 168700 25200
rect 168600 25200 168700 25300
rect 168600 25300 168700 25400
rect 168600 25400 168700 25500
rect 168600 25500 168700 25600
rect 168600 25600 168700 25700
rect 168600 25700 168700 25800
rect 168600 25800 168700 25900
rect 168600 25900 168700 26000
rect 168600 26000 168700 26100
rect 168600 26100 168700 26200
rect 168600 26200 168700 26300
rect 168600 26300 168700 26400
rect 168600 26400 168700 26500
rect 168600 26500 168700 26600
rect 168600 26600 168700 26700
rect 168600 26700 168700 26800
rect 168600 26800 168700 26900
rect 168600 26900 168700 27000
rect 168600 27000 168700 27100
rect 168600 27100 168700 27200
rect 168600 27200 168700 27300
rect 168600 27300 168700 27400
rect 168600 27400 168700 27500
rect 168600 27500 168700 27600
rect 168600 27600 168700 27700
rect 168600 27700 168700 27800
rect 168600 27800 168700 27900
rect 168600 27900 168700 28000
rect 168600 28000 168700 28100
rect 168600 28100 168700 28200
rect 168600 28200 168700 28300
rect 168600 28300 168700 28400
rect 168600 28400 168700 28500
rect 168600 28500 168700 28600
rect 168700 22000 168800 22100
rect 168700 22100 168800 22200
rect 168700 22200 168800 22300
rect 168700 22300 168800 22400
rect 168700 22400 168800 22500
rect 168700 22500 168800 22600
rect 168700 22600 168800 22700
rect 168700 22700 168800 22800
rect 168700 22800 168800 22900
rect 168700 22900 168800 23000
rect 168700 23000 168800 23100
rect 168700 23100 168800 23200
rect 168700 23200 168800 23300
rect 168700 23300 168800 23400
rect 168700 23400 168800 23500
rect 168700 23500 168800 23600
rect 168700 23600 168800 23700
rect 168700 23700 168800 23800
rect 168700 23800 168800 23900
rect 168700 23900 168800 24000
rect 168700 24000 168800 24100
rect 168700 24100 168800 24200
rect 168700 24200 168800 24300
rect 168700 24300 168800 24400
rect 168700 24400 168800 24500
rect 168700 24500 168800 24600
rect 168700 24600 168800 24700
rect 168700 24700 168800 24800
rect 168700 24800 168800 24900
rect 168700 24900 168800 25000
rect 168700 25000 168800 25100
rect 168700 25100 168800 25200
rect 168700 25200 168800 25300
rect 168700 25300 168800 25400
rect 168700 25400 168800 25500
rect 168700 25500 168800 25600
rect 168700 25600 168800 25700
rect 168700 25700 168800 25800
rect 168700 25800 168800 25900
rect 168700 25900 168800 26000
rect 168700 26000 168800 26100
rect 168700 26100 168800 26200
rect 168700 26200 168800 26300
rect 168700 26300 168800 26400
rect 168700 26400 168800 26500
rect 168700 26500 168800 26600
rect 168700 26600 168800 26700
rect 168700 26700 168800 26800
rect 168700 26800 168800 26900
rect 168700 26900 168800 27000
rect 168700 27000 168800 27100
rect 168700 27100 168800 27200
rect 168700 27200 168800 27300
rect 168700 27300 168800 27400
rect 168700 27400 168800 27500
rect 168700 27500 168800 27600
rect 168700 27600 168800 27700
rect 168700 27700 168800 27800
rect 168700 27800 168800 27900
rect 168700 27900 168800 28000
rect 168700 28000 168800 28100
rect 168700 28100 168800 28200
rect 168700 28200 168800 28300
rect 168700 28300 168800 28400
rect 168700 28400 168800 28500
rect 168700 28500 168800 28600
rect 168700 28600 168800 28700
rect 168700 28700 168800 28800
rect 168800 22100 168900 22200
rect 168800 22200 168900 22300
rect 168800 22300 168900 22400
rect 168800 22400 168900 22500
rect 168800 22500 168900 22600
rect 168800 22600 168900 22700
rect 168800 22700 168900 22800
rect 168800 22800 168900 22900
rect 168800 22900 168900 23000
rect 168800 23000 168900 23100
rect 168800 23100 168900 23200
rect 168800 23200 168900 23300
rect 168800 23300 168900 23400
rect 168800 23400 168900 23500
rect 168800 23500 168900 23600
rect 168800 23600 168900 23700
rect 168800 23700 168900 23800
rect 168800 23800 168900 23900
rect 168800 23900 168900 24000
rect 168800 24000 168900 24100
rect 168800 24100 168900 24200
rect 168800 24200 168900 24300
rect 168800 24300 168900 24400
rect 168800 24400 168900 24500
rect 168800 24500 168900 24600
rect 168800 24600 168900 24700
rect 168800 24700 168900 24800
rect 168800 24800 168900 24900
rect 168800 24900 168900 25000
rect 168800 25000 168900 25100
rect 168800 25100 168900 25200
rect 168800 25200 168900 25300
rect 168800 25300 168900 25400
rect 168800 25400 168900 25500
rect 168800 25500 168900 25600
rect 168800 25600 168900 25700
rect 168800 25700 168900 25800
rect 168800 25800 168900 25900
rect 168800 25900 168900 26000
rect 168800 26000 168900 26100
rect 168800 26100 168900 26200
rect 168800 26200 168900 26300
rect 168800 26300 168900 26400
rect 168800 26400 168900 26500
rect 168800 26500 168900 26600
rect 168800 26600 168900 26700
rect 168800 26700 168900 26800
rect 168800 26800 168900 26900
rect 168800 26900 168900 27000
rect 168800 27000 168900 27100
rect 168800 27100 168900 27200
rect 168800 27200 168900 27300
rect 168800 27300 168900 27400
rect 168800 27400 168900 27500
rect 168800 27500 168900 27600
rect 168800 27600 168900 27700
rect 168800 27700 168900 27800
rect 168800 27800 168900 27900
rect 168800 27900 168900 28000
rect 168800 28000 168900 28100
rect 168800 28100 168900 28200
rect 168800 28200 168900 28300
rect 168800 28300 168900 28400
rect 168800 28400 168900 28500
rect 168800 28500 168900 28600
rect 168800 28600 168900 28700
rect 168800 28700 168900 28800
rect 168800 28800 168900 28900
rect 168800 28900 168900 29000
rect 168800 29000 168900 29100
rect 168900 22200 169000 22300
rect 168900 22300 169000 22400
rect 168900 22400 169000 22500
rect 168900 22500 169000 22600
rect 168900 22600 169000 22700
rect 168900 22700 169000 22800
rect 168900 22800 169000 22900
rect 168900 22900 169000 23000
rect 168900 23000 169000 23100
rect 168900 23100 169000 23200
rect 168900 23200 169000 23300
rect 168900 23300 169000 23400
rect 168900 23400 169000 23500
rect 168900 23500 169000 23600
rect 168900 23600 169000 23700
rect 168900 23700 169000 23800
rect 168900 23800 169000 23900
rect 168900 23900 169000 24000
rect 168900 24000 169000 24100
rect 168900 24100 169000 24200
rect 168900 24200 169000 24300
rect 168900 24300 169000 24400
rect 168900 24400 169000 24500
rect 168900 24500 169000 24600
rect 168900 24600 169000 24700
rect 168900 24700 169000 24800
rect 168900 24800 169000 24900
rect 168900 24900 169000 25000
rect 168900 25000 169000 25100
rect 168900 25100 169000 25200
rect 168900 25200 169000 25300
rect 168900 25300 169000 25400
rect 168900 25400 169000 25500
rect 168900 25500 169000 25600
rect 168900 25600 169000 25700
rect 168900 25700 169000 25800
rect 168900 25800 169000 25900
rect 168900 25900 169000 26000
rect 168900 26000 169000 26100
rect 168900 26100 169000 26200
rect 168900 26200 169000 26300
rect 168900 26300 169000 26400
rect 168900 26400 169000 26500
rect 168900 26500 169000 26600
rect 168900 26600 169000 26700
rect 168900 26700 169000 26800
rect 168900 26800 169000 26900
rect 168900 26900 169000 27000
rect 168900 27000 169000 27100
rect 168900 27100 169000 27200
rect 168900 27200 169000 27300
rect 168900 27300 169000 27400
rect 168900 27400 169000 27500
rect 168900 27500 169000 27600
rect 168900 27600 169000 27700
rect 168900 27700 169000 27800
rect 168900 27800 169000 27900
rect 168900 27900 169000 28000
rect 168900 28000 169000 28100
rect 168900 28100 169000 28200
rect 168900 28200 169000 28300
rect 168900 28300 169000 28400
rect 168900 28400 169000 28500
rect 168900 28500 169000 28600
rect 168900 28600 169000 28700
rect 168900 28700 169000 28800
rect 168900 28800 169000 28900
rect 168900 28900 169000 29000
rect 168900 29000 169000 29100
rect 168900 29100 169000 29200
rect 168900 29200 169000 29300
rect 168900 29300 169000 29400
rect 169000 22400 169100 22500
rect 169000 22500 169100 22600
rect 169000 22600 169100 22700
rect 169000 22700 169100 22800
rect 169000 22800 169100 22900
rect 169000 22900 169100 23000
rect 169000 23000 169100 23100
rect 169000 23500 169100 23600
rect 169000 23600 169100 23700
rect 169000 23700 169100 23800
rect 169000 23800 169100 23900
rect 169000 23900 169100 24000
rect 169000 24000 169100 24100
rect 169000 24100 169100 24200
rect 169000 24200 169100 24300
rect 169000 24300 169100 24400
rect 169000 24400 169100 24500
rect 169000 24500 169100 24600
rect 169000 24600 169100 24700
rect 169000 24700 169100 24800
rect 169000 24800 169100 24900
rect 169000 24900 169100 25000
rect 169000 25000 169100 25100
rect 169000 25100 169100 25200
rect 169000 25200 169100 25300
rect 169000 25300 169100 25400
rect 169000 25400 169100 25500
rect 169000 25500 169100 25600
rect 169000 25600 169100 25700
rect 169000 25700 169100 25800
rect 169000 25800 169100 25900
rect 169000 25900 169100 26000
rect 169000 26000 169100 26100
rect 169000 26100 169100 26200
rect 169000 26200 169100 26300
rect 169000 26300 169100 26400
rect 169000 26400 169100 26500
rect 169000 26500 169100 26600
rect 169000 26600 169100 26700
rect 169000 26700 169100 26800
rect 169000 26800 169100 26900
rect 169000 26900 169100 27000
rect 169000 27000 169100 27100
rect 169000 27100 169100 27200
rect 169000 27200 169100 27300
rect 169000 27300 169100 27400
rect 169000 27400 169100 27500
rect 169000 27500 169100 27600
rect 169000 27600 169100 27700
rect 169000 27700 169100 27800
rect 169000 27800 169100 27900
rect 169000 27900 169100 28000
rect 169000 28000 169100 28100
rect 169000 28100 169100 28200
rect 169000 28200 169100 28300
rect 169000 28300 169100 28400
rect 169000 28400 169100 28500
rect 169000 28500 169100 28600
rect 169000 28600 169100 28700
rect 169000 28700 169100 28800
rect 169000 28800 169100 28900
rect 169000 28900 169100 29000
rect 169000 29000 169100 29100
rect 169000 29100 169100 29200
rect 169000 29200 169100 29300
rect 169000 29300 169100 29400
rect 169000 29400 169100 29500
rect 169000 29500 169100 29600
rect 169000 29600 169100 29700
rect 169100 23800 169200 23900
rect 169100 23900 169200 24000
rect 169100 24000 169200 24100
rect 169100 24100 169200 24200
rect 169100 24200 169200 24300
rect 169100 24300 169200 24400
rect 169100 24400 169200 24500
rect 169100 24500 169200 24600
rect 169100 24600 169200 24700
rect 169100 24700 169200 24800
rect 169100 24800 169200 24900
rect 169100 24900 169200 25000
rect 169100 25000 169200 25100
rect 169100 25100 169200 25200
rect 169100 25200 169200 25300
rect 169100 25300 169200 25400
rect 169100 25400 169200 25500
rect 169100 25500 169200 25600
rect 169100 25600 169200 25700
rect 169100 25700 169200 25800
rect 169100 25800 169200 25900
rect 169100 25900 169200 26000
rect 169100 26000 169200 26100
rect 169100 26100 169200 26200
rect 169100 26200 169200 26300
rect 169100 26300 169200 26400
rect 169100 26400 169200 26500
rect 169100 26500 169200 26600
rect 169100 26600 169200 26700
rect 169100 26700 169200 26800
rect 169100 26800 169200 26900
rect 169100 26900 169200 27000
rect 169100 27000 169200 27100
rect 169100 27100 169200 27200
rect 169100 27200 169200 27300
rect 169100 27300 169200 27400
rect 169100 27400 169200 27500
rect 169100 27500 169200 27600
rect 169100 27600 169200 27700
rect 169100 27700 169200 27800
rect 169100 27800 169200 27900
rect 169100 27900 169200 28000
rect 169100 28000 169200 28100
rect 169100 28100 169200 28200
rect 169100 28200 169200 28300
rect 169100 28300 169200 28400
rect 169100 28400 169200 28500
rect 169100 28500 169200 28600
rect 169100 28600 169200 28700
rect 169100 28700 169200 28800
rect 169100 28800 169200 28900
rect 169100 28900 169200 29000
rect 169100 29000 169200 29100
rect 169100 29100 169200 29200
rect 169100 29200 169200 29300
rect 169100 29300 169200 29400
rect 169100 29400 169200 29500
rect 169100 29500 169200 29600
rect 169100 29600 169200 29700
rect 169100 29700 169200 29800
rect 169100 29800 169200 29900
rect 169100 29900 169200 30000
rect 169200 24200 169300 24300
rect 169200 24300 169300 24400
rect 169200 24400 169300 24500
rect 169200 24500 169300 24600
rect 169200 24600 169300 24700
rect 169200 24700 169300 24800
rect 169200 24800 169300 24900
rect 169200 24900 169300 25000
rect 169200 25000 169300 25100
rect 169200 25100 169300 25200
rect 169200 25200 169300 25300
rect 169200 25300 169300 25400
rect 169200 25400 169300 25500
rect 169200 25500 169300 25600
rect 169200 25600 169300 25700
rect 169200 25700 169300 25800
rect 169200 25800 169300 25900
rect 169200 25900 169300 26000
rect 169200 26000 169300 26100
rect 169200 26100 169300 26200
rect 169200 26200 169300 26300
rect 169200 26300 169300 26400
rect 169200 26400 169300 26500
rect 169200 26500 169300 26600
rect 169200 26600 169300 26700
rect 169200 26700 169300 26800
rect 169200 26800 169300 26900
rect 169200 26900 169300 27000
rect 169200 27000 169300 27100
rect 169200 27100 169300 27200
rect 169200 27200 169300 27300
rect 169200 27300 169300 27400
rect 169200 27400 169300 27500
rect 169200 27500 169300 27600
rect 169200 27600 169300 27700
rect 169200 27700 169300 27800
rect 169200 27800 169300 27900
rect 169200 27900 169300 28000
rect 169200 28000 169300 28100
rect 169200 28100 169300 28200
rect 169200 28200 169300 28300
rect 169200 28300 169300 28400
rect 169200 28400 169300 28500
rect 169200 28500 169300 28600
rect 169200 28600 169300 28700
rect 169200 28700 169300 28800
rect 169200 28800 169300 28900
rect 169200 28900 169300 29000
rect 169200 29000 169300 29100
rect 169200 29100 169300 29200
rect 169200 29200 169300 29300
rect 169200 29300 169300 29400
rect 169200 29400 169300 29500
rect 169200 29500 169300 29600
rect 169200 29600 169300 29700
rect 169200 29700 169300 29800
rect 169200 29800 169300 29900
rect 169200 29900 169300 30000
rect 169200 30000 169300 30100
rect 169200 30100 169300 30200
rect 169200 30200 169300 30300
rect 169300 24400 169400 24500
rect 169300 24500 169400 24600
rect 169300 24600 169400 24700
rect 169300 24700 169400 24800
rect 169300 24800 169400 24900
rect 169300 24900 169400 25000
rect 169300 25000 169400 25100
rect 169300 25100 169400 25200
rect 169300 25200 169400 25300
rect 169300 25300 169400 25400
rect 169300 25400 169400 25500
rect 169300 25500 169400 25600
rect 169300 25600 169400 25700
rect 169300 25700 169400 25800
rect 169300 25800 169400 25900
rect 169300 25900 169400 26000
rect 169300 26000 169400 26100
rect 169300 26100 169400 26200
rect 169300 26200 169400 26300
rect 169300 26300 169400 26400
rect 169300 26400 169400 26500
rect 169300 26500 169400 26600
rect 169300 26600 169400 26700
rect 169300 26700 169400 26800
rect 169300 26800 169400 26900
rect 169300 26900 169400 27000
rect 169300 27000 169400 27100
rect 169300 27100 169400 27200
rect 169300 27200 169400 27300
rect 169300 27300 169400 27400
rect 169300 27400 169400 27500
rect 169300 27500 169400 27600
rect 169300 27600 169400 27700
rect 169300 27700 169400 27800
rect 169300 27800 169400 27900
rect 169300 27900 169400 28000
rect 169300 28000 169400 28100
rect 169300 28100 169400 28200
rect 169300 28200 169400 28300
rect 169300 28300 169400 28400
rect 169300 28400 169400 28500
rect 169300 28500 169400 28600
rect 169300 28600 169400 28700
rect 169300 28700 169400 28800
rect 169300 28800 169400 28900
rect 169300 28900 169400 29000
rect 169300 29000 169400 29100
rect 169300 29100 169400 29200
rect 169300 29200 169400 29300
rect 169300 29300 169400 29400
rect 169300 29400 169400 29500
rect 169300 29500 169400 29600
rect 169300 29600 169400 29700
rect 169300 29700 169400 29800
rect 169300 29800 169400 29900
rect 169300 29900 169400 30000
rect 169300 30000 169400 30100
rect 169300 30100 169400 30200
rect 169300 30200 169400 30300
rect 169300 30300 169400 30400
rect 169300 30400 169400 30500
rect 169300 30500 169400 30600
rect 169400 24700 169500 24800
rect 169400 24800 169500 24900
rect 169400 24900 169500 25000
rect 169400 25000 169500 25100
rect 169400 25100 169500 25200
rect 169400 25200 169500 25300
rect 169400 25300 169500 25400
rect 169400 25400 169500 25500
rect 169400 25500 169500 25600
rect 169400 25600 169500 25700
rect 169400 25700 169500 25800
rect 169400 25800 169500 25900
rect 169400 25900 169500 26000
rect 169400 26000 169500 26100
rect 169400 26100 169500 26200
rect 169400 26200 169500 26300
rect 169400 26300 169500 26400
rect 169400 26400 169500 26500
rect 169400 26500 169500 26600
rect 169400 26600 169500 26700
rect 169400 26700 169500 26800
rect 169400 26800 169500 26900
rect 169400 26900 169500 27000
rect 169400 27000 169500 27100
rect 169400 27100 169500 27200
rect 169400 27200 169500 27300
rect 169400 27300 169500 27400
rect 169400 27400 169500 27500
rect 169400 27500 169500 27600
rect 169400 27600 169500 27700
rect 169400 27700 169500 27800
rect 169400 27800 169500 27900
rect 169400 27900 169500 28000
rect 169400 28000 169500 28100
rect 169400 28100 169500 28200
rect 169400 28200 169500 28300
rect 169400 28300 169500 28400
rect 169400 28400 169500 28500
rect 169400 28500 169500 28600
rect 169400 28600 169500 28700
rect 169400 28700 169500 28800
rect 169400 28800 169500 28900
rect 169400 28900 169500 29000
rect 169400 29000 169500 29100
rect 169400 29100 169500 29200
rect 169400 29200 169500 29300
rect 169400 29300 169500 29400
rect 169400 29400 169500 29500
rect 169400 29500 169500 29600
rect 169400 29600 169500 29700
rect 169400 29700 169500 29800
rect 169400 29800 169500 29900
rect 169400 29900 169500 30000
rect 169400 30000 169500 30100
rect 169400 30100 169500 30200
rect 169400 30200 169500 30300
rect 169400 30300 169500 30400
rect 169400 30400 169500 30500
rect 169400 30500 169500 30600
rect 169400 30600 169500 30700
rect 169400 30700 169500 30800
rect 169400 30800 169500 30900
rect 169500 25000 169600 25100
rect 169500 25100 169600 25200
rect 169500 25200 169600 25300
rect 169500 25300 169600 25400
rect 169500 25400 169600 25500
rect 169500 25500 169600 25600
rect 169500 25600 169600 25700
rect 169500 25700 169600 25800
rect 169500 25800 169600 25900
rect 169500 25900 169600 26000
rect 169500 26000 169600 26100
rect 169500 26100 169600 26200
rect 169500 26200 169600 26300
rect 169500 26300 169600 26400
rect 169500 26400 169600 26500
rect 169500 26500 169600 26600
rect 169500 26600 169600 26700
rect 169500 26700 169600 26800
rect 169500 26800 169600 26900
rect 169500 26900 169600 27000
rect 169500 27000 169600 27100
rect 169500 27100 169600 27200
rect 169500 27200 169600 27300
rect 169500 27300 169600 27400
rect 169500 27400 169600 27500
rect 169500 27500 169600 27600
rect 169500 27600 169600 27700
rect 169500 27700 169600 27800
rect 169500 27800 169600 27900
rect 169500 27900 169600 28000
rect 169500 28000 169600 28100
rect 169500 28100 169600 28200
rect 169500 28200 169600 28300
rect 169500 28300 169600 28400
rect 169500 28400 169600 28500
rect 169500 28500 169600 28600
rect 169500 28600 169600 28700
rect 169500 28700 169600 28800
rect 169500 28800 169600 28900
rect 169500 28900 169600 29000
rect 169500 29000 169600 29100
rect 169500 29100 169600 29200
rect 169500 29200 169600 29300
rect 169500 29300 169600 29400
rect 169500 29400 169600 29500
rect 169500 29500 169600 29600
rect 169500 29600 169600 29700
rect 169500 29700 169600 29800
rect 169500 29800 169600 29900
rect 169500 29900 169600 30000
rect 169500 30000 169600 30100
rect 169500 30100 169600 30200
rect 169500 30200 169600 30300
rect 169500 30300 169600 30400
rect 169500 30400 169600 30500
rect 169500 30500 169600 30600
rect 169500 30600 169600 30700
rect 169500 30700 169600 30800
rect 169500 30800 169600 30900
rect 169500 30900 169600 31000
rect 169500 31000 169600 31100
rect 169500 31100 169600 31200
rect 169600 25300 169700 25400
rect 169600 25400 169700 25500
rect 169600 25500 169700 25600
rect 169600 25600 169700 25700
rect 169600 25700 169700 25800
rect 169600 25800 169700 25900
rect 169600 25900 169700 26000
rect 169600 26000 169700 26100
rect 169600 26100 169700 26200
rect 169600 26200 169700 26300
rect 169600 26300 169700 26400
rect 169600 26400 169700 26500
rect 169600 26500 169700 26600
rect 169600 26600 169700 26700
rect 169600 26700 169700 26800
rect 169600 26800 169700 26900
rect 169600 26900 169700 27000
rect 169600 27000 169700 27100
rect 169600 27100 169700 27200
rect 169600 27200 169700 27300
rect 169600 27300 169700 27400
rect 169600 27400 169700 27500
rect 169600 27500 169700 27600
rect 169600 27600 169700 27700
rect 169600 27700 169700 27800
rect 169600 27800 169700 27900
rect 169600 27900 169700 28000
rect 169600 28000 169700 28100
rect 169600 28100 169700 28200
rect 169600 28200 169700 28300
rect 169600 28300 169700 28400
rect 169600 28400 169700 28500
rect 169600 28500 169700 28600
rect 169600 28600 169700 28700
rect 169600 28700 169700 28800
rect 169600 28800 169700 28900
rect 169600 28900 169700 29000
rect 169600 29000 169700 29100
rect 169600 29100 169700 29200
rect 169600 29200 169700 29300
rect 169600 29300 169700 29400
rect 169600 29400 169700 29500
rect 169600 29500 169700 29600
rect 169600 29600 169700 29700
rect 169600 29700 169700 29800
rect 169600 29800 169700 29900
rect 169600 29900 169700 30000
rect 169600 30000 169700 30100
rect 169600 30100 169700 30200
rect 169600 30200 169700 30300
rect 169600 30300 169700 30400
rect 169600 30400 169700 30500
rect 169600 30500 169700 30600
rect 169600 30600 169700 30700
rect 169600 30700 169700 30800
rect 169600 30800 169700 30900
rect 169600 30900 169700 31000
rect 169600 31000 169700 31100
rect 169600 31100 169700 31200
rect 169600 31200 169700 31300
rect 169600 31300 169700 31400
rect 169600 31400 169700 31500
rect 169600 31500 169700 31600
rect 169700 25600 169800 25700
rect 169700 25700 169800 25800
rect 169700 25800 169800 25900
rect 169700 25900 169800 26000
rect 169700 26000 169800 26100
rect 169700 26100 169800 26200
rect 169700 26200 169800 26300
rect 169700 26300 169800 26400
rect 169700 26400 169800 26500
rect 169700 26500 169800 26600
rect 169700 26600 169800 26700
rect 169700 26700 169800 26800
rect 169700 26800 169800 26900
rect 169700 26900 169800 27000
rect 169700 27000 169800 27100
rect 169700 27100 169800 27200
rect 169700 27200 169800 27300
rect 169700 27300 169800 27400
rect 169700 27400 169800 27500
rect 169700 27500 169800 27600
rect 169700 27600 169800 27700
rect 169700 27700 169800 27800
rect 169700 27800 169800 27900
rect 169700 27900 169800 28000
rect 169700 28000 169800 28100
rect 169700 28100 169800 28200
rect 169700 28200 169800 28300
rect 169700 28300 169800 28400
rect 169700 28400 169800 28500
rect 169700 28500 169800 28600
rect 169700 28600 169800 28700
rect 169700 28700 169800 28800
rect 169700 28800 169800 28900
rect 169700 28900 169800 29000
rect 169700 29000 169800 29100
rect 169700 29100 169800 29200
rect 169700 29200 169800 29300
rect 169700 29300 169800 29400
rect 169700 29400 169800 29500
rect 169700 29500 169800 29600
rect 169700 29600 169800 29700
rect 169700 29700 169800 29800
rect 169700 29800 169800 29900
rect 169700 29900 169800 30000
rect 169700 30000 169800 30100
rect 169700 30100 169800 30200
rect 169700 30200 169800 30300
rect 169700 30300 169800 30400
rect 169700 30400 169800 30500
rect 169700 30500 169800 30600
rect 169700 30600 169800 30700
rect 169700 30700 169800 30800
rect 169700 30800 169800 30900
rect 169700 30900 169800 31000
rect 169700 31000 169800 31100
rect 169700 31100 169800 31200
rect 169700 31200 169800 31300
rect 169700 31300 169800 31400
rect 169700 31400 169800 31500
rect 169700 31500 169800 31600
rect 169700 31600 169800 31700
rect 169700 31700 169800 31800
rect 169700 31800 169800 31900
rect 169800 25800 169900 25900
rect 169800 25900 169900 26000
rect 169800 26000 169900 26100
rect 169800 26100 169900 26200
rect 169800 26200 169900 26300
rect 169800 26300 169900 26400
rect 169800 26400 169900 26500
rect 169800 26500 169900 26600
rect 169800 26600 169900 26700
rect 169800 26700 169900 26800
rect 169800 26800 169900 26900
rect 169800 26900 169900 27000
rect 169800 27000 169900 27100
rect 169800 27100 169900 27200
rect 169800 27200 169900 27300
rect 169800 27300 169900 27400
rect 169800 27400 169900 27500
rect 169800 27500 169900 27600
rect 169800 27600 169900 27700
rect 169800 27700 169900 27800
rect 169800 27800 169900 27900
rect 169800 27900 169900 28000
rect 169800 28000 169900 28100
rect 169800 28100 169900 28200
rect 169800 28200 169900 28300
rect 169800 28300 169900 28400
rect 169800 28400 169900 28500
rect 169800 28500 169900 28600
rect 169800 28600 169900 28700
rect 169800 28700 169900 28800
rect 169800 28800 169900 28900
rect 169800 28900 169900 29000
rect 169800 29000 169900 29100
rect 169800 29100 169900 29200
rect 169800 29200 169900 29300
rect 169800 29300 169900 29400
rect 169800 29400 169900 29500
rect 169800 29500 169900 29600
rect 169800 29600 169900 29700
rect 169800 29700 169900 29800
rect 169800 29800 169900 29900
rect 169800 29900 169900 30000
rect 169800 30000 169900 30100
rect 169800 30100 169900 30200
rect 169800 30200 169900 30300
rect 169800 30300 169900 30400
rect 169800 30400 169900 30500
rect 169800 30500 169900 30600
rect 169800 30600 169900 30700
rect 169800 30700 169900 30800
rect 169800 30800 169900 30900
rect 169800 30900 169900 31000
rect 169800 31000 169900 31100
rect 169800 31100 169900 31200
rect 169800 31200 169900 31300
rect 169800 31300 169900 31400
rect 169800 31400 169900 31500
rect 169800 31500 169900 31600
rect 169800 31600 169900 31700
rect 169800 31700 169900 31800
rect 169800 31800 169900 31900
rect 169800 31900 169900 32000
rect 169800 32000 169900 32100
rect 169800 32100 169900 32200
rect 169900 26100 170000 26200
rect 169900 26200 170000 26300
rect 169900 26300 170000 26400
rect 169900 26400 170000 26500
rect 169900 26500 170000 26600
rect 169900 26600 170000 26700
rect 169900 26700 170000 26800
rect 169900 26800 170000 26900
rect 169900 26900 170000 27000
rect 169900 27000 170000 27100
rect 169900 27100 170000 27200
rect 169900 27200 170000 27300
rect 169900 27300 170000 27400
rect 169900 27400 170000 27500
rect 169900 27500 170000 27600
rect 169900 27600 170000 27700
rect 169900 27700 170000 27800
rect 169900 27800 170000 27900
rect 169900 27900 170000 28000
rect 169900 28000 170000 28100
rect 169900 28100 170000 28200
rect 169900 28200 170000 28300
rect 169900 28300 170000 28400
rect 169900 28400 170000 28500
rect 169900 28500 170000 28600
rect 169900 28600 170000 28700
rect 169900 28700 170000 28800
rect 169900 28800 170000 28900
rect 169900 28900 170000 29000
rect 169900 29000 170000 29100
rect 169900 29100 170000 29200
rect 169900 29200 170000 29300
rect 169900 29300 170000 29400
rect 169900 29400 170000 29500
rect 169900 29500 170000 29600
rect 169900 29600 170000 29700
rect 169900 29700 170000 29800
rect 169900 29800 170000 29900
rect 169900 29900 170000 30000
rect 169900 30000 170000 30100
rect 169900 30100 170000 30200
rect 169900 30200 170000 30300
rect 169900 30300 170000 30400
rect 169900 30400 170000 30500
rect 169900 30500 170000 30600
rect 169900 30600 170000 30700
rect 169900 30700 170000 30800
rect 169900 30800 170000 30900
rect 169900 30900 170000 31000
rect 169900 31000 170000 31100
rect 169900 31100 170000 31200
rect 169900 31200 170000 31300
rect 169900 31300 170000 31400
rect 169900 31400 170000 31500
rect 169900 31500 170000 31600
rect 169900 31600 170000 31700
rect 169900 31700 170000 31800
rect 169900 31800 170000 31900
rect 169900 31900 170000 32000
rect 169900 32000 170000 32100
rect 169900 32100 170000 32200
rect 169900 32200 170000 32300
rect 169900 32300 170000 32400
rect 169900 32400 170000 32500
rect 170000 26300 170100 26400
rect 170000 26400 170100 26500
rect 170000 26500 170100 26600
rect 170000 26600 170100 26700
rect 170000 26700 170100 26800
rect 170000 26800 170100 26900
rect 170000 26900 170100 27000
rect 170000 27000 170100 27100
rect 170000 27100 170100 27200
rect 170000 27200 170100 27300
rect 170000 27300 170100 27400
rect 170000 27400 170100 27500
rect 170000 27500 170100 27600
rect 170000 27600 170100 27700
rect 170000 27700 170100 27800
rect 170000 27800 170100 27900
rect 170000 27900 170100 28000
rect 170000 28000 170100 28100
rect 170000 28100 170100 28200
rect 170000 28200 170100 28300
rect 170000 28300 170100 28400
rect 170000 28400 170100 28500
rect 170000 28500 170100 28600
rect 170000 28600 170100 28700
rect 170000 28700 170100 28800
rect 170000 28800 170100 28900
rect 170000 28900 170100 29000
rect 170000 29000 170100 29100
rect 170000 29100 170100 29200
rect 170000 29200 170100 29300
rect 170000 29300 170100 29400
rect 170000 29400 170100 29500
rect 170000 29500 170100 29600
rect 170000 29600 170100 29700
rect 170000 29700 170100 29800
rect 170000 29800 170100 29900
rect 170000 29900 170100 30000
rect 170000 30000 170100 30100
rect 170000 30100 170100 30200
rect 170000 30200 170100 30300
rect 170000 30300 170100 30400
rect 170000 30400 170100 30500
rect 170000 30500 170100 30600
rect 170000 30600 170100 30700
rect 170000 30700 170100 30800
rect 170000 30800 170100 30900
rect 170000 30900 170100 31000
rect 170000 31000 170100 31100
rect 170000 31100 170100 31200
rect 170000 31200 170100 31300
rect 170000 31300 170100 31400
rect 170000 31400 170100 31500
rect 170000 31500 170100 31600
rect 170000 31600 170100 31700
rect 170000 31700 170100 31800
rect 170000 31800 170100 31900
rect 170000 31900 170100 32000
rect 170000 32000 170100 32100
rect 170000 32100 170100 32200
rect 170000 32200 170100 32300
rect 170000 32300 170100 32400
rect 170000 32400 170100 32500
rect 170000 32500 170100 32600
rect 170000 32600 170100 32700
rect 170000 32700 170100 32800
rect 170100 26500 170200 26600
rect 170100 26600 170200 26700
rect 170100 26700 170200 26800
rect 170100 26800 170200 26900
rect 170100 26900 170200 27000
rect 170100 27000 170200 27100
rect 170100 27100 170200 27200
rect 170100 27200 170200 27300
rect 170100 27300 170200 27400
rect 170100 27400 170200 27500
rect 170100 27500 170200 27600
rect 170100 27600 170200 27700
rect 170100 27700 170200 27800
rect 170100 27800 170200 27900
rect 170100 27900 170200 28000
rect 170100 28000 170200 28100
rect 170100 28100 170200 28200
rect 170100 28200 170200 28300
rect 170100 28300 170200 28400
rect 170100 28400 170200 28500
rect 170100 28500 170200 28600
rect 170100 28600 170200 28700
rect 170100 28700 170200 28800
rect 170100 28800 170200 28900
rect 170100 28900 170200 29000
rect 170100 29000 170200 29100
rect 170100 29100 170200 29200
rect 170100 29200 170200 29300
rect 170100 29300 170200 29400
rect 170100 29400 170200 29500
rect 170100 29500 170200 29600
rect 170100 29600 170200 29700
rect 170100 29700 170200 29800
rect 170100 29800 170200 29900
rect 170100 29900 170200 30000
rect 170100 30000 170200 30100
rect 170100 30100 170200 30200
rect 170100 30200 170200 30300
rect 170100 30300 170200 30400
rect 170100 30400 170200 30500
rect 170100 30500 170200 30600
rect 170100 30600 170200 30700
rect 170100 30700 170200 30800
rect 170100 30800 170200 30900
rect 170100 30900 170200 31000
rect 170100 31000 170200 31100
rect 170100 31100 170200 31200
rect 170100 31200 170200 31300
rect 170100 31300 170200 31400
rect 170100 31400 170200 31500
rect 170100 31500 170200 31600
rect 170100 31600 170200 31700
rect 170100 31700 170200 31800
rect 170100 31800 170200 31900
rect 170100 31900 170200 32000
rect 170100 32000 170200 32100
rect 170100 32100 170200 32200
rect 170100 32200 170200 32300
rect 170100 32300 170200 32400
rect 170100 32400 170200 32500
rect 170100 32500 170200 32600
rect 170100 32600 170200 32700
rect 170100 32700 170200 32800
rect 170100 32800 170200 32900
rect 170100 32900 170200 33000
rect 170100 33000 170200 33100
rect 170100 33100 170200 33200
rect 170200 26800 170300 26900
rect 170200 26900 170300 27000
rect 170200 27000 170300 27100
rect 170200 27100 170300 27200
rect 170200 27200 170300 27300
rect 170200 27300 170300 27400
rect 170200 27400 170300 27500
rect 170200 27500 170300 27600
rect 170200 27600 170300 27700
rect 170200 27700 170300 27800
rect 170200 27800 170300 27900
rect 170200 27900 170300 28000
rect 170200 28000 170300 28100
rect 170200 28100 170300 28200
rect 170200 28200 170300 28300
rect 170200 28300 170300 28400
rect 170200 28400 170300 28500
rect 170200 28500 170300 28600
rect 170200 28600 170300 28700
rect 170200 28700 170300 28800
rect 170200 28800 170300 28900
rect 170200 28900 170300 29000
rect 170200 29000 170300 29100
rect 170200 29100 170300 29200
rect 170200 29200 170300 29300
rect 170200 29300 170300 29400
rect 170200 29400 170300 29500
rect 170200 29500 170300 29600
rect 170200 29600 170300 29700
rect 170200 29700 170300 29800
rect 170200 29800 170300 29900
rect 170200 29900 170300 30000
rect 170200 30000 170300 30100
rect 170200 30100 170300 30200
rect 170200 30200 170300 30300
rect 170200 30300 170300 30400
rect 170200 30400 170300 30500
rect 170200 30500 170300 30600
rect 170200 30600 170300 30700
rect 170200 30700 170300 30800
rect 170200 30800 170300 30900
rect 170200 30900 170300 31000
rect 170200 31000 170300 31100
rect 170200 31100 170300 31200
rect 170200 31200 170300 31300
rect 170200 31300 170300 31400
rect 170200 31400 170300 31500
rect 170200 31500 170300 31600
rect 170200 31600 170300 31700
rect 170200 31700 170300 31800
rect 170200 31800 170300 31900
rect 170200 31900 170300 32000
rect 170200 32000 170300 32100
rect 170200 32100 170300 32200
rect 170200 32200 170300 32300
rect 170200 32300 170300 32400
rect 170200 32400 170300 32500
rect 170200 32500 170300 32600
rect 170200 32600 170300 32700
rect 170200 32700 170300 32800
rect 170200 32800 170300 32900
rect 170200 32900 170300 33000
rect 170200 33000 170300 33100
rect 170200 33100 170300 33200
rect 170200 33200 170300 33300
rect 170200 33300 170300 33400
rect 170200 33400 170300 33500
rect 170300 27000 170400 27100
rect 170300 27100 170400 27200
rect 170300 27200 170400 27300
rect 170300 27300 170400 27400
rect 170300 27400 170400 27500
rect 170300 27500 170400 27600
rect 170300 27600 170400 27700
rect 170300 27700 170400 27800
rect 170300 27800 170400 27900
rect 170300 27900 170400 28000
rect 170300 28000 170400 28100
rect 170300 28100 170400 28200
rect 170300 28200 170400 28300
rect 170300 28300 170400 28400
rect 170300 28400 170400 28500
rect 170300 28500 170400 28600
rect 170300 28600 170400 28700
rect 170300 28700 170400 28800
rect 170300 28800 170400 28900
rect 170300 28900 170400 29000
rect 170300 29000 170400 29100
rect 170300 29100 170400 29200
rect 170300 29200 170400 29300
rect 170300 29300 170400 29400
rect 170300 29400 170400 29500
rect 170300 29500 170400 29600
rect 170300 29600 170400 29700
rect 170300 29700 170400 29800
rect 170300 29800 170400 29900
rect 170300 29900 170400 30000
rect 170300 30000 170400 30100
rect 170300 30100 170400 30200
rect 170300 30200 170400 30300
rect 170300 30300 170400 30400
rect 170300 30400 170400 30500
rect 170300 30500 170400 30600
rect 170300 30600 170400 30700
rect 170300 30700 170400 30800
rect 170300 30800 170400 30900
rect 170300 30900 170400 31000
rect 170300 31000 170400 31100
rect 170300 31100 170400 31200
rect 170300 31200 170400 31300
rect 170300 31300 170400 31400
rect 170300 31400 170400 31500
rect 170300 31500 170400 31600
rect 170300 31600 170400 31700
rect 170300 31700 170400 31800
rect 170300 31800 170400 31900
rect 170300 31900 170400 32000
rect 170300 32000 170400 32100
rect 170300 32100 170400 32200
rect 170300 32200 170400 32300
rect 170300 32300 170400 32400
rect 170300 32400 170400 32500
rect 170300 32500 170400 32600
rect 170300 32600 170400 32700
rect 170300 32700 170400 32800
rect 170300 32800 170400 32900
rect 170300 32900 170400 33000
rect 170300 33000 170400 33100
rect 170300 33100 170400 33200
rect 170300 33200 170400 33300
rect 170300 33300 170400 33400
rect 170300 33400 170400 33500
rect 170300 33500 170400 33600
rect 170300 33600 170400 33700
rect 170300 33700 170400 33800
rect 170400 27200 170500 27300
rect 170400 27300 170500 27400
rect 170400 27400 170500 27500
rect 170400 27500 170500 27600
rect 170400 27600 170500 27700
rect 170400 27700 170500 27800
rect 170400 27800 170500 27900
rect 170400 27900 170500 28000
rect 170400 28000 170500 28100
rect 170400 28100 170500 28200
rect 170400 28200 170500 28300
rect 170400 28300 170500 28400
rect 170400 28400 170500 28500
rect 170400 28500 170500 28600
rect 170400 28600 170500 28700
rect 170400 28700 170500 28800
rect 170400 28800 170500 28900
rect 170400 28900 170500 29000
rect 170400 29000 170500 29100
rect 170400 29100 170500 29200
rect 170400 29200 170500 29300
rect 170400 29300 170500 29400
rect 170400 29400 170500 29500
rect 170400 29500 170500 29600
rect 170400 29600 170500 29700
rect 170400 29700 170500 29800
rect 170400 29800 170500 29900
rect 170400 29900 170500 30000
rect 170400 30000 170500 30100
rect 170400 30100 170500 30200
rect 170400 30200 170500 30300
rect 170400 30300 170500 30400
rect 170400 30400 170500 30500
rect 170400 30500 170500 30600
rect 170400 30600 170500 30700
rect 170400 30700 170500 30800
rect 170400 30800 170500 30900
rect 170400 30900 170500 31000
rect 170400 31000 170500 31100
rect 170400 31100 170500 31200
rect 170400 31200 170500 31300
rect 170400 31300 170500 31400
rect 170400 31400 170500 31500
rect 170400 31500 170500 31600
rect 170400 31600 170500 31700
rect 170400 31700 170500 31800
rect 170400 31800 170500 31900
rect 170400 31900 170500 32000
rect 170400 32000 170500 32100
rect 170400 32100 170500 32200
rect 170400 32200 170500 32300
rect 170400 32300 170500 32400
rect 170400 32400 170500 32500
rect 170400 32500 170500 32600
rect 170400 32600 170500 32700
rect 170400 32700 170500 32800
rect 170400 32800 170500 32900
rect 170400 32900 170500 33000
rect 170400 33000 170500 33100
rect 170400 33100 170500 33200
rect 170400 33200 170500 33300
rect 170400 33300 170500 33400
rect 170400 33400 170500 33500
rect 170400 33500 170500 33600
rect 170400 33600 170500 33700
rect 170400 33700 170500 33800
rect 170400 33800 170500 33900
rect 170400 33900 170500 34000
rect 170400 34000 170500 34100
rect 170500 27500 170600 27600
rect 170500 27600 170600 27700
rect 170500 27700 170600 27800
rect 170500 27800 170600 27900
rect 170500 27900 170600 28000
rect 170500 28000 170600 28100
rect 170500 28100 170600 28200
rect 170500 28200 170600 28300
rect 170500 28300 170600 28400
rect 170500 28400 170600 28500
rect 170500 28500 170600 28600
rect 170500 28600 170600 28700
rect 170500 28700 170600 28800
rect 170500 28800 170600 28900
rect 170500 28900 170600 29000
rect 170500 29000 170600 29100
rect 170500 29100 170600 29200
rect 170500 29200 170600 29300
rect 170500 29300 170600 29400
rect 170500 29400 170600 29500
rect 170500 29500 170600 29600
rect 170500 29600 170600 29700
rect 170500 29700 170600 29800
rect 170500 29800 170600 29900
rect 170500 29900 170600 30000
rect 170500 30000 170600 30100
rect 170500 30100 170600 30200
rect 170500 30200 170600 30300
rect 170500 30300 170600 30400
rect 170500 30400 170600 30500
rect 170500 30500 170600 30600
rect 170500 30600 170600 30700
rect 170500 30700 170600 30800
rect 170500 30800 170600 30900
rect 170500 30900 170600 31000
rect 170500 31000 170600 31100
rect 170500 31100 170600 31200
rect 170500 31200 170600 31300
rect 170500 31300 170600 31400
rect 170500 31400 170600 31500
rect 170500 31500 170600 31600
rect 170500 31600 170600 31700
rect 170500 31700 170600 31800
rect 170500 31800 170600 31900
rect 170500 31900 170600 32000
rect 170500 32000 170600 32100
rect 170500 32100 170600 32200
rect 170500 32200 170600 32300
rect 170500 32300 170600 32400
rect 170500 32400 170600 32500
rect 170500 32500 170600 32600
rect 170500 32600 170600 32700
rect 170500 32700 170600 32800
rect 170500 32800 170600 32900
rect 170500 32900 170600 33000
rect 170500 33000 170600 33100
rect 170500 33100 170600 33200
rect 170500 33200 170600 33300
rect 170500 33300 170600 33400
rect 170500 33400 170600 33500
rect 170500 33500 170600 33600
rect 170500 33600 170600 33700
rect 170500 33700 170600 33800
rect 170500 33800 170600 33900
rect 170500 33900 170600 34000
rect 170500 34000 170600 34100
rect 170500 34100 170600 34200
rect 170500 34200 170600 34300
rect 170500 34300 170600 34400
rect 170600 27700 170700 27800
rect 170600 27800 170700 27900
rect 170600 27900 170700 28000
rect 170600 28000 170700 28100
rect 170600 28100 170700 28200
rect 170600 28200 170700 28300
rect 170600 28300 170700 28400
rect 170600 28400 170700 28500
rect 170600 28500 170700 28600
rect 170600 28600 170700 28700
rect 170600 28700 170700 28800
rect 170600 28800 170700 28900
rect 170600 28900 170700 29000
rect 170600 29000 170700 29100
rect 170600 29100 170700 29200
rect 170600 29200 170700 29300
rect 170600 29300 170700 29400
rect 170600 29400 170700 29500
rect 170600 29500 170700 29600
rect 170600 29600 170700 29700
rect 170600 29700 170700 29800
rect 170600 29800 170700 29900
rect 170600 29900 170700 30000
rect 170600 30000 170700 30100
rect 170600 30100 170700 30200
rect 170600 30200 170700 30300
rect 170600 30300 170700 30400
rect 170600 30400 170700 30500
rect 170600 30500 170700 30600
rect 170600 30600 170700 30700
rect 170600 30700 170700 30800
rect 170600 30800 170700 30900
rect 170600 30900 170700 31000
rect 170600 31000 170700 31100
rect 170600 31100 170700 31200
rect 170600 31200 170700 31300
rect 170600 31300 170700 31400
rect 170600 31400 170700 31500
rect 170600 31500 170700 31600
rect 170600 31600 170700 31700
rect 170600 31700 170700 31800
rect 170600 31800 170700 31900
rect 170600 31900 170700 32000
rect 170600 32000 170700 32100
rect 170600 32100 170700 32200
rect 170600 32200 170700 32300
rect 170600 32300 170700 32400
rect 170600 32400 170700 32500
rect 170600 32500 170700 32600
rect 170600 32600 170700 32700
rect 170600 32700 170700 32800
rect 170600 32800 170700 32900
rect 170600 32900 170700 33000
rect 170600 33000 170700 33100
rect 170600 33100 170700 33200
rect 170600 33200 170700 33300
rect 170600 33300 170700 33400
rect 170600 33400 170700 33500
rect 170600 33500 170700 33600
rect 170600 33600 170700 33700
rect 170600 33700 170700 33800
rect 170600 33800 170700 33900
rect 170600 33900 170700 34000
rect 170600 34000 170700 34100
rect 170600 34100 170700 34200
rect 170600 34200 170700 34300
rect 170600 34300 170700 34400
rect 170600 34400 170700 34500
rect 170600 34500 170700 34600
rect 170600 34600 170700 34700
rect 170700 27900 170800 28000
rect 170700 28000 170800 28100
rect 170700 28100 170800 28200
rect 170700 28200 170800 28300
rect 170700 28300 170800 28400
rect 170700 28400 170800 28500
rect 170700 28500 170800 28600
rect 170700 28600 170800 28700
rect 170700 28700 170800 28800
rect 170700 28800 170800 28900
rect 170700 28900 170800 29000
rect 170700 29000 170800 29100
rect 170700 29100 170800 29200
rect 170700 29200 170800 29300
rect 170700 29300 170800 29400
rect 170700 29400 170800 29500
rect 170700 29500 170800 29600
rect 170700 29600 170800 29700
rect 170700 29700 170800 29800
rect 170700 29800 170800 29900
rect 170700 29900 170800 30000
rect 170700 30000 170800 30100
rect 170700 30100 170800 30200
rect 170700 30200 170800 30300
rect 170700 30300 170800 30400
rect 170700 30400 170800 30500
rect 170700 30500 170800 30600
rect 170700 30600 170800 30700
rect 170700 30700 170800 30800
rect 170700 30800 170800 30900
rect 170700 30900 170800 31000
rect 170700 31000 170800 31100
rect 170700 31100 170800 31200
rect 170700 31200 170800 31300
rect 170700 31300 170800 31400
rect 170700 31400 170800 31500
rect 170700 31500 170800 31600
rect 170700 31600 170800 31700
rect 170700 31700 170800 31800
rect 170700 31800 170800 31900
rect 170700 31900 170800 32000
rect 170700 32000 170800 32100
rect 170700 32100 170800 32200
rect 170700 32200 170800 32300
rect 170700 32300 170800 32400
rect 170700 32400 170800 32500
rect 170700 32500 170800 32600
rect 170700 32600 170800 32700
rect 170700 32700 170800 32800
rect 170700 32800 170800 32900
rect 170700 32900 170800 33000
rect 170700 33000 170800 33100
rect 170700 33100 170800 33200
rect 170700 33200 170800 33300
rect 170700 33300 170800 33400
rect 170700 33400 170800 33500
rect 170700 33500 170800 33600
rect 170700 33600 170800 33700
rect 170700 33700 170800 33800
rect 170700 33800 170800 33900
rect 170700 33900 170800 34000
rect 170700 34000 170800 34100
rect 170700 34100 170800 34200
rect 170700 34200 170800 34300
rect 170700 34300 170800 34400
rect 170700 34400 170800 34500
rect 170700 34500 170800 34600
rect 170700 34600 170800 34700
rect 170700 34700 170800 34800
rect 170700 34800 170800 34900
rect 170700 34900 170800 35000
rect 170800 28200 170900 28300
rect 170800 28300 170900 28400
rect 170800 28400 170900 28500
rect 170800 28500 170900 28600
rect 170800 28600 170900 28700
rect 170800 28700 170900 28800
rect 170800 28800 170900 28900
rect 170800 28900 170900 29000
rect 170800 29000 170900 29100
rect 170800 29100 170900 29200
rect 170800 29200 170900 29300
rect 170800 29300 170900 29400
rect 170800 29400 170900 29500
rect 170800 29500 170900 29600
rect 170800 29600 170900 29700
rect 170800 29700 170900 29800
rect 170800 29800 170900 29900
rect 170800 29900 170900 30000
rect 170800 30000 170900 30100
rect 170800 30100 170900 30200
rect 170800 30200 170900 30300
rect 170800 30300 170900 30400
rect 170800 30400 170900 30500
rect 170800 30500 170900 30600
rect 170800 30600 170900 30700
rect 170800 30700 170900 30800
rect 170800 30800 170900 30900
rect 170800 30900 170900 31000
rect 170800 31000 170900 31100
rect 170800 31100 170900 31200
rect 170800 31200 170900 31300
rect 170800 31300 170900 31400
rect 170800 31400 170900 31500
rect 170800 31500 170900 31600
rect 170800 31600 170900 31700
rect 170800 31700 170900 31800
rect 170800 31800 170900 31900
rect 170800 31900 170900 32000
rect 170800 32000 170900 32100
rect 170800 32100 170900 32200
rect 170800 32200 170900 32300
rect 170800 32300 170900 32400
rect 170800 32400 170900 32500
rect 170800 32500 170900 32600
rect 170800 32600 170900 32700
rect 170800 32700 170900 32800
rect 170800 32800 170900 32900
rect 170800 32900 170900 33000
rect 170800 33000 170900 33100
rect 170800 33100 170900 33200
rect 170800 33200 170900 33300
rect 170800 33300 170900 33400
rect 170800 33400 170900 33500
rect 170800 33500 170900 33600
rect 170800 33600 170900 33700
rect 170800 33700 170900 33800
rect 170800 33800 170900 33900
rect 170800 33900 170900 34000
rect 170800 34000 170900 34100
rect 170800 34100 170900 34200
rect 170800 34200 170900 34300
rect 170800 34300 170900 34400
rect 170800 34400 170900 34500
rect 170800 34500 170900 34600
rect 170800 34600 170900 34700
rect 170800 34700 170900 34800
rect 170800 34800 170900 34900
rect 170800 34900 170900 35000
rect 170800 35000 170900 35100
rect 170800 35100 170900 35200
rect 170800 35200 170900 35300
rect 170900 28400 171000 28500
rect 170900 28500 171000 28600
rect 170900 28600 171000 28700
rect 170900 28700 171000 28800
rect 170900 28800 171000 28900
rect 170900 28900 171000 29000
rect 170900 29000 171000 29100
rect 170900 29100 171000 29200
rect 170900 29200 171000 29300
rect 170900 29300 171000 29400
rect 170900 29400 171000 29500
rect 170900 29500 171000 29600
rect 170900 29600 171000 29700
rect 170900 29700 171000 29800
rect 170900 29800 171000 29900
rect 170900 29900 171000 30000
rect 170900 30000 171000 30100
rect 170900 30100 171000 30200
rect 170900 30200 171000 30300
rect 170900 30300 171000 30400
rect 170900 30400 171000 30500
rect 170900 30500 171000 30600
rect 170900 30600 171000 30700
rect 170900 30700 171000 30800
rect 170900 30800 171000 30900
rect 170900 30900 171000 31000
rect 170900 31000 171000 31100
rect 170900 31100 171000 31200
rect 170900 31200 171000 31300
rect 170900 31300 171000 31400
rect 170900 31400 171000 31500
rect 170900 31500 171000 31600
rect 170900 31600 171000 31700
rect 170900 31700 171000 31800
rect 170900 31800 171000 31900
rect 170900 31900 171000 32000
rect 170900 32000 171000 32100
rect 170900 32100 171000 32200
rect 170900 32200 171000 32300
rect 170900 32300 171000 32400
rect 170900 32400 171000 32500
rect 170900 32500 171000 32600
rect 170900 32600 171000 32700
rect 170900 32700 171000 32800
rect 170900 32800 171000 32900
rect 170900 32900 171000 33000
rect 170900 33000 171000 33100
rect 170900 33100 171000 33200
rect 170900 33200 171000 33300
rect 170900 33300 171000 33400
rect 170900 33400 171000 33500
rect 170900 33500 171000 33600
rect 170900 33600 171000 33700
rect 170900 33700 171000 33800
rect 170900 33800 171000 33900
rect 170900 33900 171000 34000
rect 170900 34000 171000 34100
rect 170900 34100 171000 34200
rect 170900 34200 171000 34300
rect 170900 34300 171000 34400
rect 170900 34400 171000 34500
rect 170900 34500 171000 34600
rect 170900 34600 171000 34700
rect 170900 34700 171000 34800
rect 170900 34800 171000 34900
rect 170900 34900 171000 35000
rect 170900 35000 171000 35100
rect 170900 35100 171000 35200
rect 170900 35200 171000 35300
rect 170900 35300 171000 35400
rect 170900 35400 171000 35500
rect 170900 35500 171000 35600
rect 171000 28700 171100 28800
rect 171000 28800 171100 28900
rect 171000 28900 171100 29000
rect 171000 29000 171100 29100
rect 171000 29100 171100 29200
rect 171000 29200 171100 29300
rect 171000 29300 171100 29400
rect 171000 29400 171100 29500
rect 171000 29500 171100 29600
rect 171000 29600 171100 29700
rect 171000 29700 171100 29800
rect 171000 29800 171100 29900
rect 171000 29900 171100 30000
rect 171000 30000 171100 30100
rect 171000 30100 171100 30200
rect 171000 30200 171100 30300
rect 171000 30300 171100 30400
rect 171000 30400 171100 30500
rect 171000 30500 171100 30600
rect 171000 30600 171100 30700
rect 171000 30700 171100 30800
rect 171000 30800 171100 30900
rect 171000 30900 171100 31000
rect 171000 31000 171100 31100
rect 171000 31100 171100 31200
rect 171000 31200 171100 31300
rect 171000 31300 171100 31400
rect 171000 31400 171100 31500
rect 171000 31500 171100 31600
rect 171000 31600 171100 31700
rect 171000 31700 171100 31800
rect 171000 31800 171100 31900
rect 171000 31900 171100 32000
rect 171000 32000 171100 32100
rect 171000 32100 171100 32200
rect 171000 32200 171100 32300
rect 171000 32300 171100 32400
rect 171000 32400 171100 32500
rect 171000 32500 171100 32600
rect 171000 32600 171100 32700
rect 171000 32700 171100 32800
rect 171000 32800 171100 32900
rect 171000 32900 171100 33000
rect 171000 33000 171100 33100
rect 171000 33100 171100 33200
rect 171000 33200 171100 33300
rect 171000 33300 171100 33400
rect 171000 33400 171100 33500
rect 171000 33500 171100 33600
rect 171000 33600 171100 33700
rect 171000 33700 171100 33800
rect 171000 33800 171100 33900
rect 171000 33900 171100 34000
rect 171000 34000 171100 34100
rect 171000 34100 171100 34200
rect 171000 34200 171100 34300
rect 171000 34300 171100 34400
rect 171000 34400 171100 34500
rect 171000 34500 171100 34600
rect 171000 34600 171100 34700
rect 171000 34700 171100 34800
rect 171000 34800 171100 34900
rect 171000 34900 171100 35000
rect 171000 35000 171100 35100
rect 171000 35100 171100 35200
rect 171000 35200 171100 35300
rect 171000 35300 171100 35400
rect 171000 35400 171100 35500
rect 171000 35500 171100 35600
rect 171000 35600 171100 35700
rect 171000 35700 171100 35800
rect 171100 28900 171200 29000
rect 171100 29000 171200 29100
rect 171100 29100 171200 29200
rect 171100 29200 171200 29300
rect 171100 29300 171200 29400
rect 171100 29400 171200 29500
rect 171100 29500 171200 29600
rect 171100 29600 171200 29700
rect 171100 29700 171200 29800
rect 171100 29800 171200 29900
rect 171100 29900 171200 30000
rect 171100 30000 171200 30100
rect 171100 30100 171200 30200
rect 171100 30200 171200 30300
rect 171100 30300 171200 30400
rect 171100 30400 171200 30500
rect 171100 30500 171200 30600
rect 171100 30600 171200 30700
rect 171100 30700 171200 30800
rect 171100 30800 171200 30900
rect 171100 30900 171200 31000
rect 171100 31000 171200 31100
rect 171100 31100 171200 31200
rect 171100 31200 171200 31300
rect 171100 31300 171200 31400
rect 171100 31400 171200 31500
rect 171100 31500 171200 31600
rect 171100 31600 171200 31700
rect 171100 31700 171200 31800
rect 171100 31800 171200 31900
rect 171100 31900 171200 32000
rect 171100 32000 171200 32100
rect 171100 32100 171200 32200
rect 171100 32200 171200 32300
rect 171100 32300 171200 32400
rect 171100 32400 171200 32500
rect 171100 32500 171200 32600
rect 171100 32600 171200 32700
rect 171100 32700 171200 32800
rect 171100 32800 171200 32900
rect 171100 32900 171200 33000
rect 171100 33000 171200 33100
rect 171100 33100 171200 33200
rect 171100 33200 171200 33300
rect 171100 33300 171200 33400
rect 171100 33400 171200 33500
rect 171100 33500 171200 33600
rect 171100 33600 171200 33700
rect 171100 33700 171200 33800
rect 171100 33800 171200 33900
rect 171100 33900 171200 34000
rect 171100 34000 171200 34100
rect 171100 34100 171200 34200
rect 171100 34200 171200 34300
rect 171100 34300 171200 34400
rect 171100 34400 171200 34500
rect 171100 34500 171200 34600
rect 171100 34600 171200 34700
rect 171100 34700 171200 34800
rect 171100 34800 171200 34900
rect 171100 34900 171200 35000
rect 171100 35000 171200 35100
rect 171100 35100 171200 35200
rect 171100 35200 171200 35300
rect 171100 35300 171200 35400
rect 171100 35400 171200 35500
rect 171100 35500 171200 35600
rect 171100 35600 171200 35700
rect 171100 35700 171200 35800
rect 171100 35800 171200 35900
rect 171100 35900 171200 36000
rect 171200 29200 171300 29300
rect 171200 29300 171300 29400
rect 171200 29400 171300 29500
rect 171200 29500 171300 29600
rect 171200 29600 171300 29700
rect 171200 29700 171300 29800
rect 171200 29800 171300 29900
rect 171200 29900 171300 30000
rect 171200 30000 171300 30100
rect 171200 30100 171300 30200
rect 171200 30200 171300 30300
rect 171200 30300 171300 30400
rect 171200 30400 171300 30500
rect 171200 30500 171300 30600
rect 171200 30600 171300 30700
rect 171200 30700 171300 30800
rect 171200 30800 171300 30900
rect 171200 30900 171300 31000
rect 171200 31000 171300 31100
rect 171200 31100 171300 31200
rect 171200 31200 171300 31300
rect 171200 31300 171300 31400
rect 171200 31400 171300 31500
rect 171200 31500 171300 31600
rect 171200 31600 171300 31700
rect 171200 31700 171300 31800
rect 171200 31800 171300 31900
rect 171200 31900 171300 32000
rect 171200 32000 171300 32100
rect 171200 32100 171300 32200
rect 171200 32200 171300 32300
rect 171200 32300 171300 32400
rect 171200 32400 171300 32500
rect 171200 32500 171300 32600
rect 171200 32600 171300 32700
rect 171200 32700 171300 32800
rect 171200 32800 171300 32900
rect 171200 32900 171300 33000
rect 171200 33000 171300 33100
rect 171200 33100 171300 33200
rect 171200 33200 171300 33300
rect 171200 33300 171300 33400
rect 171200 33400 171300 33500
rect 171200 33500 171300 33600
rect 171200 33600 171300 33700
rect 171200 33700 171300 33800
rect 171200 33800 171300 33900
rect 171200 33900 171300 34000
rect 171200 34000 171300 34100
rect 171200 34100 171300 34200
rect 171200 34200 171300 34300
rect 171200 34300 171300 34400
rect 171200 34400 171300 34500
rect 171200 34500 171300 34600
rect 171200 34600 171300 34700
rect 171200 34700 171300 34800
rect 171200 34800 171300 34900
rect 171200 34900 171300 35000
rect 171200 35000 171300 35100
rect 171200 35100 171300 35200
rect 171200 35200 171300 35300
rect 171200 35300 171300 35400
rect 171200 35400 171300 35500
rect 171200 35500 171300 35600
rect 171200 35600 171300 35700
rect 171200 35700 171300 35800
rect 171200 35800 171300 35900
rect 171200 35900 171300 36000
rect 171200 36000 171300 36100
rect 171200 36100 171300 36200
rect 171200 36200 171300 36300
rect 171300 29500 171400 29600
rect 171300 29600 171400 29700
rect 171300 29700 171400 29800
rect 171300 29800 171400 29900
rect 171300 29900 171400 30000
rect 171300 30000 171400 30100
rect 171300 30100 171400 30200
rect 171300 30200 171400 30300
rect 171300 30300 171400 30400
rect 171300 30400 171400 30500
rect 171300 30500 171400 30600
rect 171300 30600 171400 30700
rect 171300 30700 171400 30800
rect 171300 30800 171400 30900
rect 171300 30900 171400 31000
rect 171300 31000 171400 31100
rect 171300 31100 171400 31200
rect 171300 31200 171400 31300
rect 171300 31300 171400 31400
rect 171300 31400 171400 31500
rect 171300 31500 171400 31600
rect 171300 31600 171400 31700
rect 171300 31700 171400 31800
rect 171300 31800 171400 31900
rect 171300 31900 171400 32000
rect 171300 32000 171400 32100
rect 171300 32100 171400 32200
rect 171300 32200 171400 32300
rect 171300 32300 171400 32400
rect 171300 32400 171400 32500
rect 171300 32500 171400 32600
rect 171300 32600 171400 32700
rect 171300 32700 171400 32800
rect 171300 32800 171400 32900
rect 171300 32900 171400 33000
rect 171300 33000 171400 33100
rect 171300 33100 171400 33200
rect 171300 33200 171400 33300
rect 171300 33300 171400 33400
rect 171300 33400 171400 33500
rect 171300 33500 171400 33600
rect 171300 33600 171400 33700
rect 171300 33700 171400 33800
rect 171300 33800 171400 33900
rect 171300 33900 171400 34000
rect 171300 34000 171400 34100
rect 171300 34100 171400 34200
rect 171300 34200 171400 34300
rect 171300 34300 171400 34400
rect 171300 34400 171400 34500
rect 171300 34500 171400 34600
rect 171300 34600 171400 34700
rect 171300 34700 171400 34800
rect 171300 34800 171400 34900
rect 171300 34900 171400 35000
rect 171300 35000 171400 35100
rect 171300 35100 171400 35200
rect 171300 35200 171400 35300
rect 171300 35300 171400 35400
rect 171300 35400 171400 35500
rect 171300 35500 171400 35600
rect 171300 35600 171400 35700
rect 171300 35700 171400 35800
rect 171300 35800 171400 35900
rect 171300 35900 171400 36000
rect 171300 36000 171400 36100
rect 171300 36100 171400 36200
rect 171300 36200 171400 36300
rect 171300 36300 171400 36400
rect 171300 36400 171400 36500
rect 171400 29700 171500 29800
rect 171400 29800 171500 29900
rect 171400 29900 171500 30000
rect 171400 30000 171500 30100
rect 171400 30100 171500 30200
rect 171400 30200 171500 30300
rect 171400 30300 171500 30400
rect 171400 30400 171500 30500
rect 171400 30500 171500 30600
rect 171400 30600 171500 30700
rect 171400 30700 171500 30800
rect 171400 30800 171500 30900
rect 171400 30900 171500 31000
rect 171400 31000 171500 31100
rect 171400 31100 171500 31200
rect 171400 31200 171500 31300
rect 171400 31300 171500 31400
rect 171400 31400 171500 31500
rect 171400 31500 171500 31600
rect 171400 31600 171500 31700
rect 171400 31700 171500 31800
rect 171400 31800 171500 31900
rect 171400 31900 171500 32000
rect 171400 32000 171500 32100
rect 171400 32100 171500 32200
rect 171400 32200 171500 32300
rect 171400 32300 171500 32400
rect 171400 32400 171500 32500
rect 171400 32500 171500 32600
rect 171400 32600 171500 32700
rect 171400 32700 171500 32800
rect 171400 32800 171500 32900
rect 171400 32900 171500 33000
rect 171400 33000 171500 33100
rect 171400 33100 171500 33200
rect 171400 33200 171500 33300
rect 171400 33300 171500 33400
rect 171400 33400 171500 33500
rect 171400 33500 171500 33600
rect 171400 33600 171500 33700
rect 171400 33700 171500 33800
rect 171400 33800 171500 33900
rect 171400 33900 171500 34000
rect 171400 34000 171500 34100
rect 171400 34100 171500 34200
rect 171400 34200 171500 34300
rect 171400 34300 171500 34400
rect 171400 34400 171500 34500
rect 171400 34500 171500 34600
rect 171400 34600 171500 34700
rect 171400 34700 171500 34800
rect 171400 34800 171500 34900
rect 171400 34900 171500 35000
rect 171400 35000 171500 35100
rect 171400 35100 171500 35200
rect 171400 35200 171500 35300
rect 171400 35300 171500 35400
rect 171400 35400 171500 35500
rect 171400 35500 171500 35600
rect 171400 35600 171500 35700
rect 171400 35700 171500 35800
rect 171400 35800 171500 35900
rect 171400 35900 171500 36000
rect 171400 36000 171500 36100
rect 171400 36100 171500 36200
rect 171400 36200 171500 36300
rect 171400 36300 171500 36400
rect 171400 36400 171500 36500
rect 171400 36500 171500 36600
rect 171400 36600 171500 36700
rect 171500 30000 171600 30100
rect 171500 30100 171600 30200
rect 171500 30200 171600 30300
rect 171500 30300 171600 30400
rect 171500 30400 171600 30500
rect 171500 30500 171600 30600
rect 171500 30600 171600 30700
rect 171500 30700 171600 30800
rect 171500 30800 171600 30900
rect 171500 30900 171600 31000
rect 171500 31000 171600 31100
rect 171500 31100 171600 31200
rect 171500 31200 171600 31300
rect 171500 31300 171600 31400
rect 171500 31400 171600 31500
rect 171500 31500 171600 31600
rect 171500 31600 171600 31700
rect 171500 31700 171600 31800
rect 171500 31800 171600 31900
rect 171500 31900 171600 32000
rect 171500 32000 171600 32100
rect 171500 32100 171600 32200
rect 171500 32200 171600 32300
rect 171500 32300 171600 32400
rect 171500 32400 171600 32500
rect 171500 32500 171600 32600
rect 171500 32600 171600 32700
rect 171500 32700 171600 32800
rect 171500 32800 171600 32900
rect 171500 32900 171600 33000
rect 171500 33000 171600 33100
rect 171500 33100 171600 33200
rect 171500 33200 171600 33300
rect 171500 33300 171600 33400
rect 171500 33400 171600 33500
rect 171500 33500 171600 33600
rect 171500 33600 171600 33700
rect 171500 33700 171600 33800
rect 171500 33800 171600 33900
rect 171500 33900 171600 34000
rect 171500 34000 171600 34100
rect 171500 34100 171600 34200
rect 171500 34200 171600 34300
rect 171500 34300 171600 34400
rect 171500 34400 171600 34500
rect 171500 34500 171600 34600
rect 171500 34600 171600 34700
rect 171500 34700 171600 34800
rect 171500 34800 171600 34900
rect 171500 34900 171600 35000
rect 171500 35000 171600 35100
rect 171500 35100 171600 35200
rect 171500 35200 171600 35300
rect 171500 35300 171600 35400
rect 171500 35400 171600 35500
rect 171500 35500 171600 35600
rect 171500 35600 171600 35700
rect 171500 35700 171600 35800
rect 171500 35800 171600 35900
rect 171500 35900 171600 36000
rect 171500 36000 171600 36100
rect 171500 36100 171600 36200
rect 171500 36200 171600 36300
rect 171500 36300 171600 36400
rect 171500 36400 171600 36500
rect 171500 36500 171600 36600
rect 171500 36600 171600 36700
rect 171500 36700 171600 36800
rect 171600 30300 171700 30400
rect 171600 30400 171700 30500
rect 171600 30500 171700 30600
rect 171600 30600 171700 30700
rect 171600 30700 171700 30800
rect 171600 30800 171700 30900
rect 171600 30900 171700 31000
rect 171600 31000 171700 31100
rect 171600 31100 171700 31200
rect 171600 31200 171700 31300
rect 171600 31300 171700 31400
rect 171600 31400 171700 31500
rect 171600 31500 171700 31600
rect 171600 31600 171700 31700
rect 171600 31700 171700 31800
rect 171600 31800 171700 31900
rect 171600 31900 171700 32000
rect 171600 32000 171700 32100
rect 171600 32100 171700 32200
rect 171600 32200 171700 32300
rect 171600 32300 171700 32400
rect 171600 32400 171700 32500
rect 171600 32500 171700 32600
rect 171600 32600 171700 32700
rect 171600 32700 171700 32800
rect 171600 32800 171700 32900
rect 171600 32900 171700 33000
rect 171600 33000 171700 33100
rect 171600 33100 171700 33200
rect 171600 33200 171700 33300
rect 171600 33300 171700 33400
rect 171600 33400 171700 33500
rect 171600 33500 171700 33600
rect 171600 33600 171700 33700
rect 171600 33700 171700 33800
rect 171600 33800 171700 33900
rect 171600 33900 171700 34000
rect 171600 34000 171700 34100
rect 171600 34100 171700 34200
rect 171600 34200 171700 34300
rect 171600 34300 171700 34400
rect 171600 34400 171700 34500
rect 171600 34500 171700 34600
rect 171600 34600 171700 34700
rect 171600 34700 171700 34800
rect 171600 34800 171700 34900
rect 171600 34900 171700 35000
rect 171600 35000 171700 35100
rect 171600 35100 171700 35200
rect 171600 35200 171700 35300
rect 171600 35300 171700 35400
rect 171600 35400 171700 35500
rect 171600 35500 171700 35600
rect 171600 35600 171700 35700
rect 171600 35700 171700 35800
rect 171600 35800 171700 35900
rect 171600 35900 171700 36000
rect 171600 36000 171700 36100
rect 171600 36100 171700 36200
rect 171600 36200 171700 36300
rect 171600 36300 171700 36400
rect 171600 36400 171700 36500
rect 171600 36500 171700 36600
rect 171600 36600 171700 36700
rect 171600 36700 171700 36800
rect 171600 36800 171700 36900
rect 171600 36900 171700 37000
rect 171700 30600 171800 30700
rect 171700 30700 171800 30800
rect 171700 30800 171800 30900
rect 171700 30900 171800 31000
rect 171700 31000 171800 31100
rect 171700 31100 171800 31200
rect 171700 31200 171800 31300
rect 171700 31300 171800 31400
rect 171700 31400 171800 31500
rect 171700 31500 171800 31600
rect 171700 31600 171800 31700
rect 171700 31700 171800 31800
rect 171700 31800 171800 31900
rect 171700 31900 171800 32000
rect 171700 32000 171800 32100
rect 171700 32100 171800 32200
rect 171700 32200 171800 32300
rect 171700 32300 171800 32400
rect 171700 32400 171800 32500
rect 171700 32500 171800 32600
rect 171700 32600 171800 32700
rect 171700 32700 171800 32800
rect 171700 32800 171800 32900
rect 171700 32900 171800 33000
rect 171700 33000 171800 33100
rect 171700 33100 171800 33200
rect 171700 33200 171800 33300
rect 171700 33300 171800 33400
rect 171700 33400 171800 33500
rect 171700 33500 171800 33600
rect 171700 33600 171800 33700
rect 171700 33700 171800 33800
rect 171700 33800 171800 33900
rect 171700 33900 171800 34000
rect 171700 34000 171800 34100
rect 171700 34100 171800 34200
rect 171700 34200 171800 34300
rect 171700 34300 171800 34400
rect 171700 34400 171800 34500
rect 171700 34500 171800 34600
rect 171700 34600 171800 34700
rect 171700 34700 171800 34800
rect 171700 34800 171800 34900
rect 171700 34900 171800 35000
rect 171700 35000 171800 35100
rect 171700 35100 171800 35200
rect 171700 35200 171800 35300
rect 171700 35300 171800 35400
rect 171700 35400 171800 35500
rect 171700 35500 171800 35600
rect 171700 35600 171800 35700
rect 171700 35700 171800 35800
rect 171700 35800 171800 35900
rect 171700 35900 171800 36000
rect 171700 36000 171800 36100
rect 171700 36100 171800 36200
rect 171700 36200 171800 36300
rect 171700 36300 171800 36400
rect 171700 36400 171800 36500
rect 171700 36500 171800 36600
rect 171700 36600 171800 36700
rect 171700 36700 171800 36800
rect 171700 36800 171800 36900
rect 171700 36900 171800 37000
rect 171700 37000 171800 37100
rect 171700 37100 171800 37200
rect 171800 30900 171900 31000
rect 171800 31000 171900 31100
rect 171800 31100 171900 31200
rect 171800 31200 171900 31300
rect 171800 31300 171900 31400
rect 171800 31400 171900 31500
rect 171800 31500 171900 31600
rect 171800 31600 171900 31700
rect 171800 31700 171900 31800
rect 171800 31800 171900 31900
rect 171800 31900 171900 32000
rect 171800 32000 171900 32100
rect 171800 32100 171900 32200
rect 171800 32200 171900 32300
rect 171800 32300 171900 32400
rect 171800 32400 171900 32500
rect 171800 32500 171900 32600
rect 171800 32600 171900 32700
rect 171800 32700 171900 32800
rect 171800 32800 171900 32900
rect 171800 32900 171900 33000
rect 171800 33000 171900 33100
rect 171800 33100 171900 33200
rect 171800 33200 171900 33300
rect 171800 33300 171900 33400
rect 171800 33400 171900 33500
rect 171800 33500 171900 33600
rect 171800 33600 171900 33700
rect 171800 33700 171900 33800
rect 171800 33800 171900 33900
rect 171800 33900 171900 34000
rect 171800 34000 171900 34100
rect 171800 34100 171900 34200
rect 171800 34200 171900 34300
rect 171800 34300 171900 34400
rect 171800 34400 171900 34500
rect 171800 34500 171900 34600
rect 171800 34600 171900 34700
rect 171800 34700 171900 34800
rect 171800 34800 171900 34900
rect 171800 34900 171900 35000
rect 171800 35000 171900 35100
rect 171800 35100 171900 35200
rect 171800 35200 171900 35300
rect 171800 35300 171900 35400
rect 171800 35400 171900 35500
rect 171800 35500 171900 35600
rect 171800 35600 171900 35700
rect 171800 35700 171900 35800
rect 171800 35800 171900 35900
rect 171800 35900 171900 36000
rect 171800 36000 171900 36100
rect 171800 36100 171900 36200
rect 171800 36200 171900 36300
rect 171800 36300 171900 36400
rect 171800 36400 171900 36500
rect 171800 36500 171900 36600
rect 171800 36600 171900 36700
rect 171800 36700 171900 36800
rect 171800 36800 171900 36900
rect 171800 36900 171900 37000
rect 171800 37000 171900 37100
rect 171800 37100 171900 37200
rect 171800 37200 171900 37300
rect 171900 31200 172000 31300
rect 171900 31300 172000 31400
rect 171900 31400 172000 31500
rect 171900 31500 172000 31600
rect 171900 31600 172000 31700
rect 171900 31700 172000 31800
rect 171900 31800 172000 31900
rect 171900 31900 172000 32000
rect 171900 32000 172000 32100
rect 171900 32100 172000 32200
rect 171900 32200 172000 32300
rect 171900 32300 172000 32400
rect 171900 32400 172000 32500
rect 171900 32500 172000 32600
rect 171900 32600 172000 32700
rect 171900 32700 172000 32800
rect 171900 32800 172000 32900
rect 171900 32900 172000 33000
rect 171900 33000 172000 33100
rect 171900 33100 172000 33200
rect 171900 33200 172000 33300
rect 171900 33300 172000 33400
rect 171900 33400 172000 33500
rect 171900 33500 172000 33600
rect 171900 33600 172000 33700
rect 171900 33700 172000 33800
rect 171900 33800 172000 33900
rect 171900 33900 172000 34000
rect 171900 34000 172000 34100
rect 171900 34100 172000 34200
rect 171900 34200 172000 34300
rect 171900 34300 172000 34400
rect 171900 34400 172000 34500
rect 171900 34500 172000 34600
rect 171900 34600 172000 34700
rect 171900 34700 172000 34800
rect 171900 34800 172000 34900
rect 171900 34900 172000 35000
rect 171900 35000 172000 35100
rect 171900 35100 172000 35200
rect 171900 35200 172000 35300
rect 171900 35300 172000 35400
rect 171900 35400 172000 35500
rect 171900 35500 172000 35600
rect 171900 35600 172000 35700
rect 171900 35700 172000 35800
rect 171900 35800 172000 35900
rect 171900 35900 172000 36000
rect 171900 36000 172000 36100
rect 171900 36100 172000 36200
rect 171900 36200 172000 36300
rect 171900 36300 172000 36400
rect 171900 36400 172000 36500
rect 171900 36500 172000 36600
rect 171900 36600 172000 36700
rect 171900 36700 172000 36800
rect 171900 36800 172000 36900
rect 171900 36900 172000 37000
rect 171900 37000 172000 37100
rect 171900 37100 172000 37200
rect 171900 37200 172000 37300
rect 171900 37300 172000 37400
rect 172000 31600 172100 31700
rect 172000 31700 172100 31800
rect 172000 31800 172100 31900
rect 172000 31900 172100 32000
rect 172000 32000 172100 32100
rect 172000 32100 172100 32200
rect 172000 32200 172100 32300
rect 172000 32300 172100 32400
rect 172000 32400 172100 32500
rect 172000 32500 172100 32600
rect 172000 32600 172100 32700
rect 172000 32700 172100 32800
rect 172000 32800 172100 32900
rect 172000 32900 172100 33000
rect 172000 33000 172100 33100
rect 172000 33100 172100 33200
rect 172000 33200 172100 33300
rect 172000 33300 172100 33400
rect 172000 33400 172100 33500
rect 172000 33500 172100 33600
rect 172000 33600 172100 33700
rect 172000 33700 172100 33800
rect 172000 33800 172100 33900
rect 172000 33900 172100 34000
rect 172000 34000 172100 34100
rect 172000 34100 172100 34200
rect 172000 34200 172100 34300
rect 172000 34300 172100 34400
rect 172000 34400 172100 34500
rect 172000 34500 172100 34600
rect 172000 34600 172100 34700
rect 172000 34700 172100 34800
rect 172000 34800 172100 34900
rect 172000 34900 172100 35000
rect 172000 35000 172100 35100
rect 172000 35100 172100 35200
rect 172000 35200 172100 35300
rect 172000 35300 172100 35400
rect 172000 35400 172100 35500
rect 172000 35500 172100 35600
rect 172000 35600 172100 35700
rect 172000 35700 172100 35800
rect 172000 35800 172100 35900
rect 172000 35900 172100 36000
rect 172000 36000 172100 36100
rect 172000 36100 172100 36200
rect 172000 36200 172100 36300
rect 172000 36300 172100 36400
rect 172000 36400 172100 36500
rect 172000 36500 172100 36600
rect 172000 36600 172100 36700
rect 172000 36700 172100 36800
rect 172000 36800 172100 36900
rect 172000 36900 172100 37000
rect 172000 37000 172100 37100
rect 172000 37100 172100 37200
rect 172000 37200 172100 37300
rect 172000 37300 172100 37400
rect 172000 37400 172100 37500
rect 172000 37500 172100 37600
rect 172100 31900 172200 32000
rect 172100 32000 172200 32100
rect 172100 32100 172200 32200
rect 172100 32200 172200 32300
rect 172100 32300 172200 32400
rect 172100 32400 172200 32500
rect 172100 32500 172200 32600
rect 172100 32600 172200 32700
rect 172100 32700 172200 32800
rect 172100 32800 172200 32900
rect 172100 32900 172200 33000
rect 172100 33000 172200 33100
rect 172100 33100 172200 33200
rect 172100 33200 172200 33300
rect 172100 33300 172200 33400
rect 172100 33400 172200 33500
rect 172100 33500 172200 33600
rect 172100 33600 172200 33700
rect 172100 33700 172200 33800
rect 172100 33800 172200 33900
rect 172100 33900 172200 34000
rect 172100 34000 172200 34100
rect 172100 34100 172200 34200
rect 172100 34200 172200 34300
rect 172100 34300 172200 34400
rect 172100 34400 172200 34500
rect 172100 34500 172200 34600
rect 172100 34600 172200 34700
rect 172100 34700 172200 34800
rect 172100 34800 172200 34900
rect 172100 34900 172200 35000
rect 172100 35000 172200 35100
rect 172100 35100 172200 35200
rect 172100 35200 172200 35300
rect 172100 35300 172200 35400
rect 172100 35400 172200 35500
rect 172100 35500 172200 35600
rect 172100 35600 172200 35700
rect 172100 35700 172200 35800
rect 172100 35800 172200 35900
rect 172100 35900 172200 36000
rect 172100 36000 172200 36100
rect 172100 36100 172200 36200
rect 172100 36200 172200 36300
rect 172100 36300 172200 36400
rect 172100 36400 172200 36500
rect 172100 36500 172200 36600
rect 172100 36600 172200 36700
rect 172100 36700 172200 36800
rect 172100 36800 172200 36900
rect 172100 36900 172200 37000
rect 172100 37000 172200 37100
rect 172100 37100 172200 37200
rect 172100 37200 172200 37300
rect 172100 37300 172200 37400
rect 172100 37400 172200 37500
rect 172100 37500 172200 37600
rect 172100 37600 172200 37700
rect 172200 32200 172300 32300
rect 172200 32300 172300 32400
rect 172200 32400 172300 32500
rect 172200 32500 172300 32600
rect 172200 32600 172300 32700
rect 172200 32700 172300 32800
rect 172200 32800 172300 32900
rect 172200 32900 172300 33000
rect 172200 33000 172300 33100
rect 172200 33100 172300 33200
rect 172200 33200 172300 33300
rect 172200 33300 172300 33400
rect 172200 33400 172300 33500
rect 172200 33500 172300 33600
rect 172200 33600 172300 33700
rect 172200 33700 172300 33800
rect 172200 33800 172300 33900
rect 172200 33900 172300 34000
rect 172200 34000 172300 34100
rect 172200 34100 172300 34200
rect 172200 34200 172300 34300
rect 172200 34300 172300 34400
rect 172200 34400 172300 34500
rect 172200 34500 172300 34600
rect 172200 34600 172300 34700
rect 172200 34700 172300 34800
rect 172200 34800 172300 34900
rect 172200 34900 172300 35000
rect 172200 35000 172300 35100
rect 172200 35100 172300 35200
rect 172200 35200 172300 35300
rect 172200 35300 172300 35400
rect 172200 35400 172300 35500
rect 172200 35500 172300 35600
rect 172200 35600 172300 35700
rect 172200 35700 172300 35800
rect 172200 35800 172300 35900
rect 172200 35900 172300 36000
rect 172200 36000 172300 36100
rect 172200 36100 172300 36200
rect 172200 36200 172300 36300
rect 172200 36300 172300 36400
rect 172200 36400 172300 36500
rect 172200 36500 172300 36600
rect 172200 36600 172300 36700
rect 172200 36700 172300 36800
rect 172200 36800 172300 36900
rect 172200 36900 172300 37000
rect 172200 37000 172300 37100
rect 172200 37100 172300 37200
rect 172200 37200 172300 37300
rect 172200 37300 172300 37400
rect 172200 37400 172300 37500
rect 172200 37500 172300 37600
rect 172200 37600 172300 37700
rect 172300 32600 172400 32700
rect 172300 32700 172400 32800
rect 172300 32800 172400 32900
rect 172300 32900 172400 33000
rect 172300 33000 172400 33100
rect 172300 33100 172400 33200
rect 172300 33200 172400 33300
rect 172300 33300 172400 33400
rect 172300 33400 172400 33500
rect 172300 33500 172400 33600
rect 172300 33600 172400 33700
rect 172300 33700 172400 33800
rect 172300 33800 172400 33900
rect 172300 33900 172400 34000
rect 172300 34000 172400 34100
rect 172300 34100 172400 34200
rect 172300 34200 172400 34300
rect 172300 34300 172400 34400
rect 172300 34400 172400 34500
rect 172300 34500 172400 34600
rect 172300 34600 172400 34700
rect 172300 34700 172400 34800
rect 172300 34800 172400 34900
rect 172300 34900 172400 35000
rect 172300 35000 172400 35100
rect 172300 35100 172400 35200
rect 172300 35200 172400 35300
rect 172300 35300 172400 35400
rect 172300 35400 172400 35500
rect 172300 35500 172400 35600
rect 172300 35600 172400 35700
rect 172300 35700 172400 35800
rect 172300 35800 172400 35900
rect 172300 35900 172400 36000
rect 172300 36000 172400 36100
rect 172300 36100 172400 36200
rect 172300 36200 172400 36300
rect 172300 36300 172400 36400
rect 172300 36400 172400 36500
rect 172300 36500 172400 36600
rect 172300 36600 172400 36700
rect 172300 36700 172400 36800
rect 172300 36800 172400 36900
rect 172300 36900 172400 37000
rect 172300 37000 172400 37100
rect 172300 37100 172400 37200
rect 172300 37200 172400 37300
rect 172300 37300 172400 37400
rect 172300 37400 172400 37500
rect 172300 37500 172400 37600
rect 172300 37600 172400 37700
rect 172300 37700 172400 37800
rect 172400 32900 172500 33000
rect 172400 33000 172500 33100
rect 172400 33100 172500 33200
rect 172400 33200 172500 33300
rect 172400 33300 172500 33400
rect 172400 33400 172500 33500
rect 172400 33500 172500 33600
rect 172400 33600 172500 33700
rect 172400 33700 172500 33800
rect 172400 33800 172500 33900
rect 172400 33900 172500 34000
rect 172400 34000 172500 34100
rect 172400 34100 172500 34200
rect 172400 34200 172500 34300
rect 172400 34300 172500 34400
rect 172400 34400 172500 34500
rect 172400 34500 172500 34600
rect 172400 34600 172500 34700
rect 172400 34700 172500 34800
rect 172400 34800 172500 34900
rect 172400 34900 172500 35000
rect 172400 35000 172500 35100
rect 172400 35100 172500 35200
rect 172400 35200 172500 35300
rect 172400 35300 172500 35400
rect 172400 35400 172500 35500
rect 172400 35500 172500 35600
rect 172400 35600 172500 35700
rect 172400 35700 172500 35800
rect 172400 35800 172500 35900
rect 172400 35900 172500 36000
rect 172400 36000 172500 36100
rect 172400 36100 172500 36200
rect 172400 36200 172500 36300
rect 172400 36300 172500 36400
rect 172400 36400 172500 36500
rect 172400 36500 172500 36600
rect 172400 36600 172500 36700
rect 172400 36700 172500 36800
rect 172400 36800 172500 36900
rect 172400 36900 172500 37000
rect 172400 37000 172500 37100
rect 172400 37100 172500 37200
rect 172400 37200 172500 37300
rect 172400 37300 172500 37400
rect 172400 37400 172500 37500
rect 172400 37500 172500 37600
rect 172400 37600 172500 37700
rect 172400 37700 172500 37800
rect 172400 37800 172500 37900
rect 172500 33300 172600 33400
rect 172500 33400 172600 33500
rect 172500 33500 172600 33600
rect 172500 33600 172600 33700
rect 172500 33700 172600 33800
rect 172500 33800 172600 33900
rect 172500 33900 172600 34000
rect 172500 34000 172600 34100
rect 172500 34100 172600 34200
rect 172500 34200 172600 34300
rect 172500 34300 172600 34400
rect 172500 34400 172600 34500
rect 172500 34500 172600 34600
rect 172500 34600 172600 34700
rect 172500 34700 172600 34800
rect 172500 34800 172600 34900
rect 172500 34900 172600 35000
rect 172500 35000 172600 35100
rect 172500 35100 172600 35200
rect 172500 35200 172600 35300
rect 172500 35300 172600 35400
rect 172500 35400 172600 35500
rect 172500 35500 172600 35600
rect 172500 35600 172600 35700
rect 172500 35700 172600 35800
rect 172500 35800 172600 35900
rect 172500 35900 172600 36000
rect 172500 36000 172600 36100
rect 172500 36100 172600 36200
rect 172500 36200 172600 36300
rect 172500 36300 172600 36400
rect 172500 36400 172600 36500
rect 172500 36500 172600 36600
rect 172500 36600 172600 36700
rect 172500 36700 172600 36800
rect 172500 36800 172600 36900
rect 172500 36900 172600 37000
rect 172500 37000 172600 37100
rect 172500 37100 172600 37200
rect 172500 37200 172600 37300
rect 172500 37300 172600 37400
rect 172500 37400 172600 37500
rect 172500 37500 172600 37600
rect 172500 37600 172600 37700
rect 172500 37700 172600 37800
rect 172500 37800 172600 37900
rect 172600 32900 172700 33000
rect 172600 33000 172700 33100
rect 172600 33100 172700 33200
rect 172600 33200 172700 33300
rect 172600 33300 172700 33400
rect 172600 33400 172700 33500
rect 172600 33500 172700 33600
rect 172600 33600 172700 33700
rect 172600 33700 172700 33800
rect 172600 33800 172700 33900
rect 172600 33900 172700 34000
rect 172600 34000 172700 34100
rect 172600 34100 172700 34200
rect 172600 34200 172700 34300
rect 172600 34300 172700 34400
rect 172600 34400 172700 34500
rect 172600 34500 172700 34600
rect 172600 34600 172700 34700
rect 172600 34700 172700 34800
rect 172600 34800 172700 34900
rect 172600 34900 172700 35000
rect 172600 35000 172700 35100
rect 172600 35100 172700 35200
rect 172600 35200 172700 35300
rect 172600 35300 172700 35400
rect 172600 35400 172700 35500
rect 172600 35500 172700 35600
rect 172600 35600 172700 35700
rect 172600 35700 172700 35800
rect 172600 35800 172700 35900
rect 172600 35900 172700 36000
rect 172600 36000 172700 36100
rect 172600 36100 172700 36200
rect 172600 36200 172700 36300
rect 172600 36300 172700 36400
rect 172600 36400 172700 36500
rect 172600 36500 172700 36600
rect 172600 36600 172700 36700
rect 172600 36700 172700 36800
rect 172600 36800 172700 36900
rect 172600 36900 172700 37000
rect 172600 37000 172700 37100
rect 172600 37100 172700 37200
rect 172600 37200 172700 37300
rect 172600 37300 172700 37400
rect 172600 37400 172700 37500
rect 172600 37500 172700 37600
rect 172600 37600 172700 37700
rect 172600 37700 172700 37800
rect 172600 37800 172700 37900
rect 172600 37900 172700 38000
rect 172700 32200 172800 32300
rect 172700 32300 172800 32400
rect 172700 32400 172800 32500
rect 172700 32500 172800 32600
rect 172700 32600 172800 32700
rect 172700 32700 172800 32800
rect 172700 32800 172800 32900
rect 172700 32900 172800 33000
rect 172700 33000 172800 33100
rect 172700 33100 172800 33200
rect 172700 33200 172800 33300
rect 172700 33300 172800 33400
rect 172700 33400 172800 33500
rect 172700 33500 172800 33600
rect 172700 33600 172800 33700
rect 172700 33700 172800 33800
rect 172700 33800 172800 33900
rect 172700 33900 172800 34000
rect 172700 34000 172800 34100
rect 172700 34100 172800 34200
rect 172700 34200 172800 34300
rect 172700 34300 172800 34400
rect 172700 34400 172800 34500
rect 172700 34500 172800 34600
rect 172700 34600 172800 34700
rect 172700 34700 172800 34800
rect 172700 34800 172800 34900
rect 172700 34900 172800 35000
rect 172700 35000 172800 35100
rect 172700 35100 172800 35200
rect 172700 35200 172800 35300
rect 172700 35300 172800 35400
rect 172700 35400 172800 35500
rect 172700 35500 172800 35600
rect 172700 35600 172800 35700
rect 172700 35700 172800 35800
rect 172700 35800 172800 35900
rect 172700 35900 172800 36000
rect 172700 36000 172800 36100
rect 172700 36100 172800 36200
rect 172700 36200 172800 36300
rect 172700 36300 172800 36400
rect 172700 36400 172800 36500
rect 172700 36500 172800 36600
rect 172700 36600 172800 36700
rect 172700 36700 172800 36800
rect 172700 36800 172800 36900
rect 172700 36900 172800 37000
rect 172700 37000 172800 37100
rect 172700 37100 172800 37200
rect 172700 37200 172800 37300
rect 172700 37300 172800 37400
rect 172700 37400 172800 37500
rect 172700 37500 172800 37600
rect 172700 37600 172800 37700
rect 172700 37700 172800 37800
rect 172700 37800 172800 37900
rect 172700 37900 172800 38000
rect 172800 31500 172900 31600
rect 172800 31600 172900 31700
rect 172800 31700 172900 31800
rect 172800 31800 172900 31900
rect 172800 31900 172900 32000
rect 172800 32000 172900 32100
rect 172800 32100 172900 32200
rect 172800 32200 172900 32300
rect 172800 32300 172900 32400
rect 172800 32400 172900 32500
rect 172800 32500 172900 32600
rect 172800 32600 172900 32700
rect 172800 32700 172900 32800
rect 172800 32800 172900 32900
rect 172800 32900 172900 33000
rect 172800 33000 172900 33100
rect 172800 33100 172900 33200
rect 172800 33200 172900 33300
rect 172800 33300 172900 33400
rect 172800 33400 172900 33500
rect 172800 33500 172900 33600
rect 172800 33600 172900 33700
rect 172800 33700 172900 33800
rect 172800 33800 172900 33900
rect 172800 33900 172900 34000
rect 172800 34000 172900 34100
rect 172800 34100 172900 34200
rect 172800 34200 172900 34300
rect 172800 34300 172900 34400
rect 172800 34400 172900 34500
rect 172800 34500 172900 34600
rect 172800 34600 172900 34700
rect 172800 34700 172900 34800
rect 172800 34800 172900 34900
rect 172800 34900 172900 35000
rect 172800 35000 172900 35100
rect 172800 35100 172900 35200
rect 172800 35200 172900 35300
rect 172800 35300 172900 35400
rect 172800 35400 172900 35500
rect 172800 35500 172900 35600
rect 172800 35600 172900 35700
rect 172800 35700 172900 35800
rect 172800 35800 172900 35900
rect 172800 35900 172900 36000
rect 172800 36000 172900 36100
rect 172800 36100 172900 36200
rect 172800 36200 172900 36300
rect 172800 36300 172900 36400
rect 172800 36400 172900 36500
rect 172800 36500 172900 36600
rect 172800 36600 172900 36700
rect 172800 36700 172900 36800
rect 172800 36800 172900 36900
rect 172800 36900 172900 37000
rect 172800 37000 172900 37100
rect 172800 37100 172900 37200
rect 172800 37200 172900 37300
rect 172800 37300 172900 37400
rect 172800 37400 172900 37500
rect 172800 37500 172900 37600
rect 172800 37600 172900 37700
rect 172800 37700 172900 37800
rect 172800 37800 172900 37900
rect 172800 37900 172900 38000
rect 172900 30900 173000 31000
rect 172900 31000 173000 31100
rect 172900 31100 173000 31200
rect 172900 31200 173000 31300
rect 172900 31300 173000 31400
rect 172900 31400 173000 31500
rect 172900 31500 173000 31600
rect 172900 31600 173000 31700
rect 172900 31700 173000 31800
rect 172900 31800 173000 31900
rect 172900 31900 173000 32000
rect 172900 32000 173000 32100
rect 172900 32100 173000 32200
rect 172900 32200 173000 32300
rect 172900 32300 173000 32400
rect 172900 32400 173000 32500
rect 172900 32500 173000 32600
rect 172900 32600 173000 32700
rect 172900 32700 173000 32800
rect 172900 32800 173000 32900
rect 172900 32900 173000 33000
rect 172900 33000 173000 33100
rect 172900 33100 173000 33200
rect 172900 33200 173000 33300
rect 172900 33300 173000 33400
rect 172900 33400 173000 33500
rect 172900 33500 173000 33600
rect 172900 33600 173000 33700
rect 172900 33700 173000 33800
rect 172900 33800 173000 33900
rect 172900 33900 173000 34000
rect 172900 34000 173000 34100
rect 172900 34100 173000 34200
rect 172900 34200 173000 34300
rect 172900 34300 173000 34400
rect 172900 34400 173000 34500
rect 172900 34500 173000 34600
rect 172900 34600 173000 34700
rect 172900 34700 173000 34800
rect 172900 34800 173000 34900
rect 172900 34900 173000 35000
rect 172900 35000 173000 35100
rect 172900 35100 173000 35200
rect 172900 35200 173000 35300
rect 172900 35300 173000 35400
rect 172900 35400 173000 35500
rect 172900 35500 173000 35600
rect 172900 35600 173000 35700
rect 172900 35700 173000 35800
rect 172900 35800 173000 35900
rect 172900 35900 173000 36000
rect 172900 36000 173000 36100
rect 172900 36100 173000 36200
rect 172900 36200 173000 36300
rect 172900 36300 173000 36400
rect 172900 36400 173000 36500
rect 172900 36500 173000 36600
rect 172900 36600 173000 36700
rect 172900 36700 173000 36800
rect 172900 36800 173000 36900
rect 172900 36900 173000 37000
rect 172900 37000 173000 37100
rect 172900 37100 173000 37200
rect 172900 37200 173000 37300
rect 172900 37300 173000 37400
rect 172900 37400 173000 37500
rect 172900 37500 173000 37600
rect 172900 37600 173000 37700
rect 172900 37700 173000 37800
rect 172900 37800 173000 37900
rect 172900 37900 173000 38000
rect 173000 30300 173100 30400
rect 173000 30400 173100 30500
rect 173000 30500 173100 30600
rect 173000 30600 173100 30700
rect 173000 30700 173100 30800
rect 173000 30800 173100 30900
rect 173000 30900 173100 31000
rect 173000 31000 173100 31100
rect 173000 31100 173100 31200
rect 173000 31200 173100 31300
rect 173000 31300 173100 31400
rect 173000 31400 173100 31500
rect 173000 31500 173100 31600
rect 173000 31600 173100 31700
rect 173000 31700 173100 31800
rect 173000 31800 173100 31900
rect 173000 31900 173100 32000
rect 173000 32000 173100 32100
rect 173000 32100 173100 32200
rect 173000 32200 173100 32300
rect 173000 32300 173100 32400
rect 173000 32400 173100 32500
rect 173000 32500 173100 32600
rect 173000 32600 173100 32700
rect 173000 32700 173100 32800
rect 173000 32800 173100 32900
rect 173000 32900 173100 33000
rect 173000 33000 173100 33100
rect 173000 33100 173100 33200
rect 173000 33200 173100 33300
rect 173000 33300 173100 33400
rect 173000 33400 173100 33500
rect 173000 33500 173100 33600
rect 173000 33600 173100 33700
rect 173000 33700 173100 33800
rect 173000 33800 173100 33900
rect 173000 33900 173100 34000
rect 173000 34000 173100 34100
rect 173000 34100 173100 34200
rect 173000 34200 173100 34300
rect 173000 34300 173100 34400
rect 173000 34400 173100 34500
rect 173000 34500 173100 34600
rect 173000 34600 173100 34700
rect 173000 34700 173100 34800
rect 173000 34800 173100 34900
rect 173000 34900 173100 35000
rect 173000 35000 173100 35100
rect 173000 35100 173100 35200
rect 173000 35200 173100 35300
rect 173000 35300 173100 35400
rect 173000 35400 173100 35500
rect 173000 35500 173100 35600
rect 173000 35600 173100 35700
rect 173000 35700 173100 35800
rect 173000 35800 173100 35900
rect 173000 35900 173100 36000
rect 173000 36000 173100 36100
rect 173000 36100 173100 36200
rect 173000 36200 173100 36300
rect 173000 36300 173100 36400
rect 173000 36400 173100 36500
rect 173000 36500 173100 36600
rect 173000 36600 173100 36700
rect 173000 36700 173100 36800
rect 173000 36800 173100 36900
rect 173000 36900 173100 37000
rect 173000 37000 173100 37100
rect 173000 37100 173100 37200
rect 173000 37200 173100 37300
rect 173000 37300 173100 37400
rect 173000 37400 173100 37500
rect 173000 37500 173100 37600
rect 173000 37600 173100 37700
rect 173000 37700 173100 37800
rect 173000 37800 173100 37900
rect 173000 37900 173100 38000
rect 173100 29800 173200 29900
rect 173100 29900 173200 30000
rect 173100 30000 173200 30100
rect 173100 30100 173200 30200
rect 173100 30200 173200 30300
rect 173100 30300 173200 30400
rect 173100 30400 173200 30500
rect 173100 30500 173200 30600
rect 173100 30600 173200 30700
rect 173100 30700 173200 30800
rect 173100 30800 173200 30900
rect 173100 30900 173200 31000
rect 173100 31000 173200 31100
rect 173100 31100 173200 31200
rect 173100 31200 173200 31300
rect 173100 31300 173200 31400
rect 173100 31400 173200 31500
rect 173100 31500 173200 31600
rect 173100 31600 173200 31700
rect 173100 31700 173200 31800
rect 173100 31800 173200 31900
rect 173100 31900 173200 32000
rect 173100 32000 173200 32100
rect 173100 32100 173200 32200
rect 173100 32200 173200 32300
rect 173100 32300 173200 32400
rect 173100 32400 173200 32500
rect 173100 32500 173200 32600
rect 173100 32600 173200 32700
rect 173100 32700 173200 32800
rect 173100 32800 173200 32900
rect 173100 32900 173200 33000
rect 173100 33000 173200 33100
rect 173100 33100 173200 33200
rect 173100 33200 173200 33300
rect 173100 33300 173200 33400
rect 173100 33400 173200 33500
rect 173100 33500 173200 33600
rect 173100 33600 173200 33700
rect 173100 33700 173200 33800
rect 173100 33800 173200 33900
rect 173100 33900 173200 34000
rect 173100 34000 173200 34100
rect 173100 34100 173200 34200
rect 173100 34200 173200 34300
rect 173100 34300 173200 34400
rect 173100 34400 173200 34500
rect 173100 34500 173200 34600
rect 173100 34600 173200 34700
rect 173100 34700 173200 34800
rect 173100 34800 173200 34900
rect 173100 34900 173200 35000
rect 173100 35000 173200 35100
rect 173100 35100 173200 35200
rect 173100 35200 173200 35300
rect 173100 35300 173200 35400
rect 173100 35400 173200 35500
rect 173100 35500 173200 35600
rect 173100 35600 173200 35700
rect 173100 35700 173200 35800
rect 173100 35800 173200 35900
rect 173100 35900 173200 36000
rect 173100 36000 173200 36100
rect 173100 36100 173200 36200
rect 173100 36200 173200 36300
rect 173100 36300 173200 36400
rect 173100 36400 173200 36500
rect 173100 36500 173200 36600
rect 173100 36600 173200 36700
rect 173100 36700 173200 36800
rect 173100 36800 173200 36900
rect 173100 36900 173200 37000
rect 173100 37000 173200 37100
rect 173100 37100 173200 37200
rect 173100 37200 173200 37300
rect 173100 37300 173200 37400
rect 173100 37400 173200 37500
rect 173100 37500 173200 37600
rect 173100 37600 173200 37700
rect 173100 37700 173200 37800
rect 173100 37800 173200 37900
rect 173200 29200 173300 29300
rect 173200 29300 173300 29400
rect 173200 29400 173300 29500
rect 173200 29500 173300 29600
rect 173200 29600 173300 29700
rect 173200 29700 173300 29800
rect 173200 29800 173300 29900
rect 173200 29900 173300 30000
rect 173200 30000 173300 30100
rect 173200 30100 173300 30200
rect 173200 30200 173300 30300
rect 173200 30300 173300 30400
rect 173200 30400 173300 30500
rect 173200 30500 173300 30600
rect 173200 30600 173300 30700
rect 173200 30700 173300 30800
rect 173200 30800 173300 30900
rect 173200 30900 173300 31000
rect 173200 31000 173300 31100
rect 173200 31100 173300 31200
rect 173200 31200 173300 31300
rect 173200 31300 173300 31400
rect 173200 31400 173300 31500
rect 173200 31500 173300 31600
rect 173200 31600 173300 31700
rect 173200 31700 173300 31800
rect 173200 31800 173300 31900
rect 173200 31900 173300 32000
rect 173200 32000 173300 32100
rect 173200 32100 173300 32200
rect 173200 32200 173300 32300
rect 173200 32300 173300 32400
rect 173200 32400 173300 32500
rect 173200 32500 173300 32600
rect 173200 32600 173300 32700
rect 173200 32700 173300 32800
rect 173200 32800 173300 32900
rect 173200 32900 173300 33000
rect 173200 33000 173300 33100
rect 173200 33100 173300 33200
rect 173200 33200 173300 33300
rect 173200 33300 173300 33400
rect 173200 33400 173300 33500
rect 173200 33500 173300 33600
rect 173200 33600 173300 33700
rect 173200 33700 173300 33800
rect 173200 33800 173300 33900
rect 173200 33900 173300 34000
rect 173200 34000 173300 34100
rect 173200 34100 173300 34200
rect 173200 34200 173300 34300
rect 173200 34300 173300 34400
rect 173200 34400 173300 34500
rect 173200 34500 173300 34600
rect 173200 34600 173300 34700
rect 173200 34700 173300 34800
rect 173200 34800 173300 34900
rect 173200 34900 173300 35000
rect 173200 35000 173300 35100
rect 173200 35100 173300 35200
rect 173200 35200 173300 35300
rect 173200 35300 173300 35400
rect 173200 35400 173300 35500
rect 173200 35500 173300 35600
rect 173200 35600 173300 35700
rect 173200 35700 173300 35800
rect 173200 35800 173300 35900
rect 173200 35900 173300 36000
rect 173200 36000 173300 36100
rect 173200 36100 173300 36200
rect 173200 36200 173300 36300
rect 173200 36300 173300 36400
rect 173200 36400 173300 36500
rect 173200 36500 173300 36600
rect 173200 36600 173300 36700
rect 173200 36700 173300 36800
rect 173200 36800 173300 36900
rect 173200 36900 173300 37000
rect 173200 37000 173300 37100
rect 173200 37100 173300 37200
rect 173200 37200 173300 37300
rect 173200 37300 173300 37400
rect 173200 37400 173300 37500
rect 173200 37500 173300 37600
rect 173200 37600 173300 37700
rect 173200 37700 173300 37800
rect 173200 37800 173300 37900
rect 173300 28700 173400 28800
rect 173300 28800 173400 28900
rect 173300 28900 173400 29000
rect 173300 29000 173400 29100
rect 173300 29100 173400 29200
rect 173300 29200 173400 29300
rect 173300 29300 173400 29400
rect 173300 29400 173400 29500
rect 173300 29500 173400 29600
rect 173300 29600 173400 29700
rect 173300 29700 173400 29800
rect 173300 29800 173400 29900
rect 173300 29900 173400 30000
rect 173300 30000 173400 30100
rect 173300 30100 173400 30200
rect 173300 30200 173400 30300
rect 173300 30300 173400 30400
rect 173300 30400 173400 30500
rect 173300 30500 173400 30600
rect 173300 30600 173400 30700
rect 173300 30700 173400 30800
rect 173300 30800 173400 30900
rect 173300 30900 173400 31000
rect 173300 31000 173400 31100
rect 173300 31100 173400 31200
rect 173300 31200 173400 31300
rect 173300 31300 173400 31400
rect 173300 31400 173400 31500
rect 173300 31500 173400 31600
rect 173300 31600 173400 31700
rect 173300 31700 173400 31800
rect 173300 31800 173400 31900
rect 173300 31900 173400 32000
rect 173300 32000 173400 32100
rect 173300 32100 173400 32200
rect 173300 32200 173400 32300
rect 173300 32300 173400 32400
rect 173300 32400 173400 32500
rect 173300 32500 173400 32600
rect 173300 32600 173400 32700
rect 173300 32700 173400 32800
rect 173300 32800 173400 32900
rect 173300 32900 173400 33000
rect 173300 33000 173400 33100
rect 173300 33100 173400 33200
rect 173300 33200 173400 33300
rect 173300 33300 173400 33400
rect 173300 33400 173400 33500
rect 173300 33500 173400 33600
rect 173300 33600 173400 33700
rect 173300 33700 173400 33800
rect 173300 33800 173400 33900
rect 173300 33900 173400 34000
rect 173300 34000 173400 34100
rect 173300 34100 173400 34200
rect 173300 34200 173400 34300
rect 173300 34300 173400 34400
rect 173300 34400 173400 34500
rect 173300 34500 173400 34600
rect 173300 34600 173400 34700
rect 173300 34700 173400 34800
rect 173300 34800 173400 34900
rect 173300 34900 173400 35000
rect 173300 35000 173400 35100
rect 173300 35100 173400 35200
rect 173300 35200 173400 35300
rect 173300 35300 173400 35400
rect 173300 35400 173400 35500
rect 173300 35500 173400 35600
rect 173300 35600 173400 35700
rect 173300 35700 173400 35800
rect 173300 35800 173400 35900
rect 173300 35900 173400 36000
rect 173300 36000 173400 36100
rect 173300 36100 173400 36200
rect 173300 36200 173400 36300
rect 173300 36300 173400 36400
rect 173300 36400 173400 36500
rect 173300 36500 173400 36600
rect 173300 36600 173400 36700
rect 173300 36700 173400 36800
rect 173300 36800 173400 36900
rect 173300 36900 173400 37000
rect 173300 37000 173400 37100
rect 173300 37100 173400 37200
rect 173300 37200 173400 37300
rect 173300 37300 173400 37400
rect 173300 37400 173400 37500
rect 173300 37500 173400 37600
rect 173300 37600 173400 37700
rect 173300 37700 173400 37800
rect 173300 37800 173400 37900
rect 173400 28100 173500 28200
rect 173400 28200 173500 28300
rect 173400 28300 173500 28400
rect 173400 28400 173500 28500
rect 173400 28500 173500 28600
rect 173400 28600 173500 28700
rect 173400 28700 173500 28800
rect 173400 28800 173500 28900
rect 173400 28900 173500 29000
rect 173400 29000 173500 29100
rect 173400 29100 173500 29200
rect 173400 29200 173500 29300
rect 173400 29300 173500 29400
rect 173400 29400 173500 29500
rect 173400 29500 173500 29600
rect 173400 29600 173500 29700
rect 173400 29700 173500 29800
rect 173400 29800 173500 29900
rect 173400 29900 173500 30000
rect 173400 30000 173500 30100
rect 173400 30100 173500 30200
rect 173400 30200 173500 30300
rect 173400 30300 173500 30400
rect 173400 30400 173500 30500
rect 173400 30500 173500 30600
rect 173400 30600 173500 30700
rect 173400 30700 173500 30800
rect 173400 30800 173500 30900
rect 173400 30900 173500 31000
rect 173400 31000 173500 31100
rect 173400 31100 173500 31200
rect 173400 31200 173500 31300
rect 173400 31300 173500 31400
rect 173400 31400 173500 31500
rect 173400 31500 173500 31600
rect 173400 31600 173500 31700
rect 173400 31700 173500 31800
rect 173400 31800 173500 31900
rect 173400 31900 173500 32000
rect 173400 32000 173500 32100
rect 173400 32100 173500 32200
rect 173400 32200 173500 32300
rect 173400 32300 173500 32400
rect 173400 32400 173500 32500
rect 173400 32500 173500 32600
rect 173400 32600 173500 32700
rect 173400 32700 173500 32800
rect 173400 32800 173500 32900
rect 173400 32900 173500 33000
rect 173400 33000 173500 33100
rect 173400 33100 173500 33200
rect 173400 33200 173500 33300
rect 173400 33300 173500 33400
rect 173400 33400 173500 33500
rect 173400 33500 173500 33600
rect 173400 33600 173500 33700
rect 173400 33700 173500 33800
rect 173400 33800 173500 33900
rect 173400 33900 173500 34000
rect 173400 34000 173500 34100
rect 173400 34100 173500 34200
rect 173400 34200 173500 34300
rect 173400 34300 173500 34400
rect 173400 34400 173500 34500
rect 173400 34500 173500 34600
rect 173400 34600 173500 34700
rect 173400 34700 173500 34800
rect 173400 34800 173500 34900
rect 173400 34900 173500 35000
rect 173400 35000 173500 35100
rect 173400 35100 173500 35200
rect 173400 35200 173500 35300
rect 173400 35300 173500 35400
rect 173400 35400 173500 35500
rect 173400 35500 173500 35600
rect 173400 35600 173500 35700
rect 173400 35700 173500 35800
rect 173400 35800 173500 35900
rect 173400 35900 173500 36000
rect 173400 36000 173500 36100
rect 173400 36100 173500 36200
rect 173400 36200 173500 36300
rect 173400 36300 173500 36400
rect 173400 36400 173500 36500
rect 173400 36500 173500 36600
rect 173400 36600 173500 36700
rect 173400 36700 173500 36800
rect 173400 36800 173500 36900
rect 173400 36900 173500 37000
rect 173400 37000 173500 37100
rect 173400 37100 173500 37200
rect 173400 37200 173500 37300
rect 173400 37300 173500 37400
rect 173400 37400 173500 37500
rect 173400 37500 173500 37600
rect 173400 37600 173500 37700
rect 173400 37700 173500 37800
rect 173500 27600 173600 27700
rect 173500 27700 173600 27800
rect 173500 27800 173600 27900
rect 173500 27900 173600 28000
rect 173500 28000 173600 28100
rect 173500 28100 173600 28200
rect 173500 28200 173600 28300
rect 173500 28300 173600 28400
rect 173500 28400 173600 28500
rect 173500 28500 173600 28600
rect 173500 28600 173600 28700
rect 173500 28700 173600 28800
rect 173500 28800 173600 28900
rect 173500 28900 173600 29000
rect 173500 29000 173600 29100
rect 173500 29100 173600 29200
rect 173500 29200 173600 29300
rect 173500 29300 173600 29400
rect 173500 29400 173600 29500
rect 173500 29500 173600 29600
rect 173500 29600 173600 29700
rect 173500 29700 173600 29800
rect 173500 29800 173600 29900
rect 173500 29900 173600 30000
rect 173500 30000 173600 30100
rect 173500 30100 173600 30200
rect 173500 30200 173600 30300
rect 173500 30300 173600 30400
rect 173500 30400 173600 30500
rect 173500 30500 173600 30600
rect 173500 30600 173600 30700
rect 173500 30700 173600 30800
rect 173500 30800 173600 30900
rect 173500 30900 173600 31000
rect 173500 31000 173600 31100
rect 173500 31100 173600 31200
rect 173500 31200 173600 31300
rect 173500 31300 173600 31400
rect 173500 31400 173600 31500
rect 173500 31500 173600 31600
rect 173500 31600 173600 31700
rect 173500 31700 173600 31800
rect 173500 31800 173600 31900
rect 173500 31900 173600 32000
rect 173500 32000 173600 32100
rect 173500 32100 173600 32200
rect 173500 32200 173600 32300
rect 173500 32300 173600 32400
rect 173500 32400 173600 32500
rect 173500 32500 173600 32600
rect 173500 32600 173600 32700
rect 173500 32700 173600 32800
rect 173500 32800 173600 32900
rect 173500 32900 173600 33000
rect 173500 33000 173600 33100
rect 173500 33100 173600 33200
rect 173500 33200 173600 33300
rect 173500 33300 173600 33400
rect 173500 33400 173600 33500
rect 173500 33500 173600 33600
rect 173500 33600 173600 33700
rect 173500 33700 173600 33800
rect 173500 33800 173600 33900
rect 173500 33900 173600 34000
rect 173500 34000 173600 34100
rect 173500 34100 173600 34200
rect 173500 34200 173600 34300
rect 173500 34300 173600 34400
rect 173500 34400 173600 34500
rect 173500 34500 173600 34600
rect 173500 34600 173600 34700
rect 173500 34700 173600 34800
rect 173500 34800 173600 34900
rect 173500 34900 173600 35000
rect 173500 35000 173600 35100
rect 173500 35100 173600 35200
rect 173500 35200 173600 35300
rect 173500 35300 173600 35400
rect 173500 35400 173600 35500
rect 173500 35500 173600 35600
rect 173500 35600 173600 35700
rect 173500 35700 173600 35800
rect 173500 35800 173600 35900
rect 173500 35900 173600 36000
rect 173500 36000 173600 36100
rect 173500 36100 173600 36200
rect 173500 36200 173600 36300
rect 173500 36300 173600 36400
rect 173500 36400 173600 36500
rect 173500 36500 173600 36600
rect 173500 36600 173600 36700
rect 173500 36700 173600 36800
rect 173500 36800 173600 36900
rect 173500 36900 173600 37000
rect 173500 37000 173600 37100
rect 173500 37100 173600 37200
rect 173500 37200 173600 37300
rect 173500 37300 173600 37400
rect 173500 37400 173600 37500
rect 173500 37500 173600 37600
rect 173500 37600 173600 37700
rect 173600 27100 173700 27200
rect 173600 27200 173700 27300
rect 173600 27300 173700 27400
rect 173600 27400 173700 27500
rect 173600 27500 173700 27600
rect 173600 27600 173700 27700
rect 173600 27700 173700 27800
rect 173600 27800 173700 27900
rect 173600 27900 173700 28000
rect 173600 28000 173700 28100
rect 173600 28100 173700 28200
rect 173600 28200 173700 28300
rect 173600 28300 173700 28400
rect 173600 28400 173700 28500
rect 173600 28500 173700 28600
rect 173600 28600 173700 28700
rect 173600 28700 173700 28800
rect 173600 28800 173700 28900
rect 173600 28900 173700 29000
rect 173600 29000 173700 29100
rect 173600 29100 173700 29200
rect 173600 29200 173700 29300
rect 173600 29300 173700 29400
rect 173600 29400 173700 29500
rect 173600 29500 173700 29600
rect 173600 29600 173700 29700
rect 173600 29700 173700 29800
rect 173600 29800 173700 29900
rect 173600 29900 173700 30000
rect 173600 30000 173700 30100
rect 173600 30100 173700 30200
rect 173600 30200 173700 30300
rect 173600 30300 173700 30400
rect 173600 30400 173700 30500
rect 173600 30500 173700 30600
rect 173600 30600 173700 30700
rect 173600 30700 173700 30800
rect 173600 30800 173700 30900
rect 173600 30900 173700 31000
rect 173600 31000 173700 31100
rect 173600 31100 173700 31200
rect 173600 31200 173700 31300
rect 173600 31300 173700 31400
rect 173600 31400 173700 31500
rect 173600 31500 173700 31600
rect 173600 31600 173700 31700
rect 173600 31700 173700 31800
rect 173600 31800 173700 31900
rect 173600 31900 173700 32000
rect 173600 32000 173700 32100
rect 173600 32100 173700 32200
rect 173600 32200 173700 32300
rect 173600 32300 173700 32400
rect 173600 32400 173700 32500
rect 173600 32500 173700 32600
rect 173600 32600 173700 32700
rect 173600 32700 173700 32800
rect 173600 32800 173700 32900
rect 173600 32900 173700 33000
rect 173600 33000 173700 33100
rect 173600 33100 173700 33200
rect 173600 33200 173700 33300
rect 173600 33300 173700 33400
rect 173600 33400 173700 33500
rect 173600 33500 173700 33600
rect 173600 33600 173700 33700
rect 173600 33700 173700 33800
rect 173600 33800 173700 33900
rect 173600 33900 173700 34000
rect 173600 34000 173700 34100
rect 173600 34100 173700 34200
rect 173600 34200 173700 34300
rect 173600 34300 173700 34400
rect 173600 34400 173700 34500
rect 173600 34500 173700 34600
rect 173600 34600 173700 34700
rect 173600 34700 173700 34800
rect 173600 34800 173700 34900
rect 173600 34900 173700 35000
rect 173600 35000 173700 35100
rect 173600 35100 173700 35200
rect 173600 35200 173700 35300
rect 173600 35300 173700 35400
rect 173600 35400 173700 35500
rect 173600 35500 173700 35600
rect 173600 35600 173700 35700
rect 173600 35700 173700 35800
rect 173600 35800 173700 35900
rect 173600 35900 173700 36000
rect 173600 36000 173700 36100
rect 173600 36100 173700 36200
rect 173600 36200 173700 36300
rect 173600 36300 173700 36400
rect 173600 36400 173700 36500
rect 173600 36500 173700 36600
rect 173600 36600 173700 36700
rect 173600 36700 173700 36800
rect 173600 36800 173700 36900
rect 173600 36900 173700 37000
rect 173600 37000 173700 37100
rect 173600 37100 173700 37200
rect 173600 37200 173700 37300
rect 173600 37300 173700 37400
rect 173600 37400 173700 37500
rect 173600 37500 173700 37600
rect 173700 26500 173800 26600
rect 173700 26600 173800 26700
rect 173700 26700 173800 26800
rect 173700 26800 173800 26900
rect 173700 26900 173800 27000
rect 173700 27000 173800 27100
rect 173700 27100 173800 27200
rect 173700 27200 173800 27300
rect 173700 27300 173800 27400
rect 173700 27400 173800 27500
rect 173700 27500 173800 27600
rect 173700 27600 173800 27700
rect 173700 27700 173800 27800
rect 173700 27800 173800 27900
rect 173700 27900 173800 28000
rect 173700 28000 173800 28100
rect 173700 28100 173800 28200
rect 173700 28200 173800 28300
rect 173700 28300 173800 28400
rect 173700 28400 173800 28500
rect 173700 28500 173800 28600
rect 173700 28600 173800 28700
rect 173700 28700 173800 28800
rect 173700 28800 173800 28900
rect 173700 28900 173800 29000
rect 173700 29000 173800 29100
rect 173700 29100 173800 29200
rect 173700 29200 173800 29300
rect 173700 29300 173800 29400
rect 173700 29400 173800 29500
rect 173700 29500 173800 29600
rect 173700 29600 173800 29700
rect 173700 29700 173800 29800
rect 173700 29800 173800 29900
rect 173700 29900 173800 30000
rect 173700 30000 173800 30100
rect 173700 30100 173800 30200
rect 173700 30200 173800 30300
rect 173700 30300 173800 30400
rect 173700 30400 173800 30500
rect 173700 30500 173800 30600
rect 173700 30600 173800 30700
rect 173700 30700 173800 30800
rect 173700 30800 173800 30900
rect 173700 30900 173800 31000
rect 173700 31000 173800 31100
rect 173700 31100 173800 31200
rect 173700 31200 173800 31300
rect 173700 31300 173800 31400
rect 173700 31400 173800 31500
rect 173700 31500 173800 31600
rect 173700 31600 173800 31700
rect 173700 31700 173800 31800
rect 173700 31800 173800 31900
rect 173700 31900 173800 32000
rect 173700 32000 173800 32100
rect 173700 32100 173800 32200
rect 173700 32200 173800 32300
rect 173700 32300 173800 32400
rect 173700 32400 173800 32500
rect 173700 32500 173800 32600
rect 173700 32600 173800 32700
rect 173700 32700 173800 32800
rect 173700 32800 173800 32900
rect 173700 32900 173800 33000
rect 173700 33000 173800 33100
rect 173700 33100 173800 33200
rect 173700 33200 173800 33300
rect 173700 33300 173800 33400
rect 173700 33400 173800 33500
rect 173700 33500 173800 33600
rect 173700 33600 173800 33700
rect 173700 33700 173800 33800
rect 173700 33800 173800 33900
rect 173700 33900 173800 34000
rect 173700 34000 173800 34100
rect 173700 34100 173800 34200
rect 173700 34200 173800 34300
rect 173700 34300 173800 34400
rect 173700 34400 173800 34500
rect 173700 34500 173800 34600
rect 173700 34600 173800 34700
rect 173700 34700 173800 34800
rect 173700 34800 173800 34900
rect 173700 34900 173800 35000
rect 173700 35000 173800 35100
rect 173700 35100 173800 35200
rect 173700 35200 173800 35300
rect 173700 35300 173800 35400
rect 173700 35400 173800 35500
rect 173700 35500 173800 35600
rect 173700 35600 173800 35700
rect 173700 35700 173800 35800
rect 173700 35800 173800 35900
rect 173700 35900 173800 36000
rect 173700 36000 173800 36100
rect 173700 36100 173800 36200
rect 173700 36200 173800 36300
rect 173700 36300 173800 36400
rect 173700 36400 173800 36500
rect 173700 36500 173800 36600
rect 173700 36600 173800 36700
rect 173700 36700 173800 36800
rect 173700 36800 173800 36900
rect 173700 36900 173800 37000
rect 173700 37000 173800 37100
rect 173700 37100 173800 37200
rect 173700 37200 173800 37300
rect 173700 37300 173800 37400
rect 173700 37400 173800 37500
rect 173800 26000 173900 26100
rect 173800 26100 173900 26200
rect 173800 26200 173900 26300
rect 173800 26300 173900 26400
rect 173800 26400 173900 26500
rect 173800 26500 173900 26600
rect 173800 26600 173900 26700
rect 173800 26700 173900 26800
rect 173800 26800 173900 26900
rect 173800 26900 173900 27000
rect 173800 27000 173900 27100
rect 173800 27100 173900 27200
rect 173800 27200 173900 27300
rect 173800 27300 173900 27400
rect 173800 27400 173900 27500
rect 173800 27500 173900 27600
rect 173800 27600 173900 27700
rect 173800 27700 173900 27800
rect 173800 27800 173900 27900
rect 173800 27900 173900 28000
rect 173800 28000 173900 28100
rect 173800 28100 173900 28200
rect 173800 28200 173900 28300
rect 173800 28300 173900 28400
rect 173800 28400 173900 28500
rect 173800 28500 173900 28600
rect 173800 28600 173900 28700
rect 173800 28700 173900 28800
rect 173800 28800 173900 28900
rect 173800 28900 173900 29000
rect 173800 29000 173900 29100
rect 173800 29100 173900 29200
rect 173800 29200 173900 29300
rect 173800 29300 173900 29400
rect 173800 29400 173900 29500
rect 173800 29500 173900 29600
rect 173800 29600 173900 29700
rect 173800 29700 173900 29800
rect 173800 29800 173900 29900
rect 173800 29900 173900 30000
rect 173800 30000 173900 30100
rect 173800 30100 173900 30200
rect 173800 30200 173900 30300
rect 173800 30300 173900 30400
rect 173800 30400 173900 30500
rect 173800 30500 173900 30600
rect 173800 30600 173900 30700
rect 173800 30700 173900 30800
rect 173800 30800 173900 30900
rect 173800 30900 173900 31000
rect 173800 31000 173900 31100
rect 173800 31100 173900 31200
rect 173800 31200 173900 31300
rect 173800 31300 173900 31400
rect 173800 31400 173900 31500
rect 173800 31500 173900 31600
rect 173800 31600 173900 31700
rect 173800 31700 173900 31800
rect 173800 31800 173900 31900
rect 173800 31900 173900 32000
rect 173800 32000 173900 32100
rect 173800 32100 173900 32200
rect 173800 32200 173900 32300
rect 173800 32300 173900 32400
rect 173800 32400 173900 32500
rect 173800 32500 173900 32600
rect 173800 32600 173900 32700
rect 173800 32700 173900 32800
rect 173800 32800 173900 32900
rect 173800 32900 173900 33000
rect 173800 33000 173900 33100
rect 173800 33100 173900 33200
rect 173800 33200 173900 33300
rect 173800 33300 173900 33400
rect 173800 33400 173900 33500
rect 173800 33500 173900 33600
rect 173800 33600 173900 33700
rect 173800 33700 173900 33800
rect 173800 33800 173900 33900
rect 173800 33900 173900 34000
rect 173800 34000 173900 34100
rect 173800 34100 173900 34200
rect 173800 34200 173900 34300
rect 173800 34300 173900 34400
rect 173800 34400 173900 34500
rect 173800 34500 173900 34600
rect 173800 34600 173900 34700
rect 173800 34700 173900 34800
rect 173800 34800 173900 34900
rect 173800 34900 173900 35000
rect 173800 35000 173900 35100
rect 173800 35100 173900 35200
rect 173800 35200 173900 35300
rect 173800 35300 173900 35400
rect 173800 35400 173900 35500
rect 173800 35500 173900 35600
rect 173800 35600 173900 35700
rect 173800 35700 173900 35800
rect 173800 35800 173900 35900
rect 173800 35900 173900 36000
rect 173800 36000 173900 36100
rect 173800 36100 173900 36200
rect 173800 36200 173900 36300
rect 173800 36300 173900 36400
rect 173800 36400 173900 36500
rect 173800 36500 173900 36600
rect 173800 36600 173900 36700
rect 173800 36700 173900 36800
rect 173800 36800 173900 36900
rect 173800 36900 173900 37000
rect 173800 37000 173900 37100
rect 173800 37100 173900 37200
rect 173800 37200 173900 37300
rect 173900 25400 174000 25500
rect 173900 25500 174000 25600
rect 173900 25600 174000 25700
rect 173900 25700 174000 25800
rect 173900 25800 174000 25900
rect 173900 25900 174000 26000
rect 173900 26000 174000 26100
rect 173900 26100 174000 26200
rect 173900 26200 174000 26300
rect 173900 26300 174000 26400
rect 173900 26400 174000 26500
rect 173900 26500 174000 26600
rect 173900 26600 174000 26700
rect 173900 26700 174000 26800
rect 173900 26800 174000 26900
rect 173900 26900 174000 27000
rect 173900 27000 174000 27100
rect 173900 27100 174000 27200
rect 173900 27200 174000 27300
rect 173900 27300 174000 27400
rect 173900 27400 174000 27500
rect 173900 27500 174000 27600
rect 173900 27600 174000 27700
rect 173900 27700 174000 27800
rect 173900 27800 174000 27900
rect 173900 27900 174000 28000
rect 173900 28000 174000 28100
rect 173900 28100 174000 28200
rect 173900 28200 174000 28300
rect 173900 28300 174000 28400
rect 173900 28400 174000 28500
rect 173900 28500 174000 28600
rect 173900 28600 174000 28700
rect 173900 28700 174000 28800
rect 173900 28800 174000 28900
rect 173900 28900 174000 29000
rect 173900 29000 174000 29100
rect 173900 29100 174000 29200
rect 173900 29200 174000 29300
rect 173900 29300 174000 29400
rect 173900 29400 174000 29500
rect 173900 29500 174000 29600
rect 173900 29600 174000 29700
rect 173900 29700 174000 29800
rect 173900 29800 174000 29900
rect 173900 29900 174000 30000
rect 173900 30000 174000 30100
rect 173900 30100 174000 30200
rect 173900 30200 174000 30300
rect 173900 30300 174000 30400
rect 173900 30400 174000 30500
rect 173900 30500 174000 30600
rect 173900 30600 174000 30700
rect 173900 30700 174000 30800
rect 173900 30800 174000 30900
rect 173900 30900 174000 31000
rect 173900 31000 174000 31100
rect 173900 31100 174000 31200
rect 173900 31200 174000 31300
rect 173900 31300 174000 31400
rect 173900 31400 174000 31500
rect 173900 31500 174000 31600
rect 173900 31600 174000 31700
rect 173900 31700 174000 31800
rect 173900 31800 174000 31900
rect 173900 31900 174000 32000
rect 173900 32000 174000 32100
rect 173900 32100 174000 32200
rect 173900 32200 174000 32300
rect 173900 32300 174000 32400
rect 173900 32400 174000 32500
rect 173900 32500 174000 32600
rect 173900 32600 174000 32700
rect 173900 32700 174000 32800
rect 173900 32800 174000 32900
rect 173900 32900 174000 33000
rect 173900 33000 174000 33100
rect 173900 33100 174000 33200
rect 173900 33200 174000 33300
rect 173900 33300 174000 33400
rect 173900 33400 174000 33500
rect 173900 33500 174000 33600
rect 173900 33600 174000 33700
rect 173900 33700 174000 33800
rect 173900 33800 174000 33900
rect 173900 33900 174000 34000
rect 173900 34000 174000 34100
rect 173900 34100 174000 34200
rect 173900 34200 174000 34300
rect 173900 34300 174000 34400
rect 173900 34400 174000 34500
rect 173900 34500 174000 34600
rect 173900 34600 174000 34700
rect 173900 34700 174000 34800
rect 173900 34800 174000 34900
rect 173900 34900 174000 35000
rect 173900 35000 174000 35100
rect 173900 35100 174000 35200
rect 173900 35200 174000 35300
rect 173900 35300 174000 35400
rect 173900 35400 174000 35500
rect 173900 35500 174000 35600
rect 173900 35600 174000 35700
rect 173900 35700 174000 35800
rect 173900 35800 174000 35900
rect 173900 35900 174000 36000
rect 173900 36000 174000 36100
rect 173900 36100 174000 36200
rect 173900 36200 174000 36300
rect 173900 36300 174000 36400
rect 173900 36400 174000 36500
rect 173900 36500 174000 36600
rect 173900 36600 174000 36700
rect 173900 36700 174000 36800
rect 173900 36800 174000 36900
rect 173900 36900 174000 37000
rect 174000 24900 174100 25000
rect 174000 25000 174100 25100
rect 174000 25100 174100 25200
rect 174000 25200 174100 25300
rect 174000 25300 174100 25400
rect 174000 25400 174100 25500
rect 174000 25500 174100 25600
rect 174000 25600 174100 25700
rect 174000 25700 174100 25800
rect 174000 25800 174100 25900
rect 174000 25900 174100 26000
rect 174000 26000 174100 26100
rect 174000 26100 174100 26200
rect 174000 26200 174100 26300
rect 174000 26300 174100 26400
rect 174000 26400 174100 26500
rect 174000 26500 174100 26600
rect 174000 26600 174100 26700
rect 174000 26700 174100 26800
rect 174000 26800 174100 26900
rect 174000 26900 174100 27000
rect 174000 27000 174100 27100
rect 174000 27100 174100 27200
rect 174000 27200 174100 27300
rect 174000 27300 174100 27400
rect 174000 27400 174100 27500
rect 174000 27500 174100 27600
rect 174000 27600 174100 27700
rect 174000 27700 174100 27800
rect 174000 27800 174100 27900
rect 174000 27900 174100 28000
rect 174000 28000 174100 28100
rect 174000 28100 174100 28200
rect 174000 28200 174100 28300
rect 174000 28300 174100 28400
rect 174000 28400 174100 28500
rect 174000 28500 174100 28600
rect 174000 28600 174100 28700
rect 174000 28700 174100 28800
rect 174000 28800 174100 28900
rect 174000 28900 174100 29000
rect 174000 29000 174100 29100
rect 174000 29100 174100 29200
rect 174000 29200 174100 29300
rect 174000 29300 174100 29400
rect 174000 29400 174100 29500
rect 174000 29500 174100 29600
rect 174000 29600 174100 29700
rect 174000 29700 174100 29800
rect 174000 29800 174100 29900
rect 174000 29900 174100 30000
rect 174000 30000 174100 30100
rect 174000 30100 174100 30200
rect 174000 30200 174100 30300
rect 174000 30300 174100 30400
rect 174000 30400 174100 30500
rect 174000 30500 174100 30600
rect 174000 30600 174100 30700
rect 174000 30700 174100 30800
rect 174000 30800 174100 30900
rect 174000 30900 174100 31000
rect 174000 31000 174100 31100
rect 174000 31100 174100 31200
rect 174000 31200 174100 31300
rect 174000 31300 174100 31400
rect 174000 31400 174100 31500
rect 174000 31500 174100 31600
rect 174000 31600 174100 31700
rect 174000 31700 174100 31800
rect 174000 31800 174100 31900
rect 174000 31900 174100 32000
rect 174000 32000 174100 32100
rect 174000 32100 174100 32200
rect 174000 32200 174100 32300
rect 174000 32300 174100 32400
rect 174000 32400 174100 32500
rect 174000 32500 174100 32600
rect 174000 32600 174100 32700
rect 174000 32700 174100 32800
rect 174000 32800 174100 32900
rect 174000 32900 174100 33000
rect 174000 33000 174100 33100
rect 174000 33100 174100 33200
rect 174000 33200 174100 33300
rect 174000 33300 174100 33400
rect 174000 33400 174100 33500
rect 174000 33500 174100 33600
rect 174000 33600 174100 33700
rect 174000 33700 174100 33800
rect 174000 33800 174100 33900
rect 174000 33900 174100 34000
rect 174000 34000 174100 34100
rect 174000 34100 174100 34200
rect 174000 34200 174100 34300
rect 174000 34300 174100 34400
rect 174000 34400 174100 34500
rect 174000 34500 174100 34600
rect 174000 34600 174100 34700
rect 174000 34700 174100 34800
rect 174000 34800 174100 34900
rect 174000 34900 174100 35000
rect 174000 35000 174100 35100
rect 174000 35100 174100 35200
rect 174000 35200 174100 35300
rect 174000 35300 174100 35400
rect 174000 35400 174100 35500
rect 174000 35500 174100 35600
rect 174000 35600 174100 35700
rect 174000 35700 174100 35800
rect 174000 35800 174100 35900
rect 174000 35900 174100 36000
rect 174000 36000 174100 36100
rect 174000 36100 174100 36200
rect 174000 36200 174100 36300
rect 174000 36300 174100 36400
rect 174000 36400 174100 36500
rect 174000 36500 174100 36600
rect 174000 36600 174100 36700
rect 174100 24300 174200 24400
rect 174100 24400 174200 24500
rect 174100 24500 174200 24600
rect 174100 24600 174200 24700
rect 174100 24700 174200 24800
rect 174100 24800 174200 24900
rect 174100 24900 174200 25000
rect 174100 25000 174200 25100
rect 174100 25100 174200 25200
rect 174100 25200 174200 25300
rect 174100 25300 174200 25400
rect 174100 25400 174200 25500
rect 174100 25500 174200 25600
rect 174100 25600 174200 25700
rect 174100 25700 174200 25800
rect 174100 25800 174200 25900
rect 174100 25900 174200 26000
rect 174100 26000 174200 26100
rect 174100 26100 174200 26200
rect 174100 26200 174200 26300
rect 174100 26300 174200 26400
rect 174100 26400 174200 26500
rect 174100 26500 174200 26600
rect 174100 26600 174200 26700
rect 174100 26700 174200 26800
rect 174100 26800 174200 26900
rect 174100 26900 174200 27000
rect 174100 27000 174200 27100
rect 174100 27100 174200 27200
rect 174100 27200 174200 27300
rect 174100 27300 174200 27400
rect 174100 27400 174200 27500
rect 174100 27500 174200 27600
rect 174100 27600 174200 27700
rect 174100 27700 174200 27800
rect 174100 27800 174200 27900
rect 174100 27900 174200 28000
rect 174100 28000 174200 28100
rect 174100 28100 174200 28200
rect 174100 28200 174200 28300
rect 174100 28300 174200 28400
rect 174100 28400 174200 28500
rect 174100 28500 174200 28600
rect 174100 28600 174200 28700
rect 174100 28700 174200 28800
rect 174100 28800 174200 28900
rect 174100 28900 174200 29000
rect 174100 29000 174200 29100
rect 174100 29100 174200 29200
rect 174100 29200 174200 29300
rect 174100 29300 174200 29400
rect 174100 29400 174200 29500
rect 174100 29500 174200 29600
rect 174100 29600 174200 29700
rect 174100 29700 174200 29800
rect 174100 29800 174200 29900
rect 174100 29900 174200 30000
rect 174100 30000 174200 30100
rect 174100 30100 174200 30200
rect 174100 30200 174200 30300
rect 174100 30300 174200 30400
rect 174100 30400 174200 30500
rect 174100 30500 174200 30600
rect 174100 30600 174200 30700
rect 174100 30700 174200 30800
rect 174100 30800 174200 30900
rect 174100 30900 174200 31000
rect 174100 31000 174200 31100
rect 174100 31100 174200 31200
rect 174100 31200 174200 31300
rect 174100 31300 174200 31400
rect 174100 31400 174200 31500
rect 174100 31500 174200 31600
rect 174100 31600 174200 31700
rect 174100 31700 174200 31800
rect 174100 31800 174200 31900
rect 174100 31900 174200 32000
rect 174100 32000 174200 32100
rect 174100 32100 174200 32200
rect 174100 32200 174200 32300
rect 174100 32300 174200 32400
rect 174100 32400 174200 32500
rect 174100 32500 174200 32600
rect 174100 32600 174200 32700
rect 174100 32700 174200 32800
rect 174100 32800 174200 32900
rect 174100 32900 174200 33000
rect 174100 33000 174200 33100
rect 174100 33100 174200 33200
rect 174100 33200 174200 33300
rect 174100 33300 174200 33400
rect 174100 33400 174200 33500
rect 174100 33500 174200 33600
rect 174100 33600 174200 33700
rect 174100 33700 174200 33800
rect 174100 33800 174200 33900
rect 174100 33900 174200 34000
rect 174100 34000 174200 34100
rect 174100 34100 174200 34200
rect 174100 34200 174200 34300
rect 174100 34300 174200 34400
rect 174100 34400 174200 34500
rect 174100 34500 174200 34600
rect 174100 34600 174200 34700
rect 174100 34700 174200 34800
rect 174100 34800 174200 34900
rect 174100 34900 174200 35000
rect 174100 35000 174200 35100
rect 174100 35100 174200 35200
rect 174100 35200 174200 35300
rect 174100 35300 174200 35400
rect 174100 35400 174200 35500
rect 174100 35500 174200 35600
rect 174100 35600 174200 35700
rect 174100 35700 174200 35800
rect 174100 35800 174200 35900
rect 174100 35900 174200 36000
rect 174100 36000 174200 36100
rect 174100 36100 174200 36200
rect 174200 23800 174300 23900
rect 174200 23900 174300 24000
rect 174200 24000 174300 24100
rect 174200 24100 174300 24200
rect 174200 24200 174300 24300
rect 174200 24300 174300 24400
rect 174200 24400 174300 24500
rect 174200 24500 174300 24600
rect 174200 24600 174300 24700
rect 174200 24700 174300 24800
rect 174200 24800 174300 24900
rect 174200 24900 174300 25000
rect 174200 25000 174300 25100
rect 174200 25100 174300 25200
rect 174200 25200 174300 25300
rect 174200 25300 174300 25400
rect 174200 25400 174300 25500
rect 174200 25500 174300 25600
rect 174200 25600 174300 25700
rect 174200 25700 174300 25800
rect 174200 25800 174300 25900
rect 174200 25900 174300 26000
rect 174200 26000 174300 26100
rect 174200 26100 174300 26200
rect 174200 26200 174300 26300
rect 174200 26300 174300 26400
rect 174200 26400 174300 26500
rect 174200 26500 174300 26600
rect 174200 26600 174300 26700
rect 174200 26700 174300 26800
rect 174200 26800 174300 26900
rect 174200 26900 174300 27000
rect 174200 27000 174300 27100
rect 174200 27100 174300 27200
rect 174200 27200 174300 27300
rect 174200 27300 174300 27400
rect 174200 27400 174300 27500
rect 174200 27500 174300 27600
rect 174200 27600 174300 27700
rect 174200 27700 174300 27800
rect 174200 27800 174300 27900
rect 174200 27900 174300 28000
rect 174200 28000 174300 28100
rect 174200 28100 174300 28200
rect 174200 28200 174300 28300
rect 174200 28300 174300 28400
rect 174200 28400 174300 28500
rect 174200 28500 174300 28600
rect 174200 28600 174300 28700
rect 174200 28700 174300 28800
rect 174200 28800 174300 28900
rect 174200 28900 174300 29000
rect 174200 29000 174300 29100
rect 174200 29100 174300 29200
rect 174200 29200 174300 29300
rect 174200 29300 174300 29400
rect 174200 29400 174300 29500
rect 174200 29500 174300 29600
rect 174200 29600 174300 29700
rect 174200 29700 174300 29800
rect 174200 29800 174300 29900
rect 174200 29900 174300 30000
rect 174200 30000 174300 30100
rect 174200 30100 174300 30200
rect 174200 30200 174300 30300
rect 174200 30300 174300 30400
rect 174200 30400 174300 30500
rect 174200 30500 174300 30600
rect 174200 30600 174300 30700
rect 174200 30700 174300 30800
rect 174200 30800 174300 30900
rect 174200 30900 174300 31000
rect 174200 31000 174300 31100
rect 174200 31100 174300 31200
rect 174200 31200 174300 31300
rect 174200 31300 174300 31400
rect 174200 31400 174300 31500
rect 174200 31500 174300 31600
rect 174200 31600 174300 31700
rect 174200 31700 174300 31800
rect 174200 31800 174300 31900
rect 174200 31900 174300 32000
rect 174200 32000 174300 32100
rect 174200 32100 174300 32200
rect 174200 32200 174300 32300
rect 174200 32300 174300 32400
rect 174200 32400 174300 32500
rect 174200 32500 174300 32600
rect 174200 32600 174300 32700
rect 174200 32700 174300 32800
rect 174200 32800 174300 32900
rect 174200 32900 174300 33000
rect 174200 33000 174300 33100
rect 174200 33100 174300 33200
rect 174200 33200 174300 33300
rect 174200 33300 174300 33400
rect 174200 33400 174300 33500
rect 174200 33500 174300 33600
rect 174200 33600 174300 33700
rect 174200 33700 174300 33800
rect 174200 33800 174300 33900
rect 174200 33900 174300 34000
rect 174200 34000 174300 34100
rect 174200 34100 174300 34200
rect 174200 34200 174300 34300
rect 174200 34300 174300 34400
rect 174200 34400 174300 34500
rect 174200 34500 174300 34600
rect 174200 34600 174300 34700
rect 174200 34700 174300 34800
rect 174200 34800 174300 34900
rect 174200 34900 174300 35000
rect 174200 35000 174300 35100
rect 174200 35100 174300 35200
rect 174200 35200 174300 35300
rect 174200 35300 174300 35400
rect 174200 35400 174300 35500
rect 174200 35500 174300 35600
rect 174200 35600 174300 35700
rect 174300 23500 174400 23600
rect 174300 23600 174400 23700
rect 174300 23700 174400 23800
rect 174300 23800 174400 23900
rect 174300 23900 174400 24000
rect 174300 24000 174400 24100
rect 174300 24100 174400 24200
rect 174300 24200 174400 24300
rect 174300 24300 174400 24400
rect 174300 24400 174400 24500
rect 174300 24500 174400 24600
rect 174300 24600 174400 24700
rect 174300 24700 174400 24800
rect 174300 24800 174400 24900
rect 174300 24900 174400 25000
rect 174300 25000 174400 25100
rect 174300 25100 174400 25200
rect 174300 25200 174400 25300
rect 174300 25300 174400 25400
rect 174300 25400 174400 25500
rect 174300 25500 174400 25600
rect 174300 25600 174400 25700
rect 174300 25700 174400 25800
rect 174300 25800 174400 25900
rect 174300 25900 174400 26000
rect 174300 26000 174400 26100
rect 174300 26100 174400 26200
rect 174300 26200 174400 26300
rect 174300 26300 174400 26400
rect 174300 26400 174400 26500
rect 174300 26500 174400 26600
rect 174300 26600 174400 26700
rect 174300 26700 174400 26800
rect 174300 26800 174400 26900
rect 174300 26900 174400 27000
rect 174300 27000 174400 27100
rect 174300 27100 174400 27200
rect 174300 27200 174400 27300
rect 174300 27300 174400 27400
rect 174300 27400 174400 27500
rect 174300 27500 174400 27600
rect 174300 27600 174400 27700
rect 174300 27700 174400 27800
rect 174300 27800 174400 27900
rect 174300 27900 174400 28000
rect 174300 28000 174400 28100
rect 174300 28100 174400 28200
rect 174300 28200 174400 28300
rect 174300 28300 174400 28400
rect 174300 28400 174400 28500
rect 174300 28500 174400 28600
rect 174300 28600 174400 28700
rect 174300 28700 174400 28800
rect 174300 28800 174400 28900
rect 174300 28900 174400 29000
rect 174300 29000 174400 29100
rect 174300 29100 174400 29200
rect 174300 29200 174400 29300
rect 174300 29300 174400 29400
rect 174300 29400 174400 29500
rect 174300 29500 174400 29600
rect 174300 29600 174400 29700
rect 174300 29700 174400 29800
rect 174300 29800 174400 29900
rect 174300 29900 174400 30000
rect 174300 30000 174400 30100
rect 174300 30100 174400 30200
rect 174300 30200 174400 30300
rect 174300 30300 174400 30400
rect 174300 30400 174400 30500
rect 174300 30500 174400 30600
rect 174300 30600 174400 30700
rect 174300 30700 174400 30800
rect 174300 30800 174400 30900
rect 174300 30900 174400 31000
rect 174300 31000 174400 31100
rect 174300 31100 174400 31200
rect 174300 31200 174400 31300
rect 174300 31300 174400 31400
rect 174300 31400 174400 31500
rect 174300 31500 174400 31600
rect 174300 31600 174400 31700
rect 174300 31700 174400 31800
rect 174300 31800 174400 31900
rect 174300 31900 174400 32000
rect 174300 32000 174400 32100
rect 174300 32100 174400 32200
rect 174300 32200 174400 32300
rect 174300 32300 174400 32400
rect 174300 32400 174400 32500
rect 174300 32500 174400 32600
rect 174300 32600 174400 32700
rect 174300 32700 174400 32800
rect 174300 32800 174400 32900
rect 174300 32900 174400 33000
rect 174300 33000 174400 33100
rect 174300 33100 174400 33200
rect 174300 33200 174400 33300
rect 174300 33300 174400 33400
rect 174300 33400 174400 33500
rect 174300 33500 174400 33600
rect 174300 33600 174400 33700
rect 174300 33700 174400 33800
rect 174300 33800 174400 33900
rect 174300 33900 174400 34000
rect 174300 34000 174400 34100
rect 174300 34100 174400 34200
rect 174300 34200 174400 34300
rect 174300 34300 174400 34400
rect 174300 34400 174400 34500
rect 174300 34500 174400 34600
rect 174300 34600 174400 34700
rect 174300 34700 174400 34800
rect 174300 34800 174400 34900
rect 174300 34900 174400 35000
rect 174300 35000 174400 35100
rect 174400 23200 174500 23300
rect 174400 23300 174500 23400
rect 174400 23400 174500 23500
rect 174400 23500 174500 23600
rect 174400 23600 174500 23700
rect 174400 23700 174500 23800
rect 174400 23800 174500 23900
rect 174400 23900 174500 24000
rect 174400 24000 174500 24100
rect 174400 24100 174500 24200
rect 174400 24200 174500 24300
rect 174400 24300 174500 24400
rect 174400 24400 174500 24500
rect 174400 24500 174500 24600
rect 174400 24600 174500 24700
rect 174400 24700 174500 24800
rect 174400 24800 174500 24900
rect 174400 24900 174500 25000
rect 174400 25000 174500 25100
rect 174400 25100 174500 25200
rect 174400 25200 174500 25300
rect 174400 25300 174500 25400
rect 174400 25400 174500 25500
rect 174400 25500 174500 25600
rect 174400 25600 174500 25700
rect 174400 25700 174500 25800
rect 174400 25800 174500 25900
rect 174400 25900 174500 26000
rect 174400 26000 174500 26100
rect 174400 26100 174500 26200
rect 174400 26200 174500 26300
rect 174400 26300 174500 26400
rect 174400 26400 174500 26500
rect 174400 26500 174500 26600
rect 174400 26600 174500 26700
rect 174400 26700 174500 26800
rect 174400 26800 174500 26900
rect 174400 26900 174500 27000
rect 174400 27000 174500 27100
rect 174400 27100 174500 27200
rect 174400 27200 174500 27300
rect 174400 27300 174500 27400
rect 174400 27400 174500 27500
rect 174400 27500 174500 27600
rect 174400 27600 174500 27700
rect 174400 27700 174500 27800
rect 174400 27800 174500 27900
rect 174400 27900 174500 28000
rect 174400 28000 174500 28100
rect 174400 28100 174500 28200
rect 174400 28200 174500 28300
rect 174400 28300 174500 28400
rect 174400 28400 174500 28500
rect 174400 28500 174500 28600
rect 174400 28600 174500 28700
rect 174400 28700 174500 28800
rect 174400 28800 174500 28900
rect 174400 28900 174500 29000
rect 174400 29000 174500 29100
rect 174400 29100 174500 29200
rect 174400 29200 174500 29300
rect 174400 29300 174500 29400
rect 174400 29400 174500 29500
rect 174400 29500 174500 29600
rect 174400 29600 174500 29700
rect 174400 29700 174500 29800
rect 174400 29800 174500 29900
rect 174400 29900 174500 30000
rect 174400 30000 174500 30100
rect 174400 30100 174500 30200
rect 174400 30200 174500 30300
rect 174400 30300 174500 30400
rect 174400 30400 174500 30500
rect 174400 30500 174500 30600
rect 174400 30600 174500 30700
rect 174400 30700 174500 30800
rect 174400 30800 174500 30900
rect 174400 30900 174500 31000
rect 174400 31000 174500 31100
rect 174400 31100 174500 31200
rect 174400 31200 174500 31300
rect 174400 31300 174500 31400
rect 174400 31400 174500 31500
rect 174400 31500 174500 31600
rect 174400 31600 174500 31700
rect 174400 31700 174500 31800
rect 174400 31800 174500 31900
rect 174400 31900 174500 32000
rect 174400 32000 174500 32100
rect 174400 32100 174500 32200
rect 174400 32200 174500 32300
rect 174400 32300 174500 32400
rect 174400 32400 174500 32500
rect 174400 32500 174500 32600
rect 174400 32600 174500 32700
rect 174400 32700 174500 32800
rect 174400 32800 174500 32900
rect 174400 32900 174500 33000
rect 174400 33000 174500 33100
rect 174400 33100 174500 33200
rect 174400 33200 174500 33300
rect 174400 33300 174500 33400
rect 174400 33400 174500 33500
rect 174400 33500 174500 33600
rect 174400 33600 174500 33700
rect 174400 33700 174500 33800
rect 174400 33800 174500 33900
rect 174400 33900 174500 34000
rect 174400 34000 174500 34100
rect 174400 34100 174500 34200
rect 174400 34200 174500 34300
rect 174400 34300 174500 34400
rect 174500 22900 174600 23000
rect 174500 23000 174600 23100
rect 174500 23100 174600 23200
rect 174500 23200 174600 23300
rect 174500 23300 174600 23400
rect 174500 23400 174600 23500
rect 174500 23500 174600 23600
rect 174500 23600 174600 23700
rect 174500 23700 174600 23800
rect 174500 23800 174600 23900
rect 174500 23900 174600 24000
rect 174500 24000 174600 24100
rect 174500 24100 174600 24200
rect 174500 24200 174600 24300
rect 174500 24300 174600 24400
rect 174500 24400 174600 24500
rect 174500 24500 174600 24600
rect 174500 24600 174600 24700
rect 174500 24700 174600 24800
rect 174500 24800 174600 24900
rect 174500 24900 174600 25000
rect 174500 25000 174600 25100
rect 174500 25100 174600 25200
rect 174500 25200 174600 25300
rect 174500 25300 174600 25400
rect 174500 25400 174600 25500
rect 174500 25500 174600 25600
rect 174500 25600 174600 25700
rect 174500 25700 174600 25800
rect 174500 25800 174600 25900
rect 174500 25900 174600 26000
rect 174500 26000 174600 26100
rect 174500 26100 174600 26200
rect 174500 26200 174600 26300
rect 174500 26300 174600 26400
rect 174500 26400 174600 26500
rect 174500 26500 174600 26600
rect 174500 26600 174600 26700
rect 174500 26700 174600 26800
rect 174500 26800 174600 26900
rect 174500 26900 174600 27000
rect 174500 27000 174600 27100
rect 174500 27100 174600 27200
rect 174500 27200 174600 27300
rect 174500 27300 174600 27400
rect 174500 27400 174600 27500
rect 174500 27500 174600 27600
rect 174500 27600 174600 27700
rect 174500 27700 174600 27800
rect 174500 27800 174600 27900
rect 174500 27900 174600 28000
rect 174500 28000 174600 28100
rect 174500 28100 174600 28200
rect 174500 28200 174600 28300
rect 174500 28300 174600 28400
rect 174500 28400 174600 28500
rect 174500 28500 174600 28600
rect 174500 28600 174600 28700
rect 174500 28700 174600 28800
rect 174500 28800 174600 28900
rect 174500 28900 174600 29000
rect 174500 29000 174600 29100
rect 174500 29100 174600 29200
rect 174500 29200 174600 29300
rect 174500 29300 174600 29400
rect 174500 29400 174600 29500
rect 174500 29500 174600 29600
rect 174500 29600 174600 29700
rect 174500 29700 174600 29800
rect 174500 29800 174600 29900
rect 174500 29900 174600 30000
rect 174500 30000 174600 30100
rect 174500 30100 174600 30200
rect 174500 30200 174600 30300
rect 174500 30300 174600 30400
rect 174500 30400 174600 30500
rect 174500 30500 174600 30600
rect 174500 30600 174600 30700
rect 174500 30700 174600 30800
rect 174500 30800 174600 30900
rect 174500 30900 174600 31000
rect 174500 31000 174600 31100
rect 174500 31100 174600 31200
rect 174500 31200 174600 31300
rect 174500 31300 174600 31400
rect 174500 31400 174600 31500
rect 174500 31500 174600 31600
rect 174500 31600 174600 31700
rect 174500 31700 174600 31800
rect 174500 31800 174600 31900
rect 174500 31900 174600 32000
rect 174500 32000 174600 32100
rect 174500 32100 174600 32200
rect 174500 32200 174600 32300
rect 174500 32300 174600 32400
rect 174500 32400 174600 32500
rect 174500 32500 174600 32600
rect 174500 32600 174600 32700
rect 174500 32700 174600 32800
rect 174500 32800 174600 32900
rect 174500 32900 174600 33000
rect 174500 33000 174600 33100
rect 174500 33100 174600 33200
rect 174500 33200 174600 33300
rect 174500 33300 174600 33400
rect 174500 33400 174600 33500
rect 174500 33500 174600 33600
rect 174600 22600 174700 22700
rect 174600 22700 174700 22800
rect 174600 22800 174700 22900
rect 174600 22900 174700 23000
rect 174600 23000 174700 23100
rect 174600 23100 174700 23200
rect 174600 23200 174700 23300
rect 174600 23300 174700 23400
rect 174600 23400 174700 23500
rect 174600 23500 174700 23600
rect 174600 23600 174700 23700
rect 174600 23700 174700 23800
rect 174600 23800 174700 23900
rect 174600 23900 174700 24000
rect 174600 24000 174700 24100
rect 174600 24100 174700 24200
rect 174600 24200 174700 24300
rect 174600 24300 174700 24400
rect 174600 24400 174700 24500
rect 174600 24500 174700 24600
rect 174600 24600 174700 24700
rect 174600 24700 174700 24800
rect 174600 24800 174700 24900
rect 174600 24900 174700 25000
rect 174600 25000 174700 25100
rect 174600 25100 174700 25200
rect 174600 25200 174700 25300
rect 174600 25300 174700 25400
rect 174600 25400 174700 25500
rect 174600 25500 174700 25600
rect 174600 25600 174700 25700
rect 174600 25700 174700 25800
rect 174600 25800 174700 25900
rect 174600 25900 174700 26000
rect 174600 26000 174700 26100
rect 174600 26100 174700 26200
rect 174600 26200 174700 26300
rect 174600 26300 174700 26400
rect 174600 26400 174700 26500
rect 174600 26500 174700 26600
rect 174600 26600 174700 26700
rect 174600 26700 174700 26800
rect 174600 26800 174700 26900
rect 174600 26900 174700 27000
rect 174600 27000 174700 27100
rect 174600 27100 174700 27200
rect 174600 27200 174700 27300
rect 174600 27300 174700 27400
rect 174600 27400 174700 27500
rect 174600 27500 174700 27600
rect 174600 27600 174700 27700
rect 174600 27700 174700 27800
rect 174600 27800 174700 27900
rect 174600 27900 174700 28000
rect 174600 28000 174700 28100
rect 174600 28100 174700 28200
rect 174600 28200 174700 28300
rect 174600 28300 174700 28400
rect 174600 28400 174700 28500
rect 174600 28500 174700 28600
rect 174600 28600 174700 28700
rect 174600 28700 174700 28800
rect 174600 28800 174700 28900
rect 174600 28900 174700 29000
rect 174600 29000 174700 29100
rect 174600 29100 174700 29200
rect 174600 29200 174700 29300
rect 174600 29300 174700 29400
rect 174600 29400 174700 29500
rect 174600 29500 174700 29600
rect 174600 29600 174700 29700
rect 174600 29700 174700 29800
rect 174600 29800 174700 29900
rect 174600 29900 174700 30000
rect 174600 30000 174700 30100
rect 174600 30100 174700 30200
rect 174600 30200 174700 30300
rect 174600 30300 174700 30400
rect 174600 30400 174700 30500
rect 174600 30500 174700 30600
rect 174600 30600 174700 30700
rect 174600 30700 174700 30800
rect 174600 30800 174700 30900
rect 174600 30900 174700 31000
rect 174600 31000 174700 31100
rect 174600 31100 174700 31200
rect 174600 31200 174700 31300
rect 174600 31300 174700 31400
rect 174600 31400 174700 31500
rect 174600 31500 174700 31600
rect 174600 31600 174700 31700
rect 174600 31700 174700 31800
rect 174600 31800 174700 31900
rect 174600 31900 174700 32000
rect 174600 32000 174700 32100
rect 174600 32100 174700 32200
rect 174600 32200 174700 32300
rect 174600 32300 174700 32400
rect 174600 32400 174700 32500
rect 174600 32500 174700 32600
rect 174600 32600 174700 32700
rect 174600 32700 174700 32800
rect 174700 22200 174800 22300
rect 174700 22300 174800 22400
rect 174700 22400 174800 22500
rect 174700 22500 174800 22600
rect 174700 22600 174800 22700
rect 174700 22700 174800 22800
rect 174700 22800 174800 22900
rect 174700 22900 174800 23000
rect 174700 23000 174800 23100
rect 174700 23100 174800 23200
rect 174700 23200 174800 23300
rect 174700 23300 174800 23400
rect 174700 23400 174800 23500
rect 174700 23500 174800 23600
rect 174700 23600 174800 23700
rect 174700 23700 174800 23800
rect 174700 23800 174800 23900
rect 174700 23900 174800 24000
rect 174700 24000 174800 24100
rect 174700 24100 174800 24200
rect 174700 24200 174800 24300
rect 174700 24300 174800 24400
rect 174700 24400 174800 24500
rect 174700 24500 174800 24600
rect 174700 24600 174800 24700
rect 174700 24700 174800 24800
rect 174700 24800 174800 24900
rect 174700 24900 174800 25000
rect 174700 25000 174800 25100
rect 174700 25100 174800 25200
rect 174700 25200 174800 25300
rect 174700 25300 174800 25400
rect 174700 25400 174800 25500
rect 174700 25500 174800 25600
rect 174700 25600 174800 25700
rect 174700 25700 174800 25800
rect 174700 25800 174800 25900
rect 174700 25900 174800 26000
rect 174700 26000 174800 26100
rect 174700 26100 174800 26200
rect 174700 26200 174800 26300
rect 174700 26300 174800 26400
rect 174700 26400 174800 26500
rect 174700 26500 174800 26600
rect 174700 26600 174800 26700
rect 174700 26700 174800 26800
rect 174700 26800 174800 26900
rect 174700 26900 174800 27000
rect 174700 27000 174800 27100
rect 174700 27100 174800 27200
rect 174700 27200 174800 27300
rect 174700 27300 174800 27400
rect 174700 27400 174800 27500
rect 174700 27500 174800 27600
rect 174700 27600 174800 27700
rect 174700 27700 174800 27800
rect 174700 27800 174800 27900
rect 174700 27900 174800 28000
rect 174700 28000 174800 28100
rect 174700 28100 174800 28200
rect 174700 28200 174800 28300
rect 174700 28300 174800 28400
rect 174700 28400 174800 28500
rect 174700 28500 174800 28600
rect 174700 28600 174800 28700
rect 174700 28700 174800 28800
rect 174700 28800 174800 28900
rect 174700 28900 174800 29000
rect 174700 29000 174800 29100
rect 174700 29100 174800 29200
rect 174700 29200 174800 29300
rect 174700 29300 174800 29400
rect 174700 29400 174800 29500
rect 174700 29500 174800 29600
rect 174700 29600 174800 29700
rect 174700 29700 174800 29800
rect 174700 29800 174800 29900
rect 174700 29900 174800 30000
rect 174700 30000 174800 30100
rect 174700 30100 174800 30200
rect 174700 30200 174800 30300
rect 174700 30300 174800 30400
rect 174700 30400 174800 30500
rect 174700 30500 174800 30600
rect 174700 30600 174800 30700
rect 174700 30700 174800 30800
rect 174700 30800 174800 30900
rect 174700 30900 174800 31000
rect 174700 31000 174800 31100
rect 174700 31100 174800 31200
rect 174700 31200 174800 31300
rect 174700 31300 174800 31400
rect 174700 31400 174800 31500
rect 174700 31500 174800 31600
rect 174700 31600 174800 31700
rect 174700 31700 174800 31800
rect 174700 31800 174800 31900
rect 174700 31900 174800 32000
rect 174700 32000 174800 32100
rect 174800 21900 174900 22000
rect 174800 22000 174900 22100
rect 174800 22100 174900 22200
rect 174800 22200 174900 22300
rect 174800 22300 174900 22400
rect 174800 22400 174900 22500
rect 174800 22500 174900 22600
rect 174800 22600 174900 22700
rect 174800 22700 174900 22800
rect 174800 22800 174900 22900
rect 174800 22900 174900 23000
rect 174800 23000 174900 23100
rect 174800 23100 174900 23200
rect 174800 23200 174900 23300
rect 174800 23300 174900 23400
rect 174800 23400 174900 23500
rect 174800 23500 174900 23600
rect 174800 23600 174900 23700
rect 174800 23700 174900 23800
rect 174800 23800 174900 23900
rect 174800 23900 174900 24000
rect 174800 24000 174900 24100
rect 174800 24100 174900 24200
rect 174800 24200 174900 24300
rect 174800 24300 174900 24400
rect 174800 24400 174900 24500
rect 174800 24500 174900 24600
rect 174800 24600 174900 24700
rect 174800 24700 174900 24800
rect 174800 24800 174900 24900
rect 174800 24900 174900 25000
rect 174800 25000 174900 25100
rect 174800 25100 174900 25200
rect 174800 25200 174900 25300
rect 174800 25300 174900 25400
rect 174800 25400 174900 25500
rect 174800 25500 174900 25600
rect 174800 25600 174900 25700
rect 174800 25700 174900 25800
rect 174800 25800 174900 25900
rect 174800 25900 174900 26000
rect 174800 26000 174900 26100
rect 174800 26100 174900 26200
rect 174800 26200 174900 26300
rect 174800 26300 174900 26400
rect 174800 26400 174900 26500
rect 174800 26500 174900 26600
rect 174800 26600 174900 26700
rect 174800 26700 174900 26800
rect 174800 26800 174900 26900
rect 174800 26900 174900 27000
rect 174800 27000 174900 27100
rect 174800 27100 174900 27200
rect 174800 27200 174900 27300
rect 174800 27300 174900 27400
rect 174800 27400 174900 27500
rect 174800 27500 174900 27600
rect 174800 27600 174900 27700
rect 174800 27700 174900 27800
rect 174800 27800 174900 27900
rect 174800 27900 174900 28000
rect 174800 28000 174900 28100
rect 174800 28100 174900 28200
rect 174800 28200 174900 28300
rect 174800 28300 174900 28400
rect 174800 28400 174900 28500
rect 174800 28500 174900 28600
rect 174800 28600 174900 28700
rect 174800 28700 174900 28800
rect 174800 28800 174900 28900
rect 174800 28900 174900 29000
rect 174800 29000 174900 29100
rect 174800 29100 174900 29200
rect 174800 29200 174900 29300
rect 174800 29300 174900 29400
rect 174800 29400 174900 29500
rect 174800 29500 174900 29600
rect 174800 29600 174900 29700
rect 174800 29700 174900 29800
rect 174800 29800 174900 29900
rect 174800 29900 174900 30000
rect 174800 30000 174900 30100
rect 174800 30100 174900 30200
rect 174800 30200 174900 30300
rect 174800 30300 174900 30400
rect 174800 30400 174900 30500
rect 174800 30500 174900 30600
rect 174800 30600 174900 30700
rect 174800 30700 174900 30800
rect 174800 30800 174900 30900
rect 174800 30900 174900 31000
rect 174800 31000 174900 31100
rect 174800 31100 174900 31200
rect 174800 31200 174900 31300
rect 174800 31300 174900 31400
rect 174800 31400 174900 31500
rect 174900 21800 175000 21900
rect 174900 21900 175000 22000
rect 174900 22000 175000 22100
rect 174900 22100 175000 22200
rect 174900 22200 175000 22300
rect 174900 22300 175000 22400
rect 174900 22400 175000 22500
rect 174900 22500 175000 22600
rect 174900 22600 175000 22700
rect 174900 22700 175000 22800
rect 174900 22800 175000 22900
rect 174900 22900 175000 23000
rect 174900 23000 175000 23100
rect 174900 23100 175000 23200
rect 174900 23200 175000 23300
rect 174900 23300 175000 23400
rect 174900 23400 175000 23500
rect 174900 23500 175000 23600
rect 174900 23600 175000 23700
rect 174900 23700 175000 23800
rect 174900 23800 175000 23900
rect 174900 23900 175000 24000
rect 174900 24000 175000 24100
rect 174900 24100 175000 24200
rect 174900 24200 175000 24300
rect 174900 24300 175000 24400
rect 174900 24400 175000 24500
rect 174900 24500 175000 24600
rect 174900 24600 175000 24700
rect 174900 24700 175000 24800
rect 174900 24800 175000 24900
rect 174900 24900 175000 25000
rect 174900 25000 175000 25100
rect 174900 25100 175000 25200
rect 174900 25200 175000 25300
rect 174900 25300 175000 25400
rect 174900 25400 175000 25500
rect 174900 25500 175000 25600
rect 174900 25600 175000 25700
rect 174900 25700 175000 25800
rect 174900 25800 175000 25900
rect 174900 25900 175000 26000
rect 174900 26000 175000 26100
rect 174900 26100 175000 26200
rect 174900 26200 175000 26300
rect 174900 26300 175000 26400
rect 174900 26400 175000 26500
rect 174900 26500 175000 26600
rect 174900 26600 175000 26700
rect 174900 26700 175000 26800
rect 174900 26800 175000 26900
rect 174900 26900 175000 27000
rect 174900 27000 175000 27100
rect 174900 27100 175000 27200
rect 174900 27200 175000 27300
rect 174900 27300 175000 27400
rect 174900 27400 175000 27500
rect 174900 27500 175000 27600
rect 174900 27600 175000 27700
rect 174900 27700 175000 27800
rect 174900 27800 175000 27900
rect 174900 27900 175000 28000
rect 174900 28000 175000 28100
rect 174900 28100 175000 28200
rect 174900 28200 175000 28300
rect 174900 28300 175000 28400
rect 174900 28400 175000 28500
rect 174900 28500 175000 28600
rect 174900 28600 175000 28700
rect 174900 28700 175000 28800
rect 174900 28800 175000 28900
rect 174900 28900 175000 29000
rect 174900 29000 175000 29100
rect 174900 29100 175000 29200
rect 174900 29200 175000 29300
rect 174900 29300 175000 29400
rect 174900 29400 175000 29500
rect 174900 29500 175000 29600
rect 174900 29600 175000 29700
rect 174900 29700 175000 29800
rect 174900 29800 175000 29900
rect 174900 29900 175000 30000
rect 174900 30000 175000 30100
rect 174900 30100 175000 30200
rect 174900 30200 175000 30300
rect 174900 30300 175000 30400
rect 174900 30400 175000 30500
rect 174900 30500 175000 30600
rect 174900 30600 175000 30700
rect 174900 30700 175000 30800
rect 174900 30800 175000 30900
rect 175000 21700 175100 21800
rect 175000 21800 175100 21900
rect 175000 21900 175100 22000
rect 175000 22000 175100 22100
rect 175000 22100 175100 22200
rect 175000 22200 175100 22300
rect 175000 22300 175100 22400
rect 175000 22400 175100 22500
rect 175000 22500 175100 22600
rect 175000 22600 175100 22700
rect 175000 22700 175100 22800
rect 175000 22800 175100 22900
rect 175000 22900 175100 23000
rect 175000 23000 175100 23100
rect 175000 23100 175100 23200
rect 175000 23200 175100 23300
rect 175000 23300 175100 23400
rect 175000 23400 175100 23500
rect 175000 23500 175100 23600
rect 175000 23600 175100 23700
rect 175000 23700 175100 23800
rect 175000 23800 175100 23900
rect 175000 23900 175100 24000
rect 175000 24000 175100 24100
rect 175000 24100 175100 24200
rect 175000 24200 175100 24300
rect 175000 24300 175100 24400
rect 175000 24400 175100 24500
rect 175000 24500 175100 24600
rect 175000 24600 175100 24700
rect 175000 24700 175100 24800
rect 175000 24800 175100 24900
rect 175000 24900 175100 25000
rect 175000 25000 175100 25100
rect 175000 25100 175100 25200
rect 175000 25200 175100 25300
rect 175000 25300 175100 25400
rect 175000 25400 175100 25500
rect 175000 25500 175100 25600
rect 175000 25600 175100 25700
rect 175000 25700 175100 25800
rect 175000 25800 175100 25900
rect 175000 25900 175100 26000
rect 175000 26000 175100 26100
rect 175000 26100 175100 26200
rect 175000 26200 175100 26300
rect 175000 26300 175100 26400
rect 175000 26400 175100 26500
rect 175000 26500 175100 26600
rect 175000 26600 175100 26700
rect 175000 26700 175100 26800
rect 175000 26800 175100 26900
rect 175000 26900 175100 27000
rect 175000 27000 175100 27100
rect 175000 27100 175100 27200
rect 175000 27200 175100 27300
rect 175000 27300 175100 27400
rect 175000 27400 175100 27500
rect 175000 27500 175100 27600
rect 175000 27600 175100 27700
rect 175000 27700 175100 27800
rect 175000 27800 175100 27900
rect 175000 27900 175100 28000
rect 175000 28000 175100 28100
rect 175000 28100 175100 28200
rect 175000 28200 175100 28300
rect 175000 28300 175100 28400
rect 175000 28400 175100 28500
rect 175000 28500 175100 28600
rect 175000 28600 175100 28700
rect 175000 28700 175100 28800
rect 175000 28800 175100 28900
rect 175000 28900 175100 29000
rect 175000 29000 175100 29100
rect 175000 29100 175100 29200
rect 175000 29200 175100 29300
rect 175000 29300 175100 29400
rect 175000 29400 175100 29500
rect 175000 29500 175100 29600
rect 175000 29600 175100 29700
rect 175000 29700 175100 29800
rect 175000 29800 175100 29900
rect 175000 29900 175100 30000
rect 175000 30000 175100 30100
rect 175000 30100 175100 30200
rect 175000 30200 175100 30300
rect 175100 21600 175200 21700
rect 175100 21700 175200 21800
rect 175100 21800 175200 21900
rect 175100 21900 175200 22000
rect 175100 22000 175200 22100
rect 175100 22100 175200 22200
rect 175100 22200 175200 22300
rect 175100 22300 175200 22400
rect 175100 22400 175200 22500
rect 175100 22500 175200 22600
rect 175100 22600 175200 22700
rect 175100 22700 175200 22800
rect 175100 22800 175200 22900
rect 175100 22900 175200 23000
rect 175100 23000 175200 23100
rect 175100 23100 175200 23200
rect 175100 23200 175200 23300
rect 175100 23300 175200 23400
rect 175100 23400 175200 23500
rect 175100 23500 175200 23600
rect 175100 23600 175200 23700
rect 175100 23700 175200 23800
rect 175100 23800 175200 23900
rect 175100 23900 175200 24000
rect 175100 24000 175200 24100
rect 175100 24100 175200 24200
rect 175100 24200 175200 24300
rect 175100 24300 175200 24400
rect 175100 24400 175200 24500
rect 175100 24500 175200 24600
rect 175100 24600 175200 24700
rect 175100 24700 175200 24800
rect 175100 24800 175200 24900
rect 175100 24900 175200 25000
rect 175100 25000 175200 25100
rect 175100 25100 175200 25200
rect 175100 25200 175200 25300
rect 175100 25300 175200 25400
rect 175100 25400 175200 25500
rect 175100 25500 175200 25600
rect 175100 25600 175200 25700
rect 175100 25700 175200 25800
rect 175100 25800 175200 25900
rect 175100 25900 175200 26000
rect 175100 26000 175200 26100
rect 175100 26100 175200 26200
rect 175100 26200 175200 26300
rect 175100 26300 175200 26400
rect 175100 26400 175200 26500
rect 175100 26500 175200 26600
rect 175100 26600 175200 26700
rect 175100 26700 175200 26800
rect 175100 26800 175200 26900
rect 175100 26900 175200 27000
rect 175100 27000 175200 27100
rect 175100 27100 175200 27200
rect 175100 27200 175200 27300
rect 175100 27300 175200 27400
rect 175100 27400 175200 27500
rect 175100 27500 175200 27600
rect 175100 27600 175200 27700
rect 175100 27700 175200 27800
rect 175100 27800 175200 27900
rect 175100 27900 175200 28000
rect 175100 28000 175200 28100
rect 175100 28100 175200 28200
rect 175100 28200 175200 28300
rect 175100 28300 175200 28400
rect 175100 28400 175200 28500
rect 175100 28500 175200 28600
rect 175100 28600 175200 28700
rect 175100 28700 175200 28800
rect 175100 28800 175200 28900
rect 175100 28900 175200 29000
rect 175100 29000 175200 29100
rect 175100 29100 175200 29200
rect 175100 29200 175200 29300
rect 175100 29300 175200 29400
rect 175100 29400 175200 29500
rect 175100 29500 175200 29600
rect 175100 29600 175200 29700
rect 175100 29700 175200 29800
rect 175200 21500 175300 21600
rect 175200 21600 175300 21700
rect 175200 21700 175300 21800
rect 175200 21800 175300 21900
rect 175200 21900 175300 22000
rect 175200 22000 175300 22100
rect 175200 22100 175300 22200
rect 175200 22200 175300 22300
rect 175200 22300 175300 22400
rect 175200 22400 175300 22500
rect 175200 22500 175300 22600
rect 175200 22600 175300 22700
rect 175200 22700 175300 22800
rect 175200 22800 175300 22900
rect 175200 22900 175300 23000
rect 175200 23000 175300 23100
rect 175200 23100 175300 23200
rect 175200 23200 175300 23300
rect 175200 23300 175300 23400
rect 175200 23400 175300 23500
rect 175200 23500 175300 23600
rect 175200 23600 175300 23700
rect 175200 23700 175300 23800
rect 175200 23800 175300 23900
rect 175200 23900 175300 24000
rect 175200 24000 175300 24100
rect 175200 24100 175300 24200
rect 175200 24200 175300 24300
rect 175200 24300 175300 24400
rect 175200 24400 175300 24500
rect 175200 24500 175300 24600
rect 175200 24600 175300 24700
rect 175200 24700 175300 24800
rect 175200 24800 175300 24900
rect 175200 24900 175300 25000
rect 175200 25000 175300 25100
rect 175200 25100 175300 25200
rect 175200 25200 175300 25300
rect 175200 25300 175300 25400
rect 175200 25400 175300 25500
rect 175200 25500 175300 25600
rect 175200 25600 175300 25700
rect 175200 25700 175300 25800
rect 175200 25800 175300 25900
rect 175200 25900 175300 26000
rect 175200 26000 175300 26100
rect 175200 26100 175300 26200
rect 175200 26200 175300 26300
rect 175200 26300 175300 26400
rect 175200 26400 175300 26500
rect 175200 26500 175300 26600
rect 175200 26600 175300 26700
rect 175200 26700 175300 26800
rect 175200 26800 175300 26900
rect 175200 26900 175300 27000
rect 175200 27000 175300 27100
rect 175200 27100 175300 27200
rect 175200 27200 175300 27300
rect 175200 27300 175300 27400
rect 175200 27400 175300 27500
rect 175200 27500 175300 27600
rect 175200 27600 175300 27700
rect 175200 27700 175300 27800
rect 175200 27800 175300 27900
rect 175200 27900 175300 28000
rect 175200 28000 175300 28100
rect 175200 28100 175300 28200
rect 175200 28200 175300 28300
rect 175200 28300 175300 28400
rect 175200 28400 175300 28500
rect 175200 28500 175300 28600
rect 175200 28600 175300 28700
rect 175200 28700 175300 28800
rect 175200 28800 175300 28900
rect 175200 28900 175300 29000
rect 175200 29000 175300 29100
rect 175200 29100 175300 29200
rect 175200 29200 175300 29300
rect 175300 21400 175400 21500
rect 175300 21500 175400 21600
rect 175300 21600 175400 21700
rect 175300 21700 175400 21800
rect 175300 21800 175400 21900
rect 175300 21900 175400 22000
rect 175300 22000 175400 22100
rect 175300 22100 175400 22200
rect 175300 22200 175400 22300
rect 175300 22300 175400 22400
rect 175300 22400 175400 22500
rect 175300 22500 175400 22600
rect 175300 22600 175400 22700
rect 175300 22700 175400 22800
rect 175300 22800 175400 22900
rect 175300 22900 175400 23000
rect 175300 23000 175400 23100
rect 175300 23100 175400 23200
rect 175300 23200 175400 23300
rect 175300 23300 175400 23400
rect 175300 23400 175400 23500
rect 175300 23500 175400 23600
rect 175300 23600 175400 23700
rect 175300 23700 175400 23800
rect 175300 23800 175400 23900
rect 175300 23900 175400 24000
rect 175300 24000 175400 24100
rect 175300 24100 175400 24200
rect 175300 24200 175400 24300
rect 175300 24300 175400 24400
rect 175300 24400 175400 24500
rect 175300 24500 175400 24600
rect 175300 24600 175400 24700
rect 175300 24700 175400 24800
rect 175300 24800 175400 24900
rect 175300 24900 175400 25000
rect 175300 25000 175400 25100
rect 175300 25100 175400 25200
rect 175300 25200 175400 25300
rect 175300 25300 175400 25400
rect 175300 25400 175400 25500
rect 175300 25500 175400 25600
rect 175300 25600 175400 25700
rect 175300 25700 175400 25800
rect 175300 25800 175400 25900
rect 175300 25900 175400 26000
rect 175300 26000 175400 26100
rect 175300 26100 175400 26200
rect 175300 26200 175400 26300
rect 175300 26300 175400 26400
rect 175300 26400 175400 26500
rect 175300 26500 175400 26600
rect 175300 26600 175400 26700
rect 175300 26700 175400 26800
rect 175300 26800 175400 26900
rect 175300 26900 175400 27000
rect 175300 27000 175400 27100
rect 175300 27100 175400 27200
rect 175300 27200 175400 27300
rect 175300 27300 175400 27400
rect 175300 27400 175400 27500
rect 175300 27500 175400 27600
rect 175300 27600 175400 27700
rect 175300 27700 175400 27800
rect 175300 27800 175400 27900
rect 175300 27900 175400 28000
rect 175300 28000 175400 28100
rect 175300 28100 175400 28200
rect 175300 28200 175400 28300
rect 175300 28300 175400 28400
rect 175300 28400 175400 28500
rect 175300 28500 175400 28600
rect 175300 28600 175400 28700
rect 175300 28700 175400 28800
rect 175400 21400 175500 21500
rect 175400 21500 175500 21600
rect 175400 21600 175500 21700
rect 175400 21700 175500 21800
rect 175400 21800 175500 21900
rect 175400 21900 175500 22000
rect 175400 22000 175500 22100
rect 175400 22100 175500 22200
rect 175400 22200 175500 22300
rect 175400 22300 175500 22400
rect 175400 22400 175500 22500
rect 175400 22500 175500 22600
rect 175400 22600 175500 22700
rect 175400 22700 175500 22800
rect 175400 22800 175500 22900
rect 175400 22900 175500 23000
rect 175400 23000 175500 23100
rect 175400 23100 175500 23200
rect 175400 23200 175500 23300
rect 175400 23300 175500 23400
rect 175400 23400 175500 23500
rect 175400 23500 175500 23600
rect 175400 23600 175500 23700
rect 175400 23700 175500 23800
rect 175400 23800 175500 23900
rect 175400 23900 175500 24000
rect 175400 24000 175500 24100
rect 175400 24100 175500 24200
rect 175400 24200 175500 24300
rect 175400 24300 175500 24400
rect 175400 24400 175500 24500
rect 175400 24500 175500 24600
rect 175400 24600 175500 24700
rect 175400 24700 175500 24800
rect 175400 24800 175500 24900
rect 175400 24900 175500 25000
rect 175400 25000 175500 25100
rect 175400 25100 175500 25200
rect 175400 25200 175500 25300
rect 175400 25300 175500 25400
rect 175400 25400 175500 25500
rect 175400 25500 175500 25600
rect 175400 25600 175500 25700
rect 175400 25700 175500 25800
rect 175400 25800 175500 25900
rect 175400 25900 175500 26000
rect 175400 26000 175500 26100
rect 175400 26100 175500 26200
rect 175400 26200 175500 26300
rect 175400 26300 175500 26400
rect 175400 26400 175500 26500
rect 175400 26500 175500 26600
rect 175400 26600 175500 26700
rect 175400 26700 175500 26800
rect 175400 26800 175500 26900
rect 175400 26900 175500 27000
rect 175400 27000 175500 27100
rect 175400 27100 175500 27200
rect 175400 27200 175500 27300
rect 175400 27300 175500 27400
rect 175400 27400 175500 27500
rect 175400 27500 175500 27600
rect 175400 27600 175500 27700
rect 175400 27700 175500 27800
rect 175400 27800 175500 27900
rect 175400 27900 175500 28000
rect 175400 28000 175500 28100
rect 175400 28100 175500 28200
rect 175400 28200 175500 28300
rect 175500 21400 175600 21500
rect 175500 21500 175600 21600
rect 175500 21600 175600 21700
rect 175500 21700 175600 21800
rect 175500 21800 175600 21900
rect 175500 21900 175600 22000
rect 175500 22000 175600 22100
rect 175500 22100 175600 22200
rect 175500 22200 175600 22300
rect 175500 22300 175600 22400
rect 175500 22400 175600 22500
rect 175500 22500 175600 22600
rect 175500 22600 175600 22700
rect 175500 22700 175600 22800
rect 175500 22800 175600 22900
rect 175500 22900 175600 23000
rect 175500 23000 175600 23100
rect 175500 23100 175600 23200
rect 175500 23200 175600 23300
rect 175500 23300 175600 23400
rect 175500 23400 175600 23500
rect 175500 23500 175600 23600
rect 175500 23600 175600 23700
rect 175500 23700 175600 23800
rect 175500 23800 175600 23900
rect 175500 23900 175600 24000
rect 175500 24000 175600 24100
rect 175500 24100 175600 24200
rect 175500 24200 175600 24300
rect 175500 24300 175600 24400
rect 175500 24400 175600 24500
rect 175500 24500 175600 24600
rect 175500 24600 175600 24700
rect 175500 24700 175600 24800
rect 175500 24800 175600 24900
rect 175500 24900 175600 25000
rect 175500 25000 175600 25100
rect 175500 25100 175600 25200
rect 175500 25200 175600 25300
rect 175500 25300 175600 25400
rect 175500 25400 175600 25500
rect 175500 25500 175600 25600
rect 175500 25600 175600 25700
rect 175500 25700 175600 25800
rect 175500 25800 175600 25900
rect 175500 25900 175600 26000
rect 175500 26000 175600 26100
rect 175500 26100 175600 26200
rect 175500 26200 175600 26300
rect 175500 26300 175600 26400
rect 175500 26400 175600 26500
rect 175500 26500 175600 26600
rect 175500 26600 175600 26700
rect 175500 26700 175600 26800
rect 175500 26800 175600 26900
rect 175500 26900 175600 27000
rect 175500 27000 175600 27100
rect 175500 27100 175600 27200
rect 175500 27200 175600 27300
rect 175500 27300 175600 27400
rect 175500 27400 175600 27500
rect 175500 27500 175600 27600
rect 175500 27600 175600 27700
rect 175500 27700 175600 27800
rect 175500 27800 175600 27900
rect 175600 21300 175700 21400
rect 175600 21400 175700 21500
rect 175600 21500 175700 21600
rect 175600 21600 175700 21700
rect 175600 21700 175700 21800
rect 175600 21800 175700 21900
rect 175600 21900 175700 22000
rect 175600 22000 175700 22100
rect 175600 22100 175700 22200
rect 175600 22200 175700 22300
rect 175600 22300 175700 22400
rect 175600 22400 175700 22500
rect 175600 22500 175700 22600
rect 175600 22600 175700 22700
rect 175600 22700 175700 22800
rect 175600 22800 175700 22900
rect 175600 22900 175700 23000
rect 175600 23000 175700 23100
rect 175600 23100 175700 23200
rect 175600 23200 175700 23300
rect 175600 23300 175700 23400
rect 175600 23400 175700 23500
rect 175600 23500 175700 23600
rect 175600 23600 175700 23700
rect 175600 23700 175700 23800
rect 175600 23800 175700 23900
rect 175600 23900 175700 24000
rect 175600 24000 175700 24100
rect 175600 24100 175700 24200
rect 175600 24200 175700 24300
rect 175600 24300 175700 24400
rect 175600 24400 175700 24500
rect 175600 24500 175700 24600
rect 175600 24600 175700 24700
rect 175600 24700 175700 24800
rect 175600 24800 175700 24900
rect 175600 24900 175700 25000
rect 175600 25000 175700 25100
rect 175600 25100 175700 25200
rect 175600 25200 175700 25300
rect 175600 25300 175700 25400
rect 175600 25400 175700 25500
rect 175600 25500 175700 25600
rect 175600 25600 175700 25700
rect 175600 25700 175700 25800
rect 175600 25800 175700 25900
rect 175600 25900 175700 26000
rect 175600 26000 175700 26100
rect 175600 26100 175700 26200
rect 175600 26200 175700 26300
rect 175600 26300 175700 26400
rect 175600 26400 175700 26500
rect 175600 26500 175700 26600
rect 175600 26600 175700 26700
rect 175600 26700 175700 26800
rect 175600 26800 175700 26900
rect 175600 26900 175700 27000
rect 175600 27000 175700 27100
rect 175600 27100 175700 27200
rect 175600 27200 175700 27300
rect 175600 27300 175700 27400
rect 175700 21300 175800 21400
rect 175700 21400 175800 21500
rect 175700 21500 175800 21600
rect 175700 21600 175800 21700
rect 175700 21700 175800 21800
rect 175700 21800 175800 21900
rect 175700 21900 175800 22000
rect 175700 22000 175800 22100
rect 175700 22100 175800 22200
rect 175700 22200 175800 22300
rect 175700 22300 175800 22400
rect 175700 22400 175800 22500
rect 175700 22500 175800 22600
rect 175700 22600 175800 22700
rect 175700 22700 175800 22800
rect 175700 22800 175800 22900
rect 175700 22900 175800 23000
rect 175700 23000 175800 23100
rect 175700 23100 175800 23200
rect 175700 23200 175800 23300
rect 175700 23300 175800 23400
rect 175700 23400 175800 23500
rect 175700 23500 175800 23600
rect 175700 23600 175800 23700
rect 175700 23700 175800 23800
rect 175700 23800 175800 23900
rect 175700 23900 175800 24000
rect 175700 24000 175800 24100
rect 175700 24100 175800 24200
rect 175700 24200 175800 24300
rect 175700 24300 175800 24400
rect 175700 24400 175800 24500
rect 175700 24500 175800 24600
rect 175700 24600 175800 24700
rect 175700 24700 175800 24800
rect 175700 24800 175800 24900
rect 175700 24900 175800 25000
rect 175700 25000 175800 25100
rect 175700 25100 175800 25200
rect 175700 25200 175800 25300
rect 175700 25300 175800 25400
rect 175700 25400 175800 25500
rect 175700 25500 175800 25600
rect 175700 25600 175800 25700
rect 175700 25700 175800 25800
rect 175700 25800 175800 25900
rect 175700 25900 175800 26000
rect 175700 26000 175800 26100
rect 175700 26100 175800 26200
rect 175700 26200 175800 26300
rect 175700 26300 175800 26400
rect 175700 26400 175800 26500
rect 175700 26500 175800 26600
rect 175700 26600 175800 26700
rect 175700 26700 175800 26800
rect 175700 26800 175800 26900
rect 175700 26900 175800 27000
rect 175800 21300 175900 21400
rect 175800 21400 175900 21500
rect 175800 21500 175900 21600
rect 175800 21600 175900 21700
rect 175800 21700 175900 21800
rect 175800 21800 175900 21900
rect 175800 21900 175900 22000
rect 175800 22000 175900 22100
rect 175800 22100 175900 22200
rect 175800 22200 175900 22300
rect 175800 22300 175900 22400
rect 175800 22400 175900 22500
rect 175800 22500 175900 22600
rect 175800 22600 175900 22700
rect 175800 22700 175900 22800
rect 175800 22800 175900 22900
rect 175800 22900 175900 23000
rect 175800 23000 175900 23100
rect 175800 23100 175900 23200
rect 175800 23200 175900 23300
rect 175800 23300 175900 23400
rect 175800 23400 175900 23500
rect 175800 23500 175900 23600
rect 175800 23600 175900 23700
rect 175800 23700 175900 23800
rect 175800 23800 175900 23900
rect 175800 23900 175900 24000
rect 175800 24000 175900 24100
rect 175800 24100 175900 24200
rect 175800 24200 175900 24300
rect 175800 24300 175900 24400
rect 175800 24400 175900 24500
rect 175800 24500 175900 24600
rect 175800 24600 175900 24700
rect 175800 24700 175900 24800
rect 175800 24800 175900 24900
rect 175800 24900 175900 25000
rect 175800 25000 175900 25100
rect 175800 25100 175900 25200
rect 175800 25200 175900 25300
rect 175800 25300 175900 25400
rect 175800 25400 175900 25500
rect 175800 25500 175900 25600
rect 175800 25600 175900 25700
rect 175800 25700 175900 25800
rect 175800 25800 175900 25900
rect 175800 25900 175900 26000
rect 175800 26000 175900 26100
rect 175800 26100 175900 26200
rect 175800 26200 175900 26300
rect 175800 26300 175900 26400
rect 175800 26400 175900 26500
rect 175900 21300 176000 21400
rect 175900 21400 176000 21500
rect 175900 21500 176000 21600
rect 175900 21600 176000 21700
rect 175900 21700 176000 21800
rect 175900 21800 176000 21900
rect 175900 21900 176000 22000
rect 175900 22000 176000 22100
rect 175900 22100 176000 22200
rect 175900 22200 176000 22300
rect 175900 22300 176000 22400
rect 175900 22400 176000 22500
rect 175900 22500 176000 22600
rect 175900 22600 176000 22700
rect 175900 22700 176000 22800
rect 175900 22800 176000 22900
rect 175900 22900 176000 23000
rect 175900 23000 176000 23100
rect 175900 23100 176000 23200
rect 175900 23200 176000 23300
rect 175900 23300 176000 23400
rect 175900 23400 176000 23500
rect 175900 23500 176000 23600
rect 175900 23600 176000 23700
rect 175900 23700 176000 23800
rect 175900 23800 176000 23900
rect 175900 23900 176000 24000
rect 175900 24000 176000 24100
rect 175900 24100 176000 24200
rect 175900 24200 176000 24300
rect 175900 24300 176000 24400
rect 175900 24400 176000 24500
rect 175900 24500 176000 24600
rect 175900 24600 176000 24700
rect 175900 24700 176000 24800
rect 175900 24800 176000 24900
rect 175900 24900 176000 25000
rect 175900 25000 176000 25100
rect 175900 25100 176000 25200
rect 175900 25200 176000 25300
rect 175900 25300 176000 25400
rect 175900 25400 176000 25500
rect 175900 25500 176000 25600
rect 175900 25600 176000 25700
rect 175900 25700 176000 25800
rect 175900 25800 176000 25900
rect 175900 25900 176000 26000
rect 175900 26000 176000 26100
rect 176000 21300 176100 21400
rect 176000 21400 176100 21500
rect 176000 21500 176100 21600
rect 176000 21600 176100 21700
rect 176000 21700 176100 21800
rect 176000 21800 176100 21900
rect 176000 21900 176100 22000
rect 176000 22000 176100 22100
rect 176000 22100 176100 22200
rect 176000 22200 176100 22300
rect 176000 22300 176100 22400
rect 176000 22400 176100 22500
rect 176000 22500 176100 22600
rect 176000 22600 176100 22700
rect 176000 22700 176100 22800
rect 176000 22800 176100 22900
rect 176000 22900 176100 23000
rect 176000 23000 176100 23100
rect 176000 23100 176100 23200
rect 176000 23200 176100 23300
rect 176000 23300 176100 23400
rect 176000 23400 176100 23500
rect 176000 23500 176100 23600
rect 176000 23600 176100 23700
rect 176000 23700 176100 23800
rect 176000 23800 176100 23900
rect 176000 23900 176100 24000
rect 176000 24000 176100 24100
rect 176000 24100 176100 24200
rect 176000 24200 176100 24300
rect 176000 24300 176100 24400
rect 176000 24400 176100 24500
rect 176000 24500 176100 24600
rect 176000 24600 176100 24700
rect 176000 24700 176100 24800
rect 176000 24800 176100 24900
rect 176000 24900 176100 25000
rect 176000 25000 176100 25100
rect 176000 25100 176100 25200
rect 176000 25200 176100 25300
rect 176000 25300 176100 25400
rect 176000 25400 176100 25500
rect 176000 25500 176100 25600
rect 176100 21300 176200 21400
rect 176100 21400 176200 21500
rect 176100 21500 176200 21600
rect 176100 21600 176200 21700
rect 176100 21700 176200 21800
rect 176100 21800 176200 21900
rect 176100 21900 176200 22000
rect 176100 22000 176200 22100
rect 176100 22100 176200 22200
rect 176100 22200 176200 22300
rect 176100 22300 176200 22400
rect 176100 22400 176200 22500
rect 176100 22500 176200 22600
rect 176100 22600 176200 22700
rect 176100 22700 176200 22800
rect 176100 22800 176200 22900
rect 176100 22900 176200 23000
rect 176100 23000 176200 23100
rect 176100 23100 176200 23200
rect 176100 23200 176200 23300
rect 176100 23300 176200 23400
rect 176100 23400 176200 23500
rect 176100 23500 176200 23600
rect 176100 23600 176200 23700
rect 176100 23700 176200 23800
rect 176100 23800 176200 23900
rect 176100 23900 176200 24000
rect 176100 24000 176200 24100
rect 176100 24100 176200 24200
rect 176100 24200 176200 24300
rect 176100 24300 176200 24400
rect 176100 24400 176200 24500
rect 176100 24500 176200 24600
rect 176100 24600 176200 24700
rect 176100 24700 176200 24800
rect 176100 24800 176200 24900
rect 176100 24900 176200 25000
rect 176100 25000 176200 25100
rect 176200 21300 176300 21400
rect 176200 21400 176300 21500
rect 176200 21500 176300 21600
rect 176200 21600 176300 21700
rect 176200 21700 176300 21800
rect 176200 21800 176300 21900
rect 176200 21900 176300 22000
rect 176200 22000 176300 22100
rect 176200 22100 176300 22200
rect 176200 22200 176300 22300
rect 176200 22300 176300 22400
rect 176200 22400 176300 22500
rect 176200 22500 176300 22600
rect 176200 22600 176300 22700
rect 176200 22700 176300 22800
rect 176200 22800 176300 22900
rect 176200 22900 176300 23000
rect 176200 23000 176300 23100
rect 176200 23100 176300 23200
rect 176200 23200 176300 23300
rect 176200 23300 176300 23400
rect 176200 23400 176300 23500
rect 176200 23500 176300 23600
rect 176200 23600 176300 23700
rect 176200 23700 176300 23800
rect 176200 23800 176300 23900
rect 176200 23900 176300 24000
rect 176200 24000 176300 24100
rect 176200 24100 176300 24200
rect 176200 24200 176300 24300
rect 176200 24300 176300 24400
rect 176200 24400 176300 24500
rect 176200 24500 176300 24600
rect 176200 24600 176300 24700
rect 176200 24700 176300 24800
rect 176300 21300 176400 21400
rect 176300 21400 176400 21500
rect 176300 21500 176400 21600
rect 176300 21600 176400 21700
rect 176300 21700 176400 21800
rect 176300 21800 176400 21900
rect 176300 21900 176400 22000
rect 176300 22000 176400 22100
rect 176300 22100 176400 22200
rect 176300 22200 176400 22300
rect 176300 22300 176400 22400
rect 176300 22400 176400 22500
rect 176300 22500 176400 22600
rect 176300 22600 176400 22700
rect 176300 22700 176400 22800
rect 176300 22800 176400 22900
rect 176300 22900 176400 23000
rect 176300 23000 176400 23100
rect 176300 23100 176400 23200
rect 176300 23200 176400 23300
rect 176300 23300 176400 23400
rect 176300 23400 176400 23500
rect 176300 23500 176400 23600
rect 176300 23600 176400 23700
rect 176300 23700 176400 23800
rect 176300 23800 176400 23900
rect 176300 23900 176400 24000
rect 176300 24000 176400 24100
rect 176300 24100 176400 24200
rect 176300 24200 176400 24300
rect 176300 24300 176400 24400
rect 176300 24400 176400 24500
rect 176300 24500 176400 24600
rect 176300 24600 176400 24700
rect 176300 24700 176400 24800
rect 176300 24800 176400 24900
rect 176300 24900 176400 25000
rect 176400 21400 176500 21500
rect 176400 21500 176500 21600
rect 176400 21600 176500 21700
rect 176400 21700 176500 21800
rect 176400 21800 176500 21900
rect 176400 21900 176500 22000
rect 176400 22000 176500 22100
rect 176400 22100 176500 22200
rect 176400 22200 176500 22300
rect 176400 22300 176500 22400
rect 176400 22400 176500 22500
rect 176400 22500 176500 22600
rect 176400 22600 176500 22700
rect 176400 22700 176500 22800
rect 176400 22800 176500 22900
rect 176400 22900 176500 23000
rect 176400 23000 176500 23100
rect 176400 23100 176500 23200
rect 176400 23200 176500 23300
rect 176400 23300 176500 23400
rect 176400 23400 176500 23500
rect 176400 23500 176500 23600
rect 176400 23600 176500 23700
rect 176400 23700 176500 23800
rect 176400 23800 176500 23900
rect 176400 23900 176500 24000
rect 176400 24000 176500 24100
rect 176400 24100 176500 24200
rect 176400 24200 176500 24300
rect 176400 24300 176500 24400
rect 176400 24400 176500 24500
rect 176400 24500 176500 24600
rect 176400 24600 176500 24700
rect 176400 24700 176500 24800
rect 176400 24800 176500 24900
rect 176400 24900 176500 25000
rect 176400 25000 176500 25100
rect 176400 25100 176500 25200
rect 176500 21400 176600 21500
rect 176500 21500 176600 21600
rect 176500 21600 176600 21700
rect 176500 21700 176600 21800
rect 176500 21800 176600 21900
rect 176500 21900 176600 22000
rect 176500 22000 176600 22100
rect 176500 22100 176600 22200
rect 176500 22200 176600 22300
rect 176500 22300 176600 22400
rect 176500 22400 176600 22500
rect 176500 22500 176600 22600
rect 176500 22600 176600 22700
rect 176500 22700 176600 22800
rect 176500 22800 176600 22900
rect 176500 22900 176600 23000
rect 176500 23000 176600 23100
rect 176500 23100 176600 23200
rect 176500 23200 176600 23300
rect 176500 23300 176600 23400
rect 176500 23400 176600 23500
rect 176500 23500 176600 23600
rect 176500 23600 176600 23700
rect 176500 23700 176600 23800
rect 176500 23800 176600 23900
rect 176500 23900 176600 24000
rect 176500 24000 176600 24100
rect 176500 24100 176600 24200
rect 176500 24200 176600 24300
rect 176500 24300 176600 24400
rect 176500 24400 176600 24500
rect 176500 24500 176600 24600
rect 176500 24600 176600 24700
rect 176500 24700 176600 24800
rect 176500 24800 176600 24900
rect 176500 24900 176600 25000
rect 176500 25000 176600 25100
rect 176500 25100 176600 25200
rect 176500 25200 176600 25300
rect 176500 25300 176600 25400
rect 176600 21400 176700 21500
rect 176600 21500 176700 21600
rect 176600 21600 176700 21700
rect 176600 21700 176700 21800
rect 176600 21800 176700 21900
rect 176600 21900 176700 22000
rect 176600 22000 176700 22100
rect 176600 22100 176700 22200
rect 176600 22200 176700 22300
rect 176600 22300 176700 22400
rect 176600 22400 176700 22500
rect 176600 22500 176700 22600
rect 176600 22600 176700 22700
rect 176600 22700 176700 22800
rect 176600 22800 176700 22900
rect 176600 22900 176700 23000
rect 176600 23000 176700 23100
rect 176600 23100 176700 23200
rect 176600 23200 176700 23300
rect 176600 23300 176700 23400
rect 176600 23400 176700 23500
rect 176600 23500 176700 23600
rect 176600 23600 176700 23700
rect 176600 23700 176700 23800
rect 176600 23800 176700 23900
rect 176600 23900 176700 24000
rect 176600 24000 176700 24100
rect 176600 24100 176700 24200
rect 176600 24200 176700 24300
rect 176600 24300 176700 24400
rect 176600 24400 176700 24500
rect 176600 24500 176700 24600
rect 176600 24600 176700 24700
rect 176600 24700 176700 24800
rect 176600 24800 176700 24900
rect 176600 24900 176700 25000
rect 176600 25000 176700 25100
rect 176600 25100 176700 25200
rect 176600 25200 176700 25300
rect 176600 25300 176700 25400
rect 176600 25400 176700 25500
rect 176600 25500 176700 25600
rect 176600 25600 176700 25700
rect 176700 21500 176800 21600
rect 176700 21600 176800 21700
rect 176700 21700 176800 21800
rect 176700 21800 176800 21900
rect 176700 21900 176800 22000
rect 176700 22000 176800 22100
rect 176700 22100 176800 22200
rect 176700 22200 176800 22300
rect 176700 22300 176800 22400
rect 176700 22400 176800 22500
rect 176700 22500 176800 22600
rect 176700 22600 176800 22700
rect 176700 22700 176800 22800
rect 176700 22800 176800 22900
rect 176700 22900 176800 23000
rect 176700 23000 176800 23100
rect 176700 23100 176800 23200
rect 176700 23200 176800 23300
rect 176700 23300 176800 23400
rect 176700 23400 176800 23500
rect 176700 23500 176800 23600
rect 176700 23600 176800 23700
rect 176700 23700 176800 23800
rect 176700 23800 176800 23900
rect 176700 23900 176800 24000
rect 176700 24000 176800 24100
rect 176700 24100 176800 24200
rect 176700 24200 176800 24300
rect 176700 24300 176800 24400
rect 176700 24400 176800 24500
rect 176700 24500 176800 24600
rect 176700 24600 176800 24700
rect 176700 24700 176800 24800
rect 176700 24800 176800 24900
rect 176700 24900 176800 25000
rect 176700 25000 176800 25100
rect 176700 25100 176800 25200
rect 176700 25200 176800 25300
rect 176700 25300 176800 25400
rect 176700 25400 176800 25500
rect 176700 25500 176800 25600
rect 176700 25600 176800 25700
rect 176700 25700 176800 25800
rect 176700 25800 176800 25900
rect 176800 21600 176900 21700
rect 176800 21700 176900 21800
rect 176800 21800 176900 21900
rect 176800 21900 176900 22000
rect 176800 22000 176900 22100
rect 176800 22100 176900 22200
rect 176800 22200 176900 22300
rect 176800 22300 176900 22400
rect 176800 22400 176900 22500
rect 176800 22500 176900 22600
rect 176800 22600 176900 22700
rect 176800 22700 176900 22800
rect 176800 22800 176900 22900
rect 176800 22900 176900 23000
rect 176800 23000 176900 23100
rect 176800 23100 176900 23200
rect 176800 23200 176900 23300
rect 176800 23300 176900 23400
rect 176800 23400 176900 23500
rect 176800 23500 176900 23600
rect 176800 23600 176900 23700
rect 176800 23700 176900 23800
rect 176800 23800 176900 23900
rect 176800 23900 176900 24000
rect 176800 24000 176900 24100
rect 176800 24100 176900 24200
rect 176800 24200 176900 24300
rect 176800 24300 176900 24400
rect 176800 24400 176900 24500
rect 176800 24500 176900 24600
rect 176800 24600 176900 24700
rect 176800 24700 176900 24800
rect 176800 24800 176900 24900
rect 176800 24900 176900 25000
rect 176800 25000 176900 25100
rect 176800 25100 176900 25200
rect 176800 25200 176900 25300
rect 176800 25300 176900 25400
rect 176800 25400 176900 25500
rect 176800 25500 176900 25600
rect 176800 25600 176900 25700
rect 176800 25700 176900 25800
rect 176800 25800 176900 25900
rect 176800 25900 176900 26000
rect 176800 26000 176900 26100
rect 176800 26100 176900 26200
rect 176900 21700 177000 21800
rect 176900 21800 177000 21900
rect 176900 21900 177000 22000
rect 176900 22000 177000 22100
rect 176900 22100 177000 22200
rect 176900 22200 177000 22300
rect 176900 22300 177000 22400
rect 176900 22400 177000 22500
rect 176900 22500 177000 22600
rect 176900 22600 177000 22700
rect 176900 22700 177000 22800
rect 176900 22800 177000 22900
rect 176900 22900 177000 23000
rect 176900 23000 177000 23100
rect 176900 23100 177000 23200
rect 176900 23200 177000 23300
rect 176900 23300 177000 23400
rect 176900 23400 177000 23500
rect 176900 23500 177000 23600
rect 176900 23600 177000 23700
rect 176900 23700 177000 23800
rect 176900 23800 177000 23900
rect 176900 23900 177000 24000
rect 176900 24000 177000 24100
rect 176900 24100 177000 24200
rect 176900 24200 177000 24300
rect 176900 24300 177000 24400
rect 176900 24400 177000 24500
rect 176900 24500 177000 24600
rect 176900 24600 177000 24700
rect 176900 24700 177000 24800
rect 176900 24800 177000 24900
rect 176900 24900 177000 25000
rect 176900 25000 177000 25100
rect 176900 25100 177000 25200
rect 176900 25200 177000 25300
rect 176900 25300 177000 25400
rect 176900 25400 177000 25500
rect 176900 25500 177000 25600
rect 176900 25600 177000 25700
rect 176900 25700 177000 25800
rect 176900 25800 177000 25900
rect 176900 25900 177000 26000
rect 176900 26000 177000 26100
rect 176900 26100 177000 26200
rect 176900 26200 177000 26300
rect 176900 26300 177000 26400
rect 177000 21800 177100 21900
rect 177000 21900 177100 22000
rect 177000 22000 177100 22100
rect 177000 22100 177100 22200
rect 177000 22200 177100 22300
rect 177000 22300 177100 22400
rect 177000 22400 177100 22500
rect 177000 22500 177100 22600
rect 177000 22600 177100 22700
rect 177000 22700 177100 22800
rect 177000 22800 177100 22900
rect 177000 22900 177100 23000
rect 177000 23000 177100 23100
rect 177000 23100 177100 23200
rect 177000 23200 177100 23300
rect 177000 23300 177100 23400
rect 177000 23400 177100 23500
rect 177000 23500 177100 23600
rect 177000 23600 177100 23700
rect 177000 23700 177100 23800
rect 177000 23800 177100 23900
rect 177000 23900 177100 24000
rect 177000 24000 177100 24100
rect 177000 24100 177100 24200
rect 177000 24200 177100 24300
rect 177000 24300 177100 24400
rect 177000 24400 177100 24500
rect 177000 24500 177100 24600
rect 177000 24600 177100 24700
rect 177000 24700 177100 24800
rect 177000 24800 177100 24900
rect 177000 24900 177100 25000
rect 177000 25000 177100 25100
rect 177000 25100 177100 25200
rect 177000 25200 177100 25300
rect 177000 25300 177100 25400
rect 177000 25400 177100 25500
rect 177000 25500 177100 25600
rect 177000 25600 177100 25700
rect 177000 25700 177100 25800
rect 177000 25800 177100 25900
rect 177000 25900 177100 26000
rect 177000 26000 177100 26100
rect 177000 26100 177100 26200
rect 177000 26200 177100 26300
rect 177000 26300 177100 26400
rect 177000 26400 177100 26500
rect 177000 26500 177100 26600
rect 177000 26600 177100 26700
rect 177100 22000 177200 22100
rect 177100 22100 177200 22200
rect 177100 22200 177200 22300
rect 177100 22300 177200 22400
rect 177100 22400 177200 22500
rect 177100 22500 177200 22600
rect 177100 22600 177200 22700
rect 177100 22700 177200 22800
rect 177100 22800 177200 22900
rect 177100 22900 177200 23000
rect 177100 23000 177200 23100
rect 177100 23100 177200 23200
rect 177100 23200 177200 23300
rect 177100 23300 177200 23400
rect 177100 23400 177200 23500
rect 177100 23500 177200 23600
rect 177100 23600 177200 23700
rect 177100 23700 177200 23800
rect 177100 23800 177200 23900
rect 177100 23900 177200 24000
rect 177100 24000 177200 24100
rect 177100 24100 177200 24200
rect 177100 24200 177200 24300
rect 177100 24300 177200 24400
rect 177100 24400 177200 24500
rect 177100 24500 177200 24600
rect 177100 24600 177200 24700
rect 177100 24700 177200 24800
rect 177100 24800 177200 24900
rect 177100 24900 177200 25000
rect 177100 25000 177200 25100
rect 177100 25100 177200 25200
rect 177100 25200 177200 25300
rect 177100 25300 177200 25400
rect 177100 25400 177200 25500
rect 177100 25500 177200 25600
rect 177100 25600 177200 25700
rect 177100 25700 177200 25800
rect 177100 25800 177200 25900
rect 177100 25900 177200 26000
rect 177100 26000 177200 26100
rect 177100 26100 177200 26200
rect 177100 26200 177200 26300
rect 177100 26300 177200 26400
rect 177100 26400 177200 26500
rect 177100 26500 177200 26600
rect 177100 26600 177200 26700
rect 177100 26700 177200 26800
rect 177100 26800 177200 26900
rect 177200 22200 177300 22300
rect 177200 22300 177300 22400
rect 177200 22400 177300 22500
rect 177200 22500 177300 22600
rect 177200 22600 177300 22700
rect 177200 22700 177300 22800
rect 177200 22800 177300 22900
rect 177200 22900 177300 23000
rect 177200 23000 177300 23100
rect 177200 23100 177300 23200
rect 177200 23200 177300 23300
rect 177200 23300 177300 23400
rect 177200 23400 177300 23500
rect 177200 23500 177300 23600
rect 177200 23600 177300 23700
rect 177200 23700 177300 23800
rect 177200 23800 177300 23900
rect 177200 23900 177300 24000
rect 177200 24000 177300 24100
rect 177200 24100 177300 24200
rect 177200 24200 177300 24300
rect 177200 24300 177300 24400
rect 177200 24400 177300 24500
rect 177200 24500 177300 24600
rect 177200 24600 177300 24700
rect 177200 24700 177300 24800
rect 177200 24800 177300 24900
rect 177200 24900 177300 25000
rect 177200 25000 177300 25100
rect 177200 25100 177300 25200
rect 177200 25200 177300 25300
rect 177200 25300 177300 25400
rect 177200 25400 177300 25500
rect 177200 25500 177300 25600
rect 177200 25600 177300 25700
rect 177200 25700 177300 25800
rect 177200 25800 177300 25900
rect 177200 25900 177300 26000
rect 177200 26000 177300 26100
rect 177200 26100 177300 26200
rect 177200 26200 177300 26300
rect 177200 26300 177300 26400
rect 177200 26400 177300 26500
rect 177200 26500 177300 26600
rect 177200 26600 177300 26700
rect 177200 26700 177300 26800
rect 177200 26800 177300 26900
rect 177200 26900 177300 27000
rect 177200 27000 177300 27100
rect 177200 27100 177300 27200
rect 177300 22400 177400 22500
rect 177300 22500 177400 22600
rect 177300 22600 177400 22700
rect 177300 22700 177400 22800
rect 177300 22800 177400 22900
rect 177300 22900 177400 23000
rect 177300 23000 177400 23100
rect 177300 23100 177400 23200
rect 177300 23200 177400 23300
rect 177300 23300 177400 23400
rect 177300 23400 177400 23500
rect 177300 23500 177400 23600
rect 177300 23600 177400 23700
rect 177300 23700 177400 23800
rect 177300 23800 177400 23900
rect 177300 23900 177400 24000
rect 177300 24000 177400 24100
rect 177300 24100 177400 24200
rect 177300 24200 177400 24300
rect 177300 24300 177400 24400
rect 177300 24400 177400 24500
rect 177300 24500 177400 24600
rect 177300 24600 177400 24700
rect 177300 24700 177400 24800
rect 177300 24800 177400 24900
rect 177300 24900 177400 25000
rect 177300 25000 177400 25100
rect 177300 25100 177400 25200
rect 177300 25200 177400 25300
rect 177300 25300 177400 25400
rect 177300 25400 177400 25500
rect 177300 25500 177400 25600
rect 177300 25600 177400 25700
rect 177300 25700 177400 25800
rect 177300 25800 177400 25900
rect 177300 25900 177400 26000
rect 177300 26000 177400 26100
rect 177300 26100 177400 26200
rect 177300 26200 177400 26300
rect 177300 26300 177400 26400
rect 177300 26400 177400 26500
rect 177300 26500 177400 26600
rect 177300 26600 177400 26700
rect 177300 26700 177400 26800
rect 177300 26800 177400 26900
rect 177300 26900 177400 27000
rect 177300 27000 177400 27100
rect 177300 27100 177400 27200
rect 177300 27200 177400 27300
rect 177300 27300 177400 27400
rect 177300 27400 177400 27500
rect 177400 22700 177500 22800
rect 177400 22800 177500 22900
rect 177400 22900 177500 23000
rect 177400 23000 177500 23100
rect 177400 23100 177500 23200
rect 177400 23200 177500 23300
rect 177400 23300 177500 23400
rect 177400 23400 177500 23500
rect 177400 23500 177500 23600
rect 177400 23600 177500 23700
rect 177400 23700 177500 23800
rect 177400 23800 177500 23900
rect 177400 23900 177500 24000
rect 177400 24000 177500 24100
rect 177400 24100 177500 24200
rect 177400 24200 177500 24300
rect 177400 24300 177500 24400
rect 177400 24400 177500 24500
rect 177400 24500 177500 24600
rect 177400 24600 177500 24700
rect 177400 24700 177500 24800
rect 177400 24800 177500 24900
rect 177400 24900 177500 25000
rect 177400 25000 177500 25100
rect 177400 25100 177500 25200
rect 177400 25200 177500 25300
rect 177400 25300 177500 25400
rect 177400 25400 177500 25500
rect 177400 25500 177500 25600
rect 177400 25600 177500 25700
rect 177400 25700 177500 25800
rect 177400 25800 177500 25900
rect 177400 25900 177500 26000
rect 177400 26000 177500 26100
rect 177400 26100 177500 26200
rect 177400 26200 177500 26300
rect 177400 26300 177500 26400
rect 177400 26400 177500 26500
rect 177400 26500 177500 26600
rect 177400 26600 177500 26700
rect 177400 26700 177500 26800
rect 177400 26800 177500 26900
rect 177400 26900 177500 27000
rect 177400 27000 177500 27100
rect 177400 27100 177500 27200
rect 177400 27200 177500 27300
rect 177400 27300 177500 27400
rect 177400 27400 177500 27500
rect 177400 27500 177500 27600
rect 177400 27600 177500 27700
rect 177500 22900 177600 23000
rect 177500 23000 177600 23100
rect 177500 23100 177600 23200
rect 177500 23200 177600 23300
rect 177500 23300 177600 23400
rect 177500 23400 177600 23500
rect 177500 23500 177600 23600
rect 177500 23600 177600 23700
rect 177500 23700 177600 23800
rect 177500 23800 177600 23900
rect 177500 23900 177600 24000
rect 177500 24000 177600 24100
rect 177500 24100 177600 24200
rect 177500 24200 177600 24300
rect 177500 24300 177600 24400
rect 177500 24400 177600 24500
rect 177500 24500 177600 24600
rect 177500 24600 177600 24700
rect 177500 24700 177600 24800
rect 177500 24800 177600 24900
rect 177500 24900 177600 25000
rect 177500 25000 177600 25100
rect 177500 25100 177600 25200
rect 177500 25200 177600 25300
rect 177500 25300 177600 25400
rect 177500 25400 177600 25500
rect 177500 25500 177600 25600
rect 177500 25600 177600 25700
rect 177500 25700 177600 25800
rect 177500 25800 177600 25900
rect 177500 25900 177600 26000
rect 177500 26000 177600 26100
rect 177500 26100 177600 26200
rect 177500 26200 177600 26300
rect 177500 26300 177600 26400
rect 177500 26400 177600 26500
rect 177500 26500 177600 26600
rect 177500 26600 177600 26700
rect 177500 26700 177600 26800
rect 177500 26800 177600 26900
rect 177500 26900 177600 27000
rect 177500 27000 177600 27100
rect 177500 27100 177600 27200
rect 177500 27200 177600 27300
rect 177500 27300 177600 27400
rect 177500 27400 177600 27500
rect 177500 27500 177600 27600
rect 177500 27600 177600 27700
rect 177500 27700 177600 27800
rect 177500 27800 177600 27900
rect 177500 27900 177600 28000
rect 177600 23100 177700 23200
rect 177600 23200 177700 23300
rect 177600 23300 177700 23400
rect 177600 23400 177700 23500
rect 177600 23500 177700 23600
rect 177600 23600 177700 23700
rect 177600 23700 177700 23800
rect 177600 23800 177700 23900
rect 177600 23900 177700 24000
rect 177600 24000 177700 24100
rect 177600 24100 177700 24200
rect 177600 24200 177700 24300
rect 177600 24300 177700 24400
rect 177600 24400 177700 24500
rect 177600 24500 177700 24600
rect 177600 24600 177700 24700
rect 177600 24700 177700 24800
rect 177600 24800 177700 24900
rect 177600 24900 177700 25000
rect 177600 25000 177700 25100
rect 177600 25100 177700 25200
rect 177600 25200 177700 25300
rect 177600 25300 177700 25400
rect 177600 25400 177700 25500
rect 177600 25500 177700 25600
rect 177600 25600 177700 25700
rect 177600 25700 177700 25800
rect 177600 25800 177700 25900
rect 177600 25900 177700 26000
rect 177600 26000 177700 26100
rect 177600 26100 177700 26200
rect 177600 26200 177700 26300
rect 177600 26300 177700 26400
rect 177600 26400 177700 26500
rect 177600 26500 177700 26600
rect 177600 26600 177700 26700
rect 177600 26700 177700 26800
rect 177600 26800 177700 26900
rect 177600 26900 177700 27000
rect 177600 27000 177700 27100
rect 177600 27100 177700 27200
rect 177600 27200 177700 27300
rect 177600 27300 177700 27400
rect 177600 27400 177700 27500
rect 177600 27500 177700 27600
rect 177600 27600 177700 27700
rect 177600 27700 177700 27800
rect 177600 27800 177700 27900
rect 177600 27900 177700 28000
rect 177600 28000 177700 28100
rect 177600 28100 177700 28200
rect 177700 23400 177800 23500
rect 177700 23500 177800 23600
rect 177700 23600 177800 23700
rect 177700 23700 177800 23800
rect 177700 23800 177800 23900
rect 177700 23900 177800 24000
rect 177700 24000 177800 24100
rect 177700 24100 177800 24200
rect 177700 24200 177800 24300
rect 177700 24300 177800 24400
rect 177700 24400 177800 24500
rect 177700 24500 177800 24600
rect 177700 24600 177800 24700
rect 177700 24700 177800 24800
rect 177700 24800 177800 24900
rect 177700 24900 177800 25000
rect 177700 25000 177800 25100
rect 177700 25100 177800 25200
rect 177700 25200 177800 25300
rect 177700 25300 177800 25400
rect 177700 25400 177800 25500
rect 177700 25500 177800 25600
rect 177700 25600 177800 25700
rect 177700 25700 177800 25800
rect 177700 25800 177800 25900
rect 177700 25900 177800 26000
rect 177700 26000 177800 26100
rect 177700 26100 177800 26200
rect 177700 26200 177800 26300
rect 177700 26300 177800 26400
rect 177700 26400 177800 26500
rect 177700 26500 177800 26600
rect 177700 26600 177800 26700
rect 177700 26700 177800 26800
rect 177700 26800 177800 26900
rect 177700 26900 177800 27000
rect 177700 27000 177800 27100
rect 177700 27100 177800 27200
rect 177700 27200 177800 27300
rect 177700 27300 177800 27400
rect 177700 27400 177800 27500
rect 177700 27500 177800 27600
rect 177700 27600 177800 27700
rect 177700 27700 177800 27800
rect 177700 27800 177800 27900
rect 177700 27900 177800 28000
rect 177700 28000 177800 28100
rect 177700 28100 177800 28200
rect 177700 28200 177800 28300
rect 177700 28300 177800 28400
rect 177700 28400 177800 28500
rect 177800 23600 177900 23700
rect 177800 23700 177900 23800
rect 177800 23800 177900 23900
rect 177800 23900 177900 24000
rect 177800 24000 177900 24100
rect 177800 24100 177900 24200
rect 177800 24200 177900 24300
rect 177800 24300 177900 24400
rect 177800 24400 177900 24500
rect 177800 24500 177900 24600
rect 177800 24600 177900 24700
rect 177800 24700 177900 24800
rect 177800 24800 177900 24900
rect 177800 24900 177900 25000
rect 177800 25000 177900 25100
rect 177800 25100 177900 25200
rect 177800 25200 177900 25300
rect 177800 25300 177900 25400
rect 177800 25400 177900 25500
rect 177800 25500 177900 25600
rect 177800 25600 177900 25700
rect 177800 25700 177900 25800
rect 177800 25800 177900 25900
rect 177800 25900 177900 26000
rect 177800 26000 177900 26100
rect 177800 26100 177900 26200
rect 177800 26200 177900 26300
rect 177800 26300 177900 26400
rect 177800 26400 177900 26500
rect 177800 26500 177900 26600
rect 177800 26600 177900 26700
rect 177800 26700 177900 26800
rect 177800 26800 177900 26900
rect 177800 26900 177900 27000
rect 177800 27000 177900 27100
rect 177800 27100 177900 27200
rect 177800 27200 177900 27300
rect 177800 27300 177900 27400
rect 177800 27400 177900 27500
rect 177800 27500 177900 27600
rect 177800 27600 177900 27700
rect 177800 27700 177900 27800
rect 177800 27800 177900 27900
rect 177800 27900 177900 28000
rect 177800 28000 177900 28100
rect 177800 28100 177900 28200
rect 177800 28200 177900 28300
rect 177800 28300 177900 28400
rect 177800 28400 177900 28500
rect 177800 28500 177900 28600
rect 177800 28600 177900 28700
rect 177900 23900 178000 24000
rect 177900 24000 178000 24100
rect 177900 24100 178000 24200
rect 177900 24200 178000 24300
rect 177900 24300 178000 24400
rect 177900 24400 178000 24500
rect 177900 24500 178000 24600
rect 177900 24600 178000 24700
rect 177900 24700 178000 24800
rect 177900 24800 178000 24900
rect 177900 24900 178000 25000
rect 177900 25000 178000 25100
rect 177900 25100 178000 25200
rect 177900 25200 178000 25300
rect 177900 25300 178000 25400
rect 177900 25400 178000 25500
rect 177900 25500 178000 25600
rect 177900 25600 178000 25700
rect 177900 25700 178000 25800
rect 177900 25800 178000 25900
rect 177900 25900 178000 26000
rect 177900 26000 178000 26100
rect 177900 26100 178000 26200
rect 177900 26200 178000 26300
rect 177900 26300 178000 26400
rect 177900 26400 178000 26500
rect 177900 26500 178000 26600
rect 177900 26600 178000 26700
rect 177900 26700 178000 26800
rect 177900 26800 178000 26900
rect 177900 26900 178000 27000
rect 177900 27000 178000 27100
rect 177900 27100 178000 27200
rect 177900 27200 178000 27300
rect 177900 27300 178000 27400
rect 177900 27400 178000 27500
rect 177900 27500 178000 27600
rect 177900 27600 178000 27700
rect 177900 27700 178000 27800
rect 177900 27800 178000 27900
rect 177900 27900 178000 28000
rect 177900 28000 178000 28100
rect 177900 28100 178000 28200
rect 177900 28200 178000 28300
rect 177900 28300 178000 28400
rect 177900 28400 178000 28500
rect 177900 28500 178000 28600
rect 177900 28600 178000 28700
rect 177900 28700 178000 28800
rect 177900 28800 178000 28900
rect 177900 28900 178000 29000
rect 178000 24100 178100 24200
rect 178000 24200 178100 24300
rect 178000 24300 178100 24400
rect 178000 24400 178100 24500
rect 178000 24500 178100 24600
rect 178000 24600 178100 24700
rect 178000 24700 178100 24800
rect 178000 24800 178100 24900
rect 178000 24900 178100 25000
rect 178000 25000 178100 25100
rect 178000 25100 178100 25200
rect 178000 25200 178100 25300
rect 178000 25300 178100 25400
rect 178000 25400 178100 25500
rect 178000 25500 178100 25600
rect 178000 25600 178100 25700
rect 178000 25700 178100 25800
rect 178000 25800 178100 25900
rect 178000 25900 178100 26000
rect 178000 26000 178100 26100
rect 178000 26100 178100 26200
rect 178000 26200 178100 26300
rect 178000 26300 178100 26400
rect 178000 26400 178100 26500
rect 178000 26500 178100 26600
rect 178000 26600 178100 26700
rect 178000 26700 178100 26800
rect 178000 26800 178100 26900
rect 178000 26900 178100 27000
rect 178000 27000 178100 27100
rect 178000 27100 178100 27200
rect 178000 27200 178100 27300
rect 178000 27300 178100 27400
rect 178000 27400 178100 27500
rect 178000 27500 178100 27600
rect 178000 27600 178100 27700
rect 178000 27700 178100 27800
rect 178000 27800 178100 27900
rect 178000 27900 178100 28000
rect 178000 28000 178100 28100
rect 178000 28100 178100 28200
rect 178000 28200 178100 28300
rect 178000 28300 178100 28400
rect 178000 28400 178100 28500
rect 178000 28500 178100 28600
rect 178000 28600 178100 28700
rect 178000 28700 178100 28800
rect 178000 28800 178100 28900
rect 178000 28900 178100 29000
rect 178000 29000 178100 29100
rect 178000 29100 178100 29200
rect 178000 29200 178100 29300
rect 178100 24300 178200 24400
rect 178100 24400 178200 24500
rect 178100 24500 178200 24600
rect 178100 24600 178200 24700
rect 178100 24700 178200 24800
rect 178100 24800 178200 24900
rect 178100 24900 178200 25000
rect 178100 25000 178200 25100
rect 178100 25100 178200 25200
rect 178100 25200 178200 25300
rect 178100 25300 178200 25400
rect 178100 25400 178200 25500
rect 178100 25500 178200 25600
rect 178100 25600 178200 25700
rect 178100 25700 178200 25800
rect 178100 25800 178200 25900
rect 178100 25900 178200 26000
rect 178100 26000 178200 26100
rect 178100 26100 178200 26200
rect 178100 26200 178200 26300
rect 178100 26300 178200 26400
rect 178100 26400 178200 26500
rect 178100 26500 178200 26600
rect 178100 26600 178200 26700
rect 178100 26700 178200 26800
rect 178100 26800 178200 26900
rect 178100 26900 178200 27000
rect 178100 27000 178200 27100
rect 178100 27100 178200 27200
rect 178100 27200 178200 27300
rect 178100 27300 178200 27400
rect 178100 27400 178200 27500
rect 178100 27500 178200 27600
rect 178100 27600 178200 27700
rect 178100 27700 178200 27800
rect 178100 27800 178200 27900
rect 178100 27900 178200 28000
rect 178100 28000 178200 28100
rect 178100 28100 178200 28200
rect 178100 28200 178200 28300
rect 178100 28300 178200 28400
rect 178100 28400 178200 28500
rect 178100 28500 178200 28600
rect 178100 28600 178200 28700
rect 178100 28700 178200 28800
rect 178100 28800 178200 28900
rect 178100 28900 178200 29000
rect 178100 29000 178200 29100
rect 178100 29100 178200 29200
rect 178100 29200 178200 29300
rect 178100 29300 178200 29400
rect 178100 29400 178200 29500
rect 178200 24600 178300 24700
rect 178200 24700 178300 24800
rect 178200 24800 178300 24900
rect 178200 24900 178300 25000
rect 178200 25000 178300 25100
rect 178200 25100 178300 25200
rect 178200 25200 178300 25300
rect 178200 25300 178300 25400
rect 178200 25400 178300 25500
rect 178200 25500 178300 25600
rect 178200 25600 178300 25700
rect 178200 25700 178300 25800
rect 178200 25800 178300 25900
rect 178200 25900 178300 26000
rect 178200 26000 178300 26100
rect 178200 26100 178300 26200
rect 178200 26200 178300 26300
rect 178200 26300 178300 26400
rect 178200 26400 178300 26500
rect 178200 26500 178300 26600
rect 178200 26600 178300 26700
rect 178200 26700 178300 26800
rect 178200 26800 178300 26900
rect 178200 26900 178300 27000
rect 178200 27000 178300 27100
rect 178200 27100 178300 27200
rect 178200 27200 178300 27300
rect 178200 27300 178300 27400
rect 178200 27400 178300 27500
rect 178200 27500 178300 27600
rect 178200 27600 178300 27700
rect 178200 27700 178300 27800
rect 178200 27800 178300 27900
rect 178200 27900 178300 28000
rect 178200 28000 178300 28100
rect 178200 28100 178300 28200
rect 178200 28200 178300 28300
rect 178200 28300 178300 28400
rect 178200 28400 178300 28500
rect 178200 28500 178300 28600
rect 178200 28600 178300 28700
rect 178200 28700 178300 28800
rect 178200 28800 178300 28900
rect 178200 28900 178300 29000
rect 178200 29000 178300 29100
rect 178200 29100 178300 29200
rect 178200 29200 178300 29300
rect 178200 29300 178300 29400
rect 178200 29400 178300 29500
rect 178200 29500 178300 29600
rect 178200 29600 178300 29700
rect 178200 29700 178300 29800
rect 178300 24900 178400 25000
rect 178300 25000 178400 25100
rect 178300 25100 178400 25200
rect 178300 25200 178400 25300
rect 178300 25300 178400 25400
rect 178300 25400 178400 25500
rect 178300 25500 178400 25600
rect 178300 25600 178400 25700
rect 178300 25700 178400 25800
rect 178300 25800 178400 25900
rect 178300 25900 178400 26000
rect 178300 26000 178400 26100
rect 178300 26100 178400 26200
rect 178300 26200 178400 26300
rect 178300 26300 178400 26400
rect 178300 26400 178400 26500
rect 178300 26500 178400 26600
rect 178300 26600 178400 26700
rect 178300 26700 178400 26800
rect 178300 26800 178400 26900
rect 178300 26900 178400 27000
rect 178300 27000 178400 27100
rect 178300 27100 178400 27200
rect 178300 27200 178400 27300
rect 178300 27300 178400 27400
rect 178300 27400 178400 27500
rect 178300 27500 178400 27600
rect 178300 27600 178400 27700
rect 178300 27700 178400 27800
rect 178300 27800 178400 27900
rect 178300 27900 178400 28000
rect 178300 28000 178400 28100
rect 178300 28100 178400 28200
rect 178300 28200 178400 28300
rect 178300 28300 178400 28400
rect 178300 28400 178400 28500
rect 178300 28500 178400 28600
rect 178300 28600 178400 28700
rect 178300 28700 178400 28800
rect 178300 28800 178400 28900
rect 178300 28900 178400 29000
rect 178300 29000 178400 29100
rect 178300 29100 178400 29200
rect 178300 29200 178400 29300
rect 178300 29300 178400 29400
rect 178300 29400 178400 29500
rect 178300 29500 178400 29600
rect 178300 29600 178400 29700
rect 178300 29700 178400 29800
rect 178300 29800 178400 29900
rect 178300 29900 178400 30000
rect 178300 30000 178400 30100
rect 178400 25100 178500 25200
rect 178400 25200 178500 25300
rect 178400 25300 178500 25400
rect 178400 25400 178500 25500
rect 178400 25500 178500 25600
rect 178400 25600 178500 25700
rect 178400 25700 178500 25800
rect 178400 25800 178500 25900
rect 178400 25900 178500 26000
rect 178400 26000 178500 26100
rect 178400 26100 178500 26200
rect 178400 26200 178500 26300
rect 178400 26300 178500 26400
rect 178400 26400 178500 26500
rect 178400 26500 178500 26600
rect 178400 26600 178500 26700
rect 178400 26700 178500 26800
rect 178400 26800 178500 26900
rect 178400 26900 178500 27000
rect 178400 27000 178500 27100
rect 178400 27100 178500 27200
rect 178400 27200 178500 27300
rect 178400 27300 178500 27400
rect 178400 27400 178500 27500
rect 178400 27500 178500 27600
rect 178400 27600 178500 27700
rect 178400 27700 178500 27800
rect 178400 27800 178500 27900
rect 178400 27900 178500 28000
rect 178400 28000 178500 28100
rect 178400 28100 178500 28200
rect 178400 28200 178500 28300
rect 178400 28300 178500 28400
rect 178400 28400 178500 28500
rect 178400 28500 178500 28600
rect 178400 28600 178500 28700
rect 178400 28700 178500 28800
rect 178400 28800 178500 28900
rect 178400 28900 178500 29000
rect 178400 29000 178500 29100
rect 178400 29100 178500 29200
rect 178400 29200 178500 29300
rect 178400 29300 178500 29400
rect 178400 29400 178500 29500
rect 178400 29500 178500 29600
rect 178400 29600 178500 29700
rect 178400 29700 178500 29800
rect 178400 29800 178500 29900
rect 178400 29900 178500 30000
rect 178400 30000 178500 30100
rect 178400 30100 178500 30200
rect 178400 30200 178500 30300
rect 178500 25400 178600 25500
rect 178500 25500 178600 25600
rect 178500 25600 178600 25700
rect 178500 25700 178600 25800
rect 178500 25800 178600 25900
rect 178500 25900 178600 26000
rect 178500 26000 178600 26100
rect 178500 26100 178600 26200
rect 178500 26200 178600 26300
rect 178500 26300 178600 26400
rect 178500 26400 178600 26500
rect 178500 26500 178600 26600
rect 178500 26600 178600 26700
rect 178500 26700 178600 26800
rect 178500 26800 178600 26900
rect 178500 26900 178600 27000
rect 178500 27000 178600 27100
rect 178500 27100 178600 27200
rect 178500 27200 178600 27300
rect 178500 27300 178600 27400
rect 178500 27400 178600 27500
rect 178500 27500 178600 27600
rect 178500 27600 178600 27700
rect 178500 27700 178600 27800
rect 178500 27800 178600 27900
rect 178500 27900 178600 28000
rect 178500 28000 178600 28100
rect 178500 28100 178600 28200
rect 178500 28200 178600 28300
rect 178500 28300 178600 28400
rect 178500 28400 178600 28500
rect 178500 28500 178600 28600
rect 178500 28600 178600 28700
rect 178500 28700 178600 28800
rect 178500 28800 178600 28900
rect 178500 28900 178600 29000
rect 178500 29000 178600 29100
rect 178500 29100 178600 29200
rect 178500 29200 178600 29300
rect 178500 29300 178600 29400
rect 178500 29400 178600 29500
rect 178500 29500 178600 29600
rect 178500 29600 178600 29700
rect 178500 29700 178600 29800
rect 178500 29800 178600 29900
rect 178500 29900 178600 30000
rect 178500 30000 178600 30100
rect 178500 30100 178600 30200
rect 178500 30200 178600 30300
rect 178500 30300 178600 30400
rect 178500 30400 178600 30500
rect 178500 30500 178600 30600
rect 178600 25700 178700 25800
rect 178600 25800 178700 25900
rect 178600 25900 178700 26000
rect 178600 26000 178700 26100
rect 178600 26100 178700 26200
rect 178600 26200 178700 26300
rect 178600 26300 178700 26400
rect 178600 26400 178700 26500
rect 178600 26500 178700 26600
rect 178600 26600 178700 26700
rect 178600 26700 178700 26800
rect 178600 26800 178700 26900
rect 178600 26900 178700 27000
rect 178600 27000 178700 27100
rect 178600 27100 178700 27200
rect 178600 27200 178700 27300
rect 178600 27300 178700 27400
rect 178600 27400 178700 27500
rect 178600 27500 178700 27600
rect 178600 27600 178700 27700
rect 178600 27700 178700 27800
rect 178600 27800 178700 27900
rect 178600 27900 178700 28000
rect 178600 28000 178700 28100
rect 178600 28100 178700 28200
rect 178600 28200 178700 28300
rect 178600 28300 178700 28400
rect 178600 28400 178700 28500
rect 178600 28500 178700 28600
rect 178600 28600 178700 28700
rect 178600 28700 178700 28800
rect 178600 28800 178700 28900
rect 178600 28900 178700 29000
rect 178600 29000 178700 29100
rect 178600 29100 178700 29200
rect 178600 29200 178700 29300
rect 178600 29300 178700 29400
rect 178600 29400 178700 29500
rect 178600 29500 178700 29600
rect 178600 29600 178700 29700
rect 178600 29700 178700 29800
rect 178600 29800 178700 29900
rect 178600 29900 178700 30000
rect 178600 30000 178700 30100
rect 178600 30100 178700 30200
rect 178600 30200 178700 30300
rect 178600 30300 178700 30400
rect 178600 30400 178700 30500
rect 178600 30500 178700 30600
rect 178600 30600 178700 30700
rect 178600 30700 178700 30800
rect 178700 25900 178800 26000
rect 178700 26000 178800 26100
rect 178700 26100 178800 26200
rect 178700 26200 178800 26300
rect 178700 26300 178800 26400
rect 178700 26400 178800 26500
rect 178700 26500 178800 26600
rect 178700 26600 178800 26700
rect 178700 26700 178800 26800
rect 178700 26800 178800 26900
rect 178700 26900 178800 27000
rect 178700 27000 178800 27100
rect 178700 27100 178800 27200
rect 178700 27200 178800 27300
rect 178700 27300 178800 27400
rect 178700 27400 178800 27500
rect 178700 27500 178800 27600
rect 178700 27600 178800 27700
rect 178700 27700 178800 27800
rect 178700 27800 178800 27900
rect 178700 27900 178800 28000
rect 178700 28000 178800 28100
rect 178700 28100 178800 28200
rect 178700 28200 178800 28300
rect 178700 28300 178800 28400
rect 178700 28400 178800 28500
rect 178700 28500 178800 28600
rect 178700 28600 178800 28700
rect 178700 28700 178800 28800
rect 178700 28800 178800 28900
rect 178700 28900 178800 29000
rect 178700 29000 178800 29100
rect 178700 29100 178800 29200
rect 178700 29200 178800 29300
rect 178700 29300 178800 29400
rect 178700 29400 178800 29500
rect 178700 29500 178800 29600
rect 178700 29600 178800 29700
rect 178700 29700 178800 29800
rect 178700 29800 178800 29900
rect 178700 29900 178800 30000
rect 178700 30000 178800 30100
rect 178700 30100 178800 30200
rect 178700 30200 178800 30300
rect 178700 30300 178800 30400
rect 178700 30400 178800 30500
rect 178700 30500 178800 30600
rect 178700 30600 178800 30700
rect 178700 30700 178800 30800
rect 178700 30800 178800 30900
rect 178700 30900 178800 31000
rect 178700 31000 178800 31100
rect 178800 26100 178900 26200
rect 178800 26200 178900 26300
rect 178800 26300 178900 26400
rect 178800 26400 178900 26500
rect 178800 26500 178900 26600
rect 178800 26600 178900 26700
rect 178800 26700 178900 26800
rect 178800 26800 178900 26900
rect 178800 26900 178900 27000
rect 178800 27000 178900 27100
rect 178800 27100 178900 27200
rect 178800 27200 178900 27300
rect 178800 27300 178900 27400
rect 178800 27400 178900 27500
rect 178800 27500 178900 27600
rect 178800 27600 178900 27700
rect 178800 27700 178900 27800
rect 178800 27800 178900 27900
rect 178800 27900 178900 28000
rect 178800 28000 178900 28100
rect 178800 28100 178900 28200
rect 178800 28200 178900 28300
rect 178800 28300 178900 28400
rect 178800 28400 178900 28500
rect 178800 28500 178900 28600
rect 178800 28600 178900 28700
rect 178800 28700 178900 28800
rect 178800 28800 178900 28900
rect 178800 28900 178900 29000
rect 178800 29000 178900 29100
rect 178800 29100 178900 29200
rect 178800 29200 178900 29300
rect 178800 29300 178900 29400
rect 178800 29400 178900 29500
rect 178800 29500 178900 29600
rect 178800 29600 178900 29700
rect 178800 29700 178900 29800
rect 178800 29800 178900 29900
rect 178800 29900 178900 30000
rect 178800 30000 178900 30100
rect 178800 30100 178900 30200
rect 178800 30200 178900 30300
rect 178800 30300 178900 30400
rect 178800 30400 178900 30500
rect 178800 30500 178900 30600
rect 178800 30600 178900 30700
rect 178800 30700 178900 30800
rect 178800 30800 178900 30900
rect 178800 30900 178900 31000
rect 178800 31000 178900 31100
rect 178800 31100 178900 31200
rect 178800 31200 178900 31300
rect 178800 31300 178900 31400
rect 178900 26400 179000 26500
rect 178900 26500 179000 26600
rect 178900 26600 179000 26700
rect 178900 26700 179000 26800
rect 178900 26800 179000 26900
rect 178900 26900 179000 27000
rect 178900 27000 179000 27100
rect 178900 27100 179000 27200
rect 178900 27200 179000 27300
rect 178900 27300 179000 27400
rect 178900 27400 179000 27500
rect 178900 27500 179000 27600
rect 178900 27600 179000 27700
rect 178900 27700 179000 27800
rect 178900 27800 179000 27900
rect 178900 27900 179000 28000
rect 178900 28000 179000 28100
rect 178900 28100 179000 28200
rect 178900 28200 179000 28300
rect 178900 28300 179000 28400
rect 178900 28400 179000 28500
rect 178900 28500 179000 28600
rect 178900 28600 179000 28700
rect 178900 28700 179000 28800
rect 178900 28800 179000 28900
rect 178900 28900 179000 29000
rect 178900 29000 179000 29100
rect 178900 29100 179000 29200
rect 178900 29200 179000 29300
rect 178900 29300 179000 29400
rect 178900 29400 179000 29500
rect 178900 29500 179000 29600
rect 178900 29600 179000 29700
rect 178900 29700 179000 29800
rect 178900 29800 179000 29900
rect 178900 29900 179000 30000
rect 178900 30000 179000 30100
rect 178900 30100 179000 30200
rect 178900 30200 179000 30300
rect 178900 30300 179000 30400
rect 178900 30400 179000 30500
rect 178900 30500 179000 30600
rect 178900 30600 179000 30700
rect 178900 30700 179000 30800
rect 178900 30800 179000 30900
rect 178900 30900 179000 31000
rect 178900 31000 179000 31100
rect 178900 31100 179000 31200
rect 178900 31200 179000 31300
rect 178900 31300 179000 31400
rect 178900 31400 179000 31500
rect 178900 31500 179000 31600
rect 179000 26600 179100 26700
rect 179000 26700 179100 26800
rect 179000 26800 179100 26900
rect 179000 26900 179100 27000
rect 179000 27000 179100 27100
rect 179000 27100 179100 27200
rect 179000 27200 179100 27300
rect 179000 27300 179100 27400
rect 179000 27400 179100 27500
rect 179000 27500 179100 27600
rect 179000 27600 179100 27700
rect 179000 27700 179100 27800
rect 179000 27800 179100 27900
rect 179000 27900 179100 28000
rect 179000 28000 179100 28100
rect 179000 28100 179100 28200
rect 179000 28200 179100 28300
rect 179000 28300 179100 28400
rect 179000 28400 179100 28500
rect 179000 28500 179100 28600
rect 179000 28600 179100 28700
rect 179000 28700 179100 28800
rect 179000 28800 179100 28900
rect 179000 28900 179100 29000
rect 179000 29000 179100 29100
rect 179000 29100 179100 29200
rect 179000 29200 179100 29300
rect 179000 29300 179100 29400
rect 179000 29400 179100 29500
rect 179000 29500 179100 29600
rect 179000 29600 179100 29700
rect 179000 29700 179100 29800
rect 179000 29800 179100 29900
rect 179000 29900 179100 30000
rect 179000 30000 179100 30100
rect 179000 30100 179100 30200
rect 179000 30200 179100 30300
rect 179000 30300 179100 30400
rect 179000 30400 179100 30500
rect 179000 30500 179100 30600
rect 179000 30600 179100 30700
rect 179000 30700 179100 30800
rect 179000 30800 179100 30900
rect 179000 30900 179100 31000
rect 179000 31000 179100 31100
rect 179000 31100 179100 31200
rect 179000 31200 179100 31300
rect 179000 31300 179100 31400
rect 179000 31400 179100 31500
rect 179000 31500 179100 31600
rect 179000 31600 179100 31700
rect 179000 31700 179100 31800
rect 179000 31800 179100 31900
rect 179100 26900 179200 27000
rect 179100 27000 179200 27100
rect 179100 27100 179200 27200
rect 179100 27200 179200 27300
rect 179100 27300 179200 27400
rect 179100 27400 179200 27500
rect 179100 27500 179200 27600
rect 179100 27600 179200 27700
rect 179100 27700 179200 27800
rect 179100 27800 179200 27900
rect 179100 27900 179200 28000
rect 179100 28000 179200 28100
rect 179100 28100 179200 28200
rect 179100 28200 179200 28300
rect 179100 28300 179200 28400
rect 179100 28400 179200 28500
rect 179100 28500 179200 28600
rect 179100 28600 179200 28700
rect 179100 28700 179200 28800
rect 179100 28800 179200 28900
rect 179100 28900 179200 29000
rect 179100 29000 179200 29100
rect 179100 29100 179200 29200
rect 179100 29200 179200 29300
rect 179100 29300 179200 29400
rect 179100 29400 179200 29500
rect 179100 29500 179200 29600
rect 179100 29600 179200 29700
rect 179100 29700 179200 29800
rect 179100 29800 179200 29900
rect 179100 29900 179200 30000
rect 179100 30000 179200 30100
rect 179100 30100 179200 30200
rect 179100 30200 179200 30300
rect 179100 30300 179200 30400
rect 179100 30400 179200 30500
rect 179100 30500 179200 30600
rect 179100 30600 179200 30700
rect 179100 30700 179200 30800
rect 179100 30800 179200 30900
rect 179100 30900 179200 31000
rect 179100 31000 179200 31100
rect 179100 31100 179200 31200
rect 179100 31200 179200 31300
rect 179100 31300 179200 31400
rect 179100 31400 179200 31500
rect 179100 31500 179200 31600
rect 179100 31600 179200 31700
rect 179100 31700 179200 31800
rect 179100 31800 179200 31900
rect 179100 31900 179200 32000
rect 179100 32000 179200 32100
rect 179100 32100 179200 32200
rect 179200 27100 179300 27200
rect 179200 27200 179300 27300
rect 179200 27300 179300 27400
rect 179200 27400 179300 27500
rect 179200 27500 179300 27600
rect 179200 27600 179300 27700
rect 179200 27700 179300 27800
rect 179200 27800 179300 27900
rect 179200 27900 179300 28000
rect 179200 28000 179300 28100
rect 179200 28100 179300 28200
rect 179200 28200 179300 28300
rect 179200 28300 179300 28400
rect 179200 28400 179300 28500
rect 179200 28500 179300 28600
rect 179200 28600 179300 28700
rect 179200 28700 179300 28800
rect 179200 28800 179300 28900
rect 179200 28900 179300 29000
rect 179200 29000 179300 29100
rect 179200 29100 179300 29200
rect 179200 29200 179300 29300
rect 179200 29300 179300 29400
rect 179200 29400 179300 29500
rect 179200 29500 179300 29600
rect 179200 29600 179300 29700
rect 179200 29700 179300 29800
rect 179200 29800 179300 29900
rect 179200 29900 179300 30000
rect 179200 30000 179300 30100
rect 179200 30100 179300 30200
rect 179200 30200 179300 30300
rect 179200 30300 179300 30400
rect 179200 30400 179300 30500
rect 179200 30500 179300 30600
rect 179200 30600 179300 30700
rect 179200 30700 179300 30800
rect 179200 30800 179300 30900
rect 179200 30900 179300 31000
rect 179200 31000 179300 31100
rect 179200 31100 179300 31200
rect 179200 31200 179300 31300
rect 179200 31300 179300 31400
rect 179200 31400 179300 31500
rect 179200 31500 179300 31600
rect 179200 31600 179300 31700
rect 179200 31700 179300 31800
rect 179200 31800 179300 31900
rect 179200 31900 179300 32000
rect 179200 32000 179300 32100
rect 179200 32100 179300 32200
rect 179200 32200 179300 32300
rect 179200 32300 179300 32400
rect 179200 32400 179300 32500
rect 179300 27400 179400 27500
rect 179300 27500 179400 27600
rect 179300 27600 179400 27700
rect 179300 27700 179400 27800
rect 179300 27800 179400 27900
rect 179300 27900 179400 28000
rect 179300 28000 179400 28100
rect 179300 28100 179400 28200
rect 179300 28200 179400 28300
rect 179300 28300 179400 28400
rect 179300 28400 179400 28500
rect 179300 28500 179400 28600
rect 179300 28600 179400 28700
rect 179300 28700 179400 28800
rect 179300 28800 179400 28900
rect 179300 28900 179400 29000
rect 179300 29000 179400 29100
rect 179300 29100 179400 29200
rect 179300 29200 179400 29300
rect 179300 29300 179400 29400
rect 179300 29400 179400 29500
rect 179300 29500 179400 29600
rect 179300 29600 179400 29700
rect 179300 29700 179400 29800
rect 179300 29800 179400 29900
rect 179300 29900 179400 30000
rect 179300 30000 179400 30100
rect 179300 30100 179400 30200
rect 179300 30200 179400 30300
rect 179300 30300 179400 30400
rect 179300 30400 179400 30500
rect 179300 30500 179400 30600
rect 179300 30600 179400 30700
rect 179300 30700 179400 30800
rect 179300 30800 179400 30900
rect 179300 30900 179400 31000
rect 179300 31000 179400 31100
rect 179300 31100 179400 31200
rect 179300 31200 179400 31300
rect 179300 31300 179400 31400
rect 179300 31400 179400 31500
rect 179300 31500 179400 31600
rect 179300 31600 179400 31700
rect 179300 31700 179400 31800
rect 179300 31800 179400 31900
rect 179300 31900 179400 32000
rect 179300 32000 179400 32100
rect 179300 32100 179400 32200
rect 179300 32200 179400 32300
rect 179300 32300 179400 32400
rect 179300 32400 179400 32500
rect 179300 32500 179400 32600
rect 179300 32600 179400 32700
rect 179400 27600 179500 27700
rect 179400 27700 179500 27800
rect 179400 27800 179500 27900
rect 179400 27900 179500 28000
rect 179400 28000 179500 28100
rect 179400 28100 179500 28200
rect 179400 28200 179500 28300
rect 179400 28300 179500 28400
rect 179400 28400 179500 28500
rect 179400 28500 179500 28600
rect 179400 28600 179500 28700
rect 179400 28700 179500 28800
rect 179400 28800 179500 28900
rect 179400 28900 179500 29000
rect 179400 29000 179500 29100
rect 179400 29100 179500 29200
rect 179400 29200 179500 29300
rect 179400 29300 179500 29400
rect 179400 29400 179500 29500
rect 179400 29500 179500 29600
rect 179400 29600 179500 29700
rect 179400 29700 179500 29800
rect 179400 29800 179500 29900
rect 179400 29900 179500 30000
rect 179400 30000 179500 30100
rect 179400 30100 179500 30200
rect 179400 30200 179500 30300
rect 179400 30300 179500 30400
rect 179400 30400 179500 30500
rect 179400 30500 179500 30600
rect 179400 30600 179500 30700
rect 179400 30700 179500 30800
rect 179400 30800 179500 30900
rect 179400 30900 179500 31000
rect 179400 31000 179500 31100
rect 179400 31100 179500 31200
rect 179400 31200 179500 31300
rect 179400 31300 179500 31400
rect 179400 31400 179500 31500
rect 179400 31500 179500 31600
rect 179400 31600 179500 31700
rect 179400 31700 179500 31800
rect 179400 31800 179500 31900
rect 179400 31900 179500 32000
rect 179400 32000 179500 32100
rect 179400 32100 179500 32200
rect 179400 32200 179500 32300
rect 179400 32300 179500 32400
rect 179400 32400 179500 32500
rect 179400 32500 179500 32600
rect 179400 32600 179500 32700
rect 179400 32700 179500 32800
rect 179400 32800 179500 32900
rect 179400 32900 179500 33000
rect 179500 27900 179600 28000
rect 179500 28000 179600 28100
rect 179500 28100 179600 28200
rect 179500 28200 179600 28300
rect 179500 28300 179600 28400
rect 179500 28400 179600 28500
rect 179500 28500 179600 28600
rect 179500 28600 179600 28700
rect 179500 28700 179600 28800
rect 179500 28800 179600 28900
rect 179500 28900 179600 29000
rect 179500 29000 179600 29100
rect 179500 29100 179600 29200
rect 179500 29200 179600 29300
rect 179500 29300 179600 29400
rect 179500 29400 179600 29500
rect 179500 29500 179600 29600
rect 179500 29600 179600 29700
rect 179500 29700 179600 29800
rect 179500 29800 179600 29900
rect 179500 29900 179600 30000
rect 179500 30000 179600 30100
rect 179500 30100 179600 30200
rect 179500 30200 179600 30300
rect 179500 30300 179600 30400
rect 179500 30400 179600 30500
rect 179500 30500 179600 30600
rect 179500 30600 179600 30700
rect 179500 30700 179600 30800
rect 179500 30800 179600 30900
rect 179500 30900 179600 31000
rect 179500 31000 179600 31100
rect 179500 31100 179600 31200
rect 179500 31200 179600 31300
rect 179500 31300 179600 31400
rect 179500 31400 179600 31500
rect 179500 31500 179600 31600
rect 179500 31600 179600 31700
rect 179500 31700 179600 31800
rect 179500 31800 179600 31900
rect 179500 31900 179600 32000
rect 179500 32000 179600 32100
rect 179500 32100 179600 32200
rect 179500 32200 179600 32300
rect 179500 32300 179600 32400
rect 179500 32400 179600 32500
rect 179500 32500 179600 32600
rect 179500 32600 179600 32700
rect 179500 32700 179600 32800
rect 179500 32800 179600 32900
rect 179500 32900 179600 33000
rect 179500 33000 179600 33100
rect 179500 33100 179600 33200
rect 179500 33200 179600 33300
rect 179600 28100 179700 28200
rect 179600 28200 179700 28300
rect 179600 28300 179700 28400
rect 179600 28400 179700 28500
rect 179600 28500 179700 28600
rect 179600 28600 179700 28700
rect 179600 28700 179700 28800
rect 179600 28800 179700 28900
rect 179600 28900 179700 29000
rect 179600 29000 179700 29100
rect 179600 29100 179700 29200
rect 179600 29200 179700 29300
rect 179600 29300 179700 29400
rect 179600 29400 179700 29500
rect 179600 29500 179700 29600
rect 179600 29600 179700 29700
rect 179600 29700 179700 29800
rect 179600 29800 179700 29900
rect 179600 29900 179700 30000
rect 179600 30000 179700 30100
rect 179600 30100 179700 30200
rect 179600 30200 179700 30300
rect 179600 30300 179700 30400
rect 179600 30400 179700 30500
rect 179600 30500 179700 30600
rect 179600 30600 179700 30700
rect 179600 30700 179700 30800
rect 179600 30800 179700 30900
rect 179600 30900 179700 31000
rect 179600 31000 179700 31100
rect 179600 31100 179700 31200
rect 179600 31200 179700 31300
rect 179600 31300 179700 31400
rect 179600 31400 179700 31500
rect 179600 31500 179700 31600
rect 179600 31600 179700 31700
rect 179600 31700 179700 31800
rect 179600 31800 179700 31900
rect 179600 31900 179700 32000
rect 179600 32000 179700 32100
rect 179600 32100 179700 32200
rect 179600 32200 179700 32300
rect 179600 32300 179700 32400
rect 179600 32400 179700 32500
rect 179600 32500 179700 32600
rect 179600 32600 179700 32700
rect 179600 32700 179700 32800
rect 179600 32800 179700 32900
rect 179600 32900 179700 33000
rect 179600 33000 179700 33100
rect 179600 33100 179700 33200
rect 179600 33200 179700 33300
rect 179600 33300 179700 33400
rect 179600 33400 179700 33500
rect 179700 28300 179800 28400
rect 179700 28400 179800 28500
rect 179700 28500 179800 28600
rect 179700 28600 179800 28700
rect 179700 28700 179800 28800
rect 179700 28800 179800 28900
rect 179700 28900 179800 29000
rect 179700 29000 179800 29100
rect 179700 29100 179800 29200
rect 179700 29200 179800 29300
rect 179700 29300 179800 29400
rect 179700 29400 179800 29500
rect 179700 29500 179800 29600
rect 179700 29600 179800 29700
rect 179700 29700 179800 29800
rect 179700 29800 179800 29900
rect 179700 29900 179800 30000
rect 179700 30000 179800 30100
rect 179700 30100 179800 30200
rect 179700 30200 179800 30300
rect 179700 30300 179800 30400
rect 179700 30400 179800 30500
rect 179700 30500 179800 30600
rect 179700 30600 179800 30700
rect 179700 30700 179800 30800
rect 179700 30800 179800 30900
rect 179700 30900 179800 31000
rect 179700 31000 179800 31100
rect 179700 31100 179800 31200
rect 179700 31200 179800 31300
rect 179700 31300 179800 31400
rect 179700 31400 179800 31500
rect 179700 31500 179800 31600
rect 179700 31600 179800 31700
rect 179700 31700 179800 31800
rect 179700 31800 179800 31900
rect 179700 31900 179800 32000
rect 179700 32000 179800 32100
rect 179700 32100 179800 32200
rect 179700 32200 179800 32300
rect 179700 32300 179800 32400
rect 179700 32400 179800 32500
rect 179700 32500 179800 32600
rect 179700 32600 179800 32700
rect 179700 32700 179800 32800
rect 179700 32800 179800 32900
rect 179700 32900 179800 33000
rect 179700 33000 179800 33100
rect 179700 33100 179800 33200
rect 179700 33200 179800 33300
rect 179700 33300 179800 33400
rect 179700 33400 179800 33500
rect 179700 33500 179800 33600
rect 179700 33600 179800 33700
rect 179700 33700 179800 33800
rect 179800 28600 179900 28700
rect 179800 28700 179900 28800
rect 179800 28800 179900 28900
rect 179800 28900 179900 29000
rect 179800 29000 179900 29100
rect 179800 29100 179900 29200
rect 179800 29200 179900 29300
rect 179800 29300 179900 29400
rect 179800 29400 179900 29500
rect 179800 29500 179900 29600
rect 179800 29600 179900 29700
rect 179800 29700 179900 29800
rect 179800 29800 179900 29900
rect 179800 29900 179900 30000
rect 179800 30000 179900 30100
rect 179800 30100 179900 30200
rect 179800 30200 179900 30300
rect 179800 30300 179900 30400
rect 179800 30400 179900 30500
rect 179800 30500 179900 30600
rect 179800 30600 179900 30700
rect 179800 30700 179900 30800
rect 179800 30800 179900 30900
rect 179800 30900 179900 31000
rect 179800 31000 179900 31100
rect 179800 31100 179900 31200
rect 179800 31200 179900 31300
rect 179800 31300 179900 31400
rect 179800 31400 179900 31500
rect 179800 31500 179900 31600
rect 179800 31600 179900 31700
rect 179800 31700 179900 31800
rect 179800 31800 179900 31900
rect 179800 31900 179900 32000
rect 179800 32000 179900 32100
rect 179800 32100 179900 32200
rect 179800 32200 179900 32300
rect 179800 32300 179900 32400
rect 179800 32400 179900 32500
rect 179800 32500 179900 32600
rect 179800 32600 179900 32700
rect 179800 32700 179900 32800
rect 179800 32800 179900 32900
rect 179800 32900 179900 33000
rect 179800 33000 179900 33100
rect 179800 33100 179900 33200
rect 179800 33200 179900 33300
rect 179800 33300 179900 33400
rect 179800 33400 179900 33500
rect 179800 33500 179900 33600
rect 179800 33600 179900 33700
rect 179800 33700 179900 33800
rect 179800 33800 179900 33900
rect 179800 33900 179900 34000
rect 179800 34000 179900 34100
rect 179800 34100 179900 34200
rect 179900 28800 180000 28900
rect 179900 28900 180000 29000
rect 179900 29000 180000 29100
rect 179900 29100 180000 29200
rect 179900 29200 180000 29300
rect 179900 29300 180000 29400
rect 179900 29400 180000 29500
rect 179900 29500 180000 29600
rect 179900 29600 180000 29700
rect 179900 29700 180000 29800
rect 179900 29800 180000 29900
rect 179900 29900 180000 30000
rect 179900 30000 180000 30100
rect 179900 30100 180000 30200
rect 179900 30200 180000 30300
rect 179900 30300 180000 30400
rect 179900 30400 180000 30500
rect 179900 30500 180000 30600
rect 179900 30600 180000 30700
rect 179900 30700 180000 30800
rect 179900 30800 180000 30900
rect 179900 30900 180000 31000
rect 179900 31000 180000 31100
rect 179900 31100 180000 31200
rect 179900 31200 180000 31300
rect 179900 31300 180000 31400
rect 179900 31400 180000 31500
rect 179900 31500 180000 31600
rect 179900 31600 180000 31700
rect 179900 31700 180000 31800
rect 179900 31800 180000 31900
rect 179900 31900 180000 32000
rect 179900 32000 180000 32100
rect 179900 32100 180000 32200
rect 179900 32200 180000 32300
rect 179900 32300 180000 32400
rect 179900 32400 180000 32500
rect 179900 32500 180000 32600
rect 179900 32600 180000 32700
rect 179900 32700 180000 32800
rect 179900 32800 180000 32900
rect 179900 32900 180000 33000
rect 179900 33000 180000 33100
rect 179900 33100 180000 33200
rect 179900 33200 180000 33300
rect 179900 33300 180000 33400
rect 179900 33400 180000 33500
rect 179900 33500 180000 33600
rect 179900 33600 180000 33700
rect 179900 33700 180000 33800
rect 179900 33800 180000 33900
rect 179900 33900 180000 34000
rect 179900 34000 180000 34100
rect 179900 34100 180000 34200
rect 179900 34200 180000 34300
rect 179900 34300 180000 34400
rect 179900 34400 180000 34500
rect 180000 29100 180100 29200
rect 180000 29200 180100 29300
rect 180000 29300 180100 29400
rect 180000 29400 180100 29500
rect 180000 29500 180100 29600
rect 180000 29600 180100 29700
rect 180000 29700 180100 29800
rect 180000 29800 180100 29900
rect 180000 29900 180100 30000
rect 180000 30000 180100 30100
rect 180000 30100 180100 30200
rect 180000 30200 180100 30300
rect 180000 30300 180100 30400
rect 180000 30400 180100 30500
rect 180000 30500 180100 30600
rect 180000 30600 180100 30700
rect 180000 30700 180100 30800
rect 180000 30800 180100 30900
rect 180000 30900 180100 31000
rect 180000 31000 180100 31100
rect 180000 31100 180100 31200
rect 180000 31200 180100 31300
rect 180000 31300 180100 31400
rect 180000 31400 180100 31500
rect 180000 31500 180100 31600
rect 180000 31600 180100 31700
rect 180000 31700 180100 31800
rect 180000 31800 180100 31900
rect 180000 31900 180100 32000
rect 180000 32000 180100 32100
rect 180000 32100 180100 32200
rect 180000 32200 180100 32300
rect 180000 32300 180100 32400
rect 180000 32400 180100 32500
rect 180000 32500 180100 32600
rect 180000 32600 180100 32700
rect 180000 32700 180100 32800
rect 180000 32800 180100 32900
rect 180000 32900 180100 33000
rect 180000 33000 180100 33100
rect 180000 33100 180100 33200
rect 180000 33200 180100 33300
rect 180000 33300 180100 33400
rect 180000 33400 180100 33500
rect 180000 33500 180100 33600
rect 180000 33600 180100 33700
rect 180000 33700 180100 33800
rect 180000 33800 180100 33900
rect 180000 33900 180100 34000
rect 180000 34000 180100 34100
rect 180000 34100 180100 34200
rect 180000 34200 180100 34300
rect 180000 34300 180100 34400
rect 180000 34400 180100 34500
rect 180000 34500 180100 34600
rect 180000 34600 180100 34700
rect 180000 34700 180100 34800
rect 180000 34800 180100 34900
rect 180100 29300 180200 29400
rect 180100 29400 180200 29500
rect 180100 29500 180200 29600
rect 180100 29600 180200 29700
rect 180100 29700 180200 29800
rect 180100 29800 180200 29900
rect 180100 29900 180200 30000
rect 180100 30000 180200 30100
rect 180100 30100 180200 30200
rect 180100 30200 180200 30300
rect 180100 30300 180200 30400
rect 180100 30400 180200 30500
rect 180100 30500 180200 30600
rect 180100 30600 180200 30700
rect 180100 30700 180200 30800
rect 180100 30800 180200 30900
rect 180100 30900 180200 31000
rect 180100 31000 180200 31100
rect 180100 31100 180200 31200
rect 180100 31200 180200 31300
rect 180100 31300 180200 31400
rect 180100 31400 180200 31500
rect 180100 31500 180200 31600
rect 180100 31600 180200 31700
rect 180100 31700 180200 31800
rect 180100 31800 180200 31900
rect 180100 31900 180200 32000
rect 180100 32000 180200 32100
rect 180100 32100 180200 32200
rect 180100 32200 180200 32300
rect 180100 32300 180200 32400
rect 180100 32400 180200 32500
rect 180100 32500 180200 32600
rect 180100 32600 180200 32700
rect 180100 32700 180200 32800
rect 180100 32800 180200 32900
rect 180100 32900 180200 33000
rect 180100 33000 180200 33100
rect 180100 33100 180200 33200
rect 180100 33200 180200 33300
rect 180100 33300 180200 33400
rect 180100 33400 180200 33500
rect 180100 33500 180200 33600
rect 180100 33600 180200 33700
rect 180100 33700 180200 33800
rect 180100 33800 180200 33900
rect 180100 33900 180200 34000
rect 180100 34000 180200 34100
rect 180100 34100 180200 34200
rect 180100 34200 180200 34300
rect 180100 34300 180200 34400
rect 180100 34400 180200 34500
rect 180100 34500 180200 34600
rect 180100 34600 180200 34700
rect 180100 34700 180200 34800
rect 180100 34800 180200 34900
rect 180100 34900 180200 35000
rect 180100 35000 180200 35100
rect 180100 35100 180200 35200
rect 180100 35200 180200 35300
rect 180200 29600 180300 29700
rect 180200 29700 180300 29800
rect 180200 29800 180300 29900
rect 180200 29900 180300 30000
rect 180200 30000 180300 30100
rect 180200 30100 180300 30200
rect 180200 30200 180300 30300
rect 180200 30300 180300 30400
rect 180200 30400 180300 30500
rect 180200 30500 180300 30600
rect 180200 30600 180300 30700
rect 180200 30700 180300 30800
rect 180200 30800 180300 30900
rect 180200 30900 180300 31000
rect 180200 31000 180300 31100
rect 180200 31100 180300 31200
rect 180200 31200 180300 31300
rect 180200 31300 180300 31400
rect 180200 31400 180300 31500
rect 180200 31500 180300 31600
rect 180200 31600 180300 31700
rect 180200 31700 180300 31800
rect 180200 31800 180300 31900
rect 180200 31900 180300 32000
rect 180200 32000 180300 32100
rect 180200 32100 180300 32200
rect 180200 32200 180300 32300
rect 180200 32300 180300 32400
rect 180200 32400 180300 32500
rect 180200 32500 180300 32600
rect 180200 32600 180300 32700
rect 180200 32700 180300 32800
rect 180200 32800 180300 32900
rect 180200 32900 180300 33000
rect 180200 33000 180300 33100
rect 180200 33100 180300 33200
rect 180200 33200 180300 33300
rect 180200 33300 180300 33400
rect 180200 33400 180300 33500
rect 180200 33500 180300 33600
rect 180200 33600 180300 33700
rect 180200 33700 180300 33800
rect 180200 33800 180300 33900
rect 180200 33900 180300 34000
rect 180200 34000 180300 34100
rect 180200 34100 180300 34200
rect 180200 34200 180300 34300
rect 180200 34300 180300 34400
rect 180200 34400 180300 34500
rect 180200 34500 180300 34600
rect 180200 34600 180300 34700
rect 180200 34700 180300 34800
rect 180200 34800 180300 34900
rect 180200 34900 180300 35000
rect 180200 35000 180300 35100
rect 180200 35100 180300 35200
rect 180200 35200 180300 35300
rect 180200 35300 180300 35400
rect 180200 35400 180300 35500
rect 180200 35500 180300 35600
rect 180200 35600 180300 35700
rect 180300 29800 180400 29900
rect 180300 29900 180400 30000
rect 180300 30000 180400 30100
rect 180300 30100 180400 30200
rect 180300 30200 180400 30300
rect 180300 30300 180400 30400
rect 180300 30400 180400 30500
rect 180300 30500 180400 30600
rect 180300 30600 180400 30700
rect 180300 30700 180400 30800
rect 180300 30800 180400 30900
rect 180300 30900 180400 31000
rect 180300 31000 180400 31100
rect 180300 31100 180400 31200
rect 180300 31200 180400 31300
rect 180300 31300 180400 31400
rect 180300 31400 180400 31500
rect 180300 31500 180400 31600
rect 180300 31600 180400 31700
rect 180300 31700 180400 31800
rect 180300 31800 180400 31900
rect 180300 31900 180400 32000
rect 180300 32000 180400 32100
rect 180300 32100 180400 32200
rect 180300 32200 180400 32300
rect 180300 32300 180400 32400
rect 180300 32400 180400 32500
rect 180300 32500 180400 32600
rect 180300 32600 180400 32700
rect 180300 32700 180400 32800
rect 180300 32800 180400 32900
rect 180300 32900 180400 33000
rect 180300 33000 180400 33100
rect 180300 33100 180400 33200
rect 180300 33200 180400 33300
rect 180300 33300 180400 33400
rect 180300 33400 180400 33500
rect 180300 33500 180400 33600
rect 180300 33600 180400 33700
rect 180300 33700 180400 33800
rect 180300 33800 180400 33900
rect 180300 33900 180400 34000
rect 180300 34000 180400 34100
rect 180300 34100 180400 34200
rect 180300 34200 180400 34300
rect 180300 34300 180400 34400
rect 180300 34400 180400 34500
rect 180300 34500 180400 34600
rect 180300 34600 180400 34700
rect 180300 34700 180400 34800
rect 180300 34800 180400 34900
rect 180300 34900 180400 35000
rect 180300 35000 180400 35100
rect 180300 35100 180400 35200
rect 180300 35200 180400 35300
rect 180300 35300 180400 35400
rect 180300 35400 180400 35500
rect 180300 35500 180400 35600
rect 180300 35600 180400 35700
rect 180300 35700 180400 35800
rect 180300 35800 180400 35900
rect 180300 35900 180400 36000
rect 180300 36000 180400 36100
rect 180400 30000 180500 30100
rect 180400 30100 180500 30200
rect 180400 30200 180500 30300
rect 180400 30300 180500 30400
rect 180400 30400 180500 30500
rect 180400 30500 180500 30600
rect 180400 30600 180500 30700
rect 180400 30700 180500 30800
rect 180400 30800 180500 30900
rect 180400 30900 180500 31000
rect 180400 31000 180500 31100
rect 180400 31100 180500 31200
rect 180400 31200 180500 31300
rect 180400 31300 180500 31400
rect 180400 31400 180500 31500
rect 180400 31500 180500 31600
rect 180400 31600 180500 31700
rect 180400 31700 180500 31800
rect 180400 31800 180500 31900
rect 180400 31900 180500 32000
rect 180400 32000 180500 32100
rect 180400 32100 180500 32200
rect 180400 32200 180500 32300
rect 180400 32300 180500 32400
rect 180400 32400 180500 32500
rect 180400 32500 180500 32600
rect 180400 32600 180500 32700
rect 180400 32700 180500 32800
rect 180400 32800 180500 32900
rect 180400 32900 180500 33000
rect 180400 33000 180500 33100
rect 180400 33100 180500 33200
rect 180400 33200 180500 33300
rect 180400 33300 180500 33400
rect 180400 33400 180500 33500
rect 180400 33500 180500 33600
rect 180400 33600 180500 33700
rect 180400 33700 180500 33800
rect 180400 33800 180500 33900
rect 180400 33900 180500 34000
rect 180400 34000 180500 34100
rect 180400 34100 180500 34200
rect 180400 34200 180500 34300
rect 180400 34300 180500 34400
rect 180400 34400 180500 34500
rect 180400 34500 180500 34600
rect 180400 34600 180500 34700
rect 180400 34700 180500 34800
rect 180400 34800 180500 34900
rect 180400 34900 180500 35000
rect 180400 35000 180500 35100
rect 180400 35100 180500 35200
rect 180400 35200 180500 35300
rect 180400 35300 180500 35400
rect 180400 35400 180500 35500
rect 180400 35500 180500 35600
rect 180400 35600 180500 35700
rect 180400 35700 180500 35800
rect 180400 35800 180500 35900
rect 180400 35900 180500 36000
rect 180400 36000 180500 36100
rect 180400 36100 180500 36200
rect 180400 36200 180500 36300
rect 180400 36300 180500 36400
rect 180500 30300 180600 30400
rect 180500 30400 180600 30500
rect 180500 30500 180600 30600
rect 180500 30600 180600 30700
rect 180500 30700 180600 30800
rect 180500 30800 180600 30900
rect 180500 30900 180600 31000
rect 180500 31000 180600 31100
rect 180500 31100 180600 31200
rect 180500 31200 180600 31300
rect 180500 31300 180600 31400
rect 180500 31400 180600 31500
rect 180500 31500 180600 31600
rect 180500 31600 180600 31700
rect 180500 31700 180600 31800
rect 180500 31800 180600 31900
rect 180500 31900 180600 32000
rect 180500 32000 180600 32100
rect 180500 32100 180600 32200
rect 180500 32200 180600 32300
rect 180500 32300 180600 32400
rect 180500 32400 180600 32500
rect 180500 32500 180600 32600
rect 180500 32600 180600 32700
rect 180500 32700 180600 32800
rect 180500 32800 180600 32900
rect 180500 32900 180600 33000
rect 180500 33000 180600 33100
rect 180500 33100 180600 33200
rect 180500 33200 180600 33300
rect 180500 33300 180600 33400
rect 180500 33400 180600 33500
rect 180500 33500 180600 33600
rect 180500 33600 180600 33700
rect 180500 33700 180600 33800
rect 180500 33800 180600 33900
rect 180500 33900 180600 34000
rect 180500 34000 180600 34100
rect 180500 34100 180600 34200
rect 180500 34200 180600 34300
rect 180500 34300 180600 34400
rect 180500 34400 180600 34500
rect 180500 34500 180600 34600
rect 180500 34600 180600 34700
rect 180500 34700 180600 34800
rect 180500 34800 180600 34900
rect 180500 34900 180600 35000
rect 180500 35000 180600 35100
rect 180500 35100 180600 35200
rect 180500 35200 180600 35300
rect 180500 35300 180600 35400
rect 180500 35400 180600 35500
rect 180500 35500 180600 35600
rect 180500 35600 180600 35700
rect 180500 35700 180600 35800
rect 180500 35800 180600 35900
rect 180500 35900 180600 36000
rect 180500 36000 180600 36100
rect 180500 36100 180600 36200
rect 180500 36200 180600 36300
rect 180500 36300 180600 36400
rect 180500 36400 180600 36500
rect 180500 36500 180600 36600
rect 180500 36600 180600 36700
rect 180600 30500 180700 30600
rect 180600 30600 180700 30700
rect 180600 30700 180700 30800
rect 180600 30800 180700 30900
rect 180600 30900 180700 31000
rect 180600 31000 180700 31100
rect 180600 31100 180700 31200
rect 180600 31200 180700 31300
rect 180600 31300 180700 31400
rect 180600 31400 180700 31500
rect 180600 31500 180700 31600
rect 180600 31600 180700 31700
rect 180600 31700 180700 31800
rect 180600 31800 180700 31900
rect 180600 31900 180700 32000
rect 180600 32000 180700 32100
rect 180600 32100 180700 32200
rect 180600 32200 180700 32300
rect 180600 32300 180700 32400
rect 180600 32400 180700 32500
rect 180600 32500 180700 32600
rect 180600 32600 180700 32700
rect 180600 32700 180700 32800
rect 180600 32800 180700 32900
rect 180600 32900 180700 33000
rect 180600 33000 180700 33100
rect 180600 33100 180700 33200
rect 180600 33200 180700 33300
rect 180600 33300 180700 33400
rect 180600 33400 180700 33500
rect 180600 33500 180700 33600
rect 180600 33600 180700 33700
rect 180600 33700 180700 33800
rect 180600 33800 180700 33900
rect 180600 33900 180700 34000
rect 180600 34000 180700 34100
rect 180600 34100 180700 34200
rect 180600 34200 180700 34300
rect 180600 34300 180700 34400
rect 180600 34400 180700 34500
rect 180600 34500 180700 34600
rect 180600 34600 180700 34700
rect 180600 34700 180700 34800
rect 180600 34800 180700 34900
rect 180600 34900 180700 35000
rect 180600 35000 180700 35100
rect 180600 35100 180700 35200
rect 180600 35200 180700 35300
rect 180600 35300 180700 35400
rect 180600 35400 180700 35500
rect 180600 35500 180700 35600
rect 180600 35600 180700 35700
rect 180600 35700 180700 35800
rect 180600 35800 180700 35900
rect 180600 35900 180700 36000
rect 180600 36000 180700 36100
rect 180600 36100 180700 36200
rect 180600 36200 180700 36300
rect 180600 36300 180700 36400
rect 180600 36400 180700 36500
rect 180600 36500 180700 36600
rect 180600 36600 180700 36700
rect 180600 36700 180700 36800
rect 180600 36800 180700 36900
rect 180600 36900 180700 37000
rect 180700 30800 180800 30900
rect 180700 30900 180800 31000
rect 180700 31000 180800 31100
rect 180700 31100 180800 31200
rect 180700 31200 180800 31300
rect 180700 31300 180800 31400
rect 180700 31400 180800 31500
rect 180700 31500 180800 31600
rect 180700 31600 180800 31700
rect 180700 31700 180800 31800
rect 180700 31800 180800 31900
rect 180700 31900 180800 32000
rect 180700 32000 180800 32100
rect 180700 32100 180800 32200
rect 180700 32200 180800 32300
rect 180700 32300 180800 32400
rect 180700 32400 180800 32500
rect 180700 32500 180800 32600
rect 180700 32600 180800 32700
rect 180700 32700 180800 32800
rect 180700 32800 180800 32900
rect 180700 32900 180800 33000
rect 180700 33000 180800 33100
rect 180700 33100 180800 33200
rect 180700 33200 180800 33300
rect 180700 33300 180800 33400
rect 180700 33400 180800 33500
rect 180700 33500 180800 33600
rect 180700 33600 180800 33700
rect 180700 33700 180800 33800
rect 180700 33800 180800 33900
rect 180700 33900 180800 34000
rect 180700 34000 180800 34100
rect 180700 34100 180800 34200
rect 180700 34200 180800 34300
rect 180700 34300 180800 34400
rect 180700 34400 180800 34500
rect 180700 34500 180800 34600
rect 180700 34600 180800 34700
rect 180700 34700 180800 34800
rect 180700 34800 180800 34900
rect 180700 34900 180800 35000
rect 180700 35000 180800 35100
rect 180700 35100 180800 35200
rect 180700 35200 180800 35300
rect 180700 35300 180800 35400
rect 180700 35400 180800 35500
rect 180700 35500 180800 35600
rect 180700 35600 180800 35700
rect 180700 35700 180800 35800
rect 180700 35800 180800 35900
rect 180700 35900 180800 36000
rect 180700 36000 180800 36100
rect 180700 36100 180800 36200
rect 180700 36200 180800 36300
rect 180700 36300 180800 36400
rect 180700 36400 180800 36500
rect 180700 36500 180800 36600
rect 180700 36600 180800 36700
rect 180700 36700 180800 36800
rect 180700 36800 180800 36900
rect 180700 36900 180800 37000
rect 180700 37000 180800 37100
rect 180700 37100 180800 37200
rect 180800 31000 180900 31100
rect 180800 31100 180900 31200
rect 180800 31200 180900 31300
rect 180800 31300 180900 31400
rect 180800 31400 180900 31500
rect 180800 31500 180900 31600
rect 180800 31600 180900 31700
rect 180800 31700 180900 31800
rect 180800 31800 180900 31900
rect 180800 31900 180900 32000
rect 180800 32000 180900 32100
rect 180800 32100 180900 32200
rect 180800 32200 180900 32300
rect 180800 32300 180900 32400
rect 180800 32400 180900 32500
rect 180800 32500 180900 32600
rect 180800 32600 180900 32700
rect 180800 32700 180900 32800
rect 180800 32800 180900 32900
rect 180800 32900 180900 33000
rect 180800 33000 180900 33100
rect 180800 33100 180900 33200
rect 180800 33200 180900 33300
rect 180800 33300 180900 33400
rect 180800 33400 180900 33500
rect 180800 33500 180900 33600
rect 180800 33600 180900 33700
rect 180800 33700 180900 33800
rect 180800 33800 180900 33900
rect 180800 33900 180900 34000
rect 180800 34000 180900 34100
rect 180800 34100 180900 34200
rect 180800 34200 180900 34300
rect 180800 34300 180900 34400
rect 180800 34400 180900 34500
rect 180800 34500 180900 34600
rect 180800 34600 180900 34700
rect 180800 34700 180900 34800
rect 180800 34800 180900 34900
rect 180800 34900 180900 35000
rect 180800 35000 180900 35100
rect 180800 35100 180900 35200
rect 180800 35200 180900 35300
rect 180800 35300 180900 35400
rect 180800 35400 180900 35500
rect 180800 35500 180900 35600
rect 180800 35600 180900 35700
rect 180800 35700 180900 35800
rect 180800 35800 180900 35900
rect 180800 35900 180900 36000
rect 180800 36000 180900 36100
rect 180800 36100 180900 36200
rect 180800 36200 180900 36300
rect 180800 36300 180900 36400
rect 180800 36400 180900 36500
rect 180800 36500 180900 36600
rect 180800 36600 180900 36700
rect 180800 36700 180900 36800
rect 180800 36800 180900 36900
rect 180800 36900 180900 37000
rect 180800 37000 180900 37100
rect 180800 37100 180900 37200
rect 180800 37200 180900 37300
rect 180800 37300 180900 37400
rect 180900 31300 181000 31400
rect 180900 31400 181000 31500
rect 180900 31500 181000 31600
rect 180900 31600 181000 31700
rect 180900 31700 181000 31800
rect 180900 31800 181000 31900
rect 180900 31900 181000 32000
rect 180900 32000 181000 32100
rect 180900 32100 181000 32200
rect 180900 32200 181000 32300
rect 180900 32300 181000 32400
rect 180900 32400 181000 32500
rect 180900 32500 181000 32600
rect 180900 32600 181000 32700
rect 180900 32700 181000 32800
rect 180900 32800 181000 32900
rect 180900 32900 181000 33000
rect 180900 33000 181000 33100
rect 180900 33100 181000 33200
rect 180900 33200 181000 33300
rect 180900 33300 181000 33400
rect 180900 33400 181000 33500
rect 180900 33500 181000 33600
rect 180900 33600 181000 33700
rect 180900 33700 181000 33800
rect 180900 33800 181000 33900
rect 180900 33900 181000 34000
rect 180900 34000 181000 34100
rect 180900 34100 181000 34200
rect 180900 34200 181000 34300
rect 180900 34300 181000 34400
rect 180900 34400 181000 34500
rect 180900 34500 181000 34600
rect 180900 34600 181000 34700
rect 180900 34700 181000 34800
rect 180900 34800 181000 34900
rect 180900 34900 181000 35000
rect 180900 35000 181000 35100
rect 180900 35100 181000 35200
rect 180900 35200 181000 35300
rect 180900 35300 181000 35400
rect 180900 35400 181000 35500
rect 180900 35500 181000 35600
rect 180900 35600 181000 35700
rect 180900 35700 181000 35800
rect 180900 35800 181000 35900
rect 180900 35900 181000 36000
rect 180900 36000 181000 36100
rect 180900 36100 181000 36200
rect 180900 36200 181000 36300
rect 180900 36300 181000 36400
rect 180900 36400 181000 36500
rect 180900 36500 181000 36600
rect 180900 36600 181000 36700
rect 180900 36700 181000 36800
rect 180900 36800 181000 36900
rect 180900 36900 181000 37000
rect 180900 37000 181000 37100
rect 180900 37100 181000 37200
rect 180900 37200 181000 37300
rect 180900 37300 181000 37400
rect 180900 37400 181000 37500
rect 180900 37500 181000 37600
rect 181000 31500 181100 31600
rect 181000 31600 181100 31700
rect 181000 31700 181100 31800
rect 181000 31800 181100 31900
rect 181000 31900 181100 32000
rect 181000 32000 181100 32100
rect 181000 32100 181100 32200
rect 181000 32200 181100 32300
rect 181000 32300 181100 32400
rect 181000 32400 181100 32500
rect 181000 32500 181100 32600
rect 181000 32600 181100 32700
rect 181000 32700 181100 32800
rect 181000 32800 181100 32900
rect 181000 32900 181100 33000
rect 181000 33000 181100 33100
rect 181000 33100 181100 33200
rect 181000 33200 181100 33300
rect 181000 33300 181100 33400
rect 181000 33400 181100 33500
rect 181000 33500 181100 33600
rect 181000 33600 181100 33700
rect 181000 33700 181100 33800
rect 181000 33800 181100 33900
rect 181000 33900 181100 34000
rect 181000 34000 181100 34100
rect 181000 34100 181100 34200
rect 181000 34200 181100 34300
rect 181000 34300 181100 34400
rect 181000 34400 181100 34500
rect 181000 34500 181100 34600
rect 181000 34600 181100 34700
rect 181000 34700 181100 34800
rect 181000 34800 181100 34900
rect 181000 34900 181100 35000
rect 181000 35000 181100 35100
rect 181000 35100 181100 35200
rect 181000 35200 181100 35300
rect 181000 35300 181100 35400
rect 181000 35400 181100 35500
rect 181000 35500 181100 35600
rect 181000 35600 181100 35700
rect 181000 35700 181100 35800
rect 181000 35800 181100 35900
rect 181000 35900 181100 36000
rect 181000 36000 181100 36100
rect 181000 36100 181100 36200
rect 181000 36200 181100 36300
rect 181000 36300 181100 36400
rect 181000 36400 181100 36500
rect 181000 36500 181100 36600
rect 181000 36600 181100 36700
rect 181000 36700 181100 36800
rect 181000 36800 181100 36900
rect 181000 36900 181100 37000
rect 181000 37000 181100 37100
rect 181000 37100 181100 37200
rect 181000 37200 181100 37300
rect 181000 37300 181100 37400
rect 181000 37400 181100 37500
rect 181000 37500 181100 37600
rect 181000 37600 181100 37700
rect 181100 31700 181200 31800
rect 181100 31800 181200 31900
rect 181100 31900 181200 32000
rect 181100 32000 181200 32100
rect 181100 32100 181200 32200
rect 181100 32200 181200 32300
rect 181100 32300 181200 32400
rect 181100 32400 181200 32500
rect 181100 32500 181200 32600
rect 181100 32600 181200 32700
rect 181100 32700 181200 32800
rect 181100 32800 181200 32900
rect 181100 32900 181200 33000
rect 181100 33000 181200 33100
rect 181100 33100 181200 33200
rect 181100 33200 181200 33300
rect 181100 33300 181200 33400
rect 181100 33400 181200 33500
rect 181100 33500 181200 33600
rect 181100 33600 181200 33700
rect 181100 33700 181200 33800
rect 181100 33800 181200 33900
rect 181100 33900 181200 34000
rect 181100 34000 181200 34100
rect 181100 34100 181200 34200
rect 181100 34200 181200 34300
rect 181100 34300 181200 34400
rect 181100 34400 181200 34500
rect 181100 34500 181200 34600
rect 181100 34600 181200 34700
rect 181100 34700 181200 34800
rect 181100 34800 181200 34900
rect 181100 34900 181200 35000
rect 181100 35000 181200 35100
rect 181100 35100 181200 35200
rect 181100 35200 181200 35300
rect 181100 35300 181200 35400
rect 181100 35400 181200 35500
rect 181100 35500 181200 35600
rect 181100 35600 181200 35700
rect 181100 35700 181200 35800
rect 181100 35800 181200 35900
rect 181100 35900 181200 36000
rect 181100 36000 181200 36100
rect 181100 36100 181200 36200
rect 181100 36200 181200 36300
rect 181100 36300 181200 36400
rect 181100 36400 181200 36500
rect 181100 36500 181200 36600
rect 181100 36600 181200 36700
rect 181100 36700 181200 36800
rect 181100 36800 181200 36900
rect 181100 36900 181200 37000
rect 181100 37000 181200 37100
rect 181100 37100 181200 37200
rect 181100 37200 181200 37300
rect 181100 37300 181200 37400
rect 181100 37400 181200 37500
rect 181100 37500 181200 37600
rect 181100 37600 181200 37700
rect 181100 37700 181200 37800
rect 181100 37800 181200 37900
rect 181200 32000 181300 32100
rect 181200 32100 181300 32200
rect 181200 32200 181300 32300
rect 181200 32300 181300 32400
rect 181200 32400 181300 32500
rect 181200 32500 181300 32600
rect 181200 32600 181300 32700
rect 181200 32700 181300 32800
rect 181200 32800 181300 32900
rect 181200 32900 181300 33000
rect 181200 33000 181300 33100
rect 181200 33100 181300 33200
rect 181200 33200 181300 33300
rect 181200 33300 181300 33400
rect 181200 33400 181300 33500
rect 181200 33500 181300 33600
rect 181200 33600 181300 33700
rect 181200 33700 181300 33800
rect 181200 33800 181300 33900
rect 181200 33900 181300 34000
rect 181200 34000 181300 34100
rect 181200 34100 181300 34200
rect 181200 34200 181300 34300
rect 181200 34300 181300 34400
rect 181200 34400 181300 34500
rect 181200 34500 181300 34600
rect 181200 34600 181300 34700
rect 181200 34700 181300 34800
rect 181200 34800 181300 34900
rect 181200 34900 181300 35000
rect 181200 35000 181300 35100
rect 181200 35100 181300 35200
rect 181200 35200 181300 35300
rect 181200 35300 181300 35400
rect 181200 35400 181300 35500
rect 181200 35500 181300 35600
rect 181200 35600 181300 35700
rect 181200 35700 181300 35800
rect 181200 35800 181300 35900
rect 181200 35900 181300 36000
rect 181200 36000 181300 36100
rect 181200 36100 181300 36200
rect 181200 36200 181300 36300
rect 181200 36300 181300 36400
rect 181200 36400 181300 36500
rect 181200 36500 181300 36600
rect 181200 36600 181300 36700
rect 181200 36700 181300 36800
rect 181200 36800 181300 36900
rect 181200 36900 181300 37000
rect 181200 37000 181300 37100
rect 181200 37100 181300 37200
rect 181200 37200 181300 37300
rect 181200 37300 181300 37400
rect 181200 37400 181300 37500
rect 181200 37500 181300 37600
rect 181200 37600 181300 37700
rect 181200 37700 181300 37800
rect 181200 37800 181300 37900
rect 181200 37900 181300 38000
rect 181300 32200 181400 32300
rect 181300 32300 181400 32400
rect 181300 32400 181400 32500
rect 181300 32500 181400 32600
rect 181300 32600 181400 32700
rect 181300 32700 181400 32800
rect 181300 32800 181400 32900
rect 181300 32900 181400 33000
rect 181300 33000 181400 33100
rect 181300 33100 181400 33200
rect 181300 33200 181400 33300
rect 181300 33300 181400 33400
rect 181300 33400 181400 33500
rect 181300 33500 181400 33600
rect 181300 33600 181400 33700
rect 181300 33700 181400 33800
rect 181300 33800 181400 33900
rect 181300 33900 181400 34000
rect 181300 34000 181400 34100
rect 181300 34100 181400 34200
rect 181300 34200 181400 34300
rect 181300 34300 181400 34400
rect 181300 34400 181400 34500
rect 181300 34500 181400 34600
rect 181300 34600 181400 34700
rect 181300 34700 181400 34800
rect 181300 34800 181400 34900
rect 181300 34900 181400 35000
rect 181300 35000 181400 35100
rect 181300 35100 181400 35200
rect 181300 35200 181400 35300
rect 181300 35300 181400 35400
rect 181300 35400 181400 35500
rect 181300 35500 181400 35600
rect 181300 35600 181400 35700
rect 181300 35700 181400 35800
rect 181300 35800 181400 35900
rect 181300 35900 181400 36000
rect 181300 36000 181400 36100
rect 181300 36100 181400 36200
rect 181300 36200 181400 36300
rect 181300 36300 181400 36400
rect 181300 36400 181400 36500
rect 181300 36500 181400 36600
rect 181300 36600 181400 36700
rect 181300 36700 181400 36800
rect 181300 36800 181400 36900
rect 181300 36900 181400 37000
rect 181300 37000 181400 37100
rect 181300 37100 181400 37200
rect 181300 37200 181400 37300
rect 181300 37300 181400 37400
rect 181300 37400 181400 37500
rect 181300 37500 181400 37600
rect 181300 37600 181400 37700
rect 181300 37700 181400 37800
rect 181300 37800 181400 37900
rect 181300 37900 181400 38000
rect 181300 38000 181400 38100
rect 181400 32500 181500 32600
rect 181400 32600 181500 32700
rect 181400 32700 181500 32800
rect 181400 32800 181500 32900
rect 181400 32900 181500 33000
rect 181400 33000 181500 33100
rect 181400 33100 181500 33200
rect 181400 33200 181500 33300
rect 181400 33300 181500 33400
rect 181400 33400 181500 33500
rect 181400 33500 181500 33600
rect 181400 33600 181500 33700
rect 181400 33700 181500 33800
rect 181400 33800 181500 33900
rect 181400 33900 181500 34000
rect 181400 34000 181500 34100
rect 181400 34100 181500 34200
rect 181400 34200 181500 34300
rect 181400 34300 181500 34400
rect 181400 34400 181500 34500
rect 181400 34500 181500 34600
rect 181400 34600 181500 34700
rect 181400 34700 181500 34800
rect 181400 34800 181500 34900
rect 181400 34900 181500 35000
rect 181400 35000 181500 35100
rect 181400 35100 181500 35200
rect 181400 35200 181500 35300
rect 181400 35300 181500 35400
rect 181400 35400 181500 35500
rect 181400 35500 181500 35600
rect 181400 35600 181500 35700
rect 181400 35700 181500 35800
rect 181400 35800 181500 35900
rect 181400 35900 181500 36000
rect 181400 36000 181500 36100
rect 181400 36100 181500 36200
rect 181400 36200 181500 36300
rect 181400 36300 181500 36400
rect 181400 36400 181500 36500
rect 181400 36500 181500 36600
rect 181400 36600 181500 36700
rect 181400 36700 181500 36800
rect 181400 36800 181500 36900
rect 181400 36900 181500 37000
rect 181400 37000 181500 37100
rect 181400 37100 181500 37200
rect 181400 37200 181500 37300
rect 181400 37300 181500 37400
rect 181400 37400 181500 37500
rect 181400 37500 181500 37600
rect 181400 37600 181500 37700
rect 181400 37700 181500 37800
rect 181400 37800 181500 37900
rect 181400 37900 181500 38000
rect 181400 38000 181500 38100
rect 181500 32700 181600 32800
rect 181500 32800 181600 32900
rect 181500 32900 181600 33000
rect 181500 33000 181600 33100
rect 181500 33100 181600 33200
rect 181500 33200 181600 33300
rect 181500 33300 181600 33400
rect 181500 33400 181600 33500
rect 181500 33500 181600 33600
rect 181500 33600 181600 33700
rect 181500 33700 181600 33800
rect 181500 33800 181600 33900
rect 181500 33900 181600 34000
rect 181500 34000 181600 34100
rect 181500 34100 181600 34200
rect 181500 34200 181600 34300
rect 181500 34300 181600 34400
rect 181500 34400 181600 34500
rect 181500 34500 181600 34600
rect 181500 34600 181600 34700
rect 181500 34700 181600 34800
rect 181500 34800 181600 34900
rect 181500 34900 181600 35000
rect 181500 35000 181600 35100
rect 181500 35100 181600 35200
rect 181500 35200 181600 35300
rect 181500 35300 181600 35400
rect 181500 35400 181600 35500
rect 181500 35500 181600 35600
rect 181500 35600 181600 35700
rect 181500 35700 181600 35800
rect 181500 35800 181600 35900
rect 181500 35900 181600 36000
rect 181500 36000 181600 36100
rect 181500 36100 181600 36200
rect 181500 36200 181600 36300
rect 181500 36300 181600 36400
rect 181500 36400 181600 36500
rect 181500 36500 181600 36600
rect 181500 36600 181600 36700
rect 181500 36700 181600 36800
rect 181500 36800 181600 36900
rect 181500 36900 181600 37000
rect 181500 37000 181600 37100
rect 181500 37100 181600 37200
rect 181500 37200 181600 37300
rect 181500 37300 181600 37400
rect 181500 37400 181600 37500
rect 181500 37500 181600 37600
rect 181500 37600 181600 37700
rect 181500 37700 181600 37800
rect 181500 37800 181600 37900
rect 181500 37900 181600 38000
rect 181500 38000 181600 38100
rect 181500 38100 181600 38200
rect 181600 33000 181700 33100
rect 181600 33100 181700 33200
rect 181600 33200 181700 33300
rect 181600 33300 181700 33400
rect 181600 33400 181700 33500
rect 181600 33500 181700 33600
rect 181600 33600 181700 33700
rect 181600 33700 181700 33800
rect 181600 33800 181700 33900
rect 181600 33900 181700 34000
rect 181600 34000 181700 34100
rect 181600 34100 181700 34200
rect 181600 34200 181700 34300
rect 181600 34300 181700 34400
rect 181600 34400 181700 34500
rect 181600 34500 181700 34600
rect 181600 34600 181700 34700
rect 181600 34700 181700 34800
rect 181600 34800 181700 34900
rect 181600 34900 181700 35000
rect 181600 35000 181700 35100
rect 181600 35100 181700 35200
rect 181600 35200 181700 35300
rect 181600 35300 181700 35400
rect 181600 35400 181700 35500
rect 181600 35500 181700 35600
rect 181600 35600 181700 35700
rect 181600 35700 181700 35800
rect 181600 35800 181700 35900
rect 181600 35900 181700 36000
rect 181600 36000 181700 36100
rect 181600 36100 181700 36200
rect 181600 36200 181700 36300
rect 181600 36300 181700 36400
rect 181600 36400 181700 36500
rect 181600 36500 181700 36600
rect 181600 36600 181700 36700
rect 181600 36700 181700 36800
rect 181600 36800 181700 36900
rect 181600 36900 181700 37000
rect 181600 37000 181700 37100
rect 181600 37100 181700 37200
rect 181600 37200 181700 37300
rect 181600 37300 181700 37400
rect 181600 37400 181700 37500
rect 181600 37500 181700 37600
rect 181600 37600 181700 37700
rect 181600 37700 181700 37800
rect 181600 37800 181700 37900
rect 181600 37900 181700 38000
rect 181600 38000 181700 38100
rect 181600 38100 181700 38200
rect 181700 33200 181800 33300
rect 181700 33300 181800 33400
rect 181700 33400 181800 33500
rect 181700 33500 181800 33600
rect 181700 33600 181800 33700
rect 181700 33700 181800 33800
rect 181700 33800 181800 33900
rect 181700 33900 181800 34000
rect 181700 34000 181800 34100
rect 181700 34100 181800 34200
rect 181700 34200 181800 34300
rect 181700 34300 181800 34400
rect 181700 34400 181800 34500
rect 181700 34500 181800 34600
rect 181700 34600 181800 34700
rect 181700 34700 181800 34800
rect 181700 34800 181800 34900
rect 181700 34900 181800 35000
rect 181700 35000 181800 35100
rect 181700 35100 181800 35200
rect 181700 35200 181800 35300
rect 181700 35300 181800 35400
rect 181700 35400 181800 35500
rect 181700 35500 181800 35600
rect 181700 35600 181800 35700
rect 181700 35700 181800 35800
rect 181700 35800 181800 35900
rect 181700 35900 181800 36000
rect 181700 36000 181800 36100
rect 181700 36100 181800 36200
rect 181700 36200 181800 36300
rect 181700 36300 181800 36400
rect 181700 36400 181800 36500
rect 181700 36500 181800 36600
rect 181700 36600 181800 36700
rect 181700 36700 181800 36800
rect 181700 36800 181800 36900
rect 181700 36900 181800 37000
rect 181700 37000 181800 37100
rect 181700 37100 181800 37200
rect 181700 37200 181800 37300
rect 181700 37300 181800 37400
rect 181700 37400 181800 37500
rect 181700 37500 181800 37600
rect 181700 37600 181800 37700
rect 181700 37700 181800 37800
rect 181700 37800 181800 37900
rect 181700 37900 181800 38000
rect 181700 38000 181800 38100
rect 181700 38100 181800 38200
rect 181700 38200 181800 38300
rect 181800 33500 181900 33600
rect 181800 33600 181900 33700
rect 181800 33700 181900 33800
rect 181800 33800 181900 33900
rect 181800 33900 181900 34000
rect 181800 34000 181900 34100
rect 181800 34100 181900 34200
rect 181800 34200 181900 34300
rect 181800 34300 181900 34400
rect 181800 34400 181900 34500
rect 181800 34500 181900 34600
rect 181800 34600 181900 34700
rect 181800 34700 181900 34800
rect 181800 34800 181900 34900
rect 181800 34900 181900 35000
rect 181800 35000 181900 35100
rect 181800 35100 181900 35200
rect 181800 35200 181900 35300
rect 181800 35300 181900 35400
rect 181800 35400 181900 35500
rect 181800 35500 181900 35600
rect 181800 35600 181900 35700
rect 181800 35700 181900 35800
rect 181800 35800 181900 35900
rect 181800 35900 181900 36000
rect 181800 36000 181900 36100
rect 181800 36100 181900 36200
rect 181800 36200 181900 36300
rect 181800 36300 181900 36400
rect 181800 36400 181900 36500
rect 181800 36500 181900 36600
rect 181800 36600 181900 36700
rect 181800 36700 181900 36800
rect 181800 36800 181900 36900
rect 181800 36900 181900 37000
rect 181800 37000 181900 37100
rect 181800 37100 181900 37200
rect 181800 37200 181900 37300
rect 181800 37300 181900 37400
rect 181800 37400 181900 37500
rect 181800 37500 181900 37600
rect 181800 37600 181900 37700
rect 181800 37700 181900 37800
rect 181800 37800 181900 37900
rect 181800 37900 181900 38000
rect 181800 38000 181900 38100
rect 181800 38100 181900 38200
rect 181800 38200 181900 38300
rect 181900 33800 182000 33900
rect 181900 33900 182000 34000
rect 181900 34000 182000 34100
rect 181900 34100 182000 34200
rect 181900 34200 182000 34300
rect 181900 34300 182000 34400
rect 181900 34400 182000 34500
rect 181900 34500 182000 34600
rect 181900 34600 182000 34700
rect 181900 34700 182000 34800
rect 181900 34800 182000 34900
rect 181900 34900 182000 35000
rect 181900 35000 182000 35100
rect 181900 35100 182000 35200
rect 181900 35200 182000 35300
rect 181900 35300 182000 35400
rect 181900 35400 182000 35500
rect 181900 35500 182000 35600
rect 181900 35600 182000 35700
rect 181900 35700 182000 35800
rect 181900 35800 182000 35900
rect 181900 35900 182000 36000
rect 181900 36000 182000 36100
rect 181900 36100 182000 36200
rect 181900 36200 182000 36300
rect 181900 36300 182000 36400
rect 181900 36400 182000 36500
rect 181900 36500 182000 36600
rect 181900 36600 182000 36700
rect 181900 36700 182000 36800
rect 181900 36800 182000 36900
rect 181900 36900 182000 37000
rect 181900 37000 182000 37100
rect 181900 37100 182000 37200
rect 181900 37200 182000 37300
rect 181900 37300 182000 37400
rect 181900 37400 182000 37500
rect 181900 37500 182000 37600
rect 181900 37600 182000 37700
rect 181900 37700 182000 37800
rect 181900 37800 182000 37900
rect 181900 37900 182000 38000
rect 181900 38000 182000 38100
rect 181900 38100 182000 38200
rect 181900 38200 182000 38300
rect 182000 34200 182100 34300
rect 182000 34300 182100 34400
rect 182000 34400 182100 34500
rect 182000 34500 182100 34600
rect 182000 34600 182100 34700
rect 182000 34700 182100 34800
rect 182000 34800 182100 34900
rect 182000 34900 182100 35000
rect 182000 35000 182100 35100
rect 182000 35100 182100 35200
rect 182000 35200 182100 35300
rect 182000 35300 182100 35400
rect 182000 35400 182100 35500
rect 182000 35500 182100 35600
rect 182000 35600 182100 35700
rect 182000 35700 182100 35800
rect 182000 35800 182100 35900
rect 182000 35900 182100 36000
rect 182000 36000 182100 36100
rect 182000 36100 182100 36200
rect 182000 36200 182100 36300
rect 182000 36300 182100 36400
rect 182000 36400 182100 36500
rect 182000 36500 182100 36600
rect 182000 36600 182100 36700
rect 182000 36700 182100 36800
rect 182000 36800 182100 36900
rect 182000 36900 182100 37000
rect 182000 37000 182100 37100
rect 182000 37100 182100 37200
rect 182000 37200 182100 37300
rect 182000 37300 182100 37400
rect 182000 37400 182100 37500
rect 182000 37500 182100 37600
rect 182000 37600 182100 37700
rect 182000 37700 182100 37800
rect 182000 37800 182100 37900
rect 182000 37900 182100 38000
rect 182000 38000 182100 38100
rect 182000 38100 182100 38200
rect 182000 38200 182100 38300
rect 182100 34500 182200 34600
rect 182100 34600 182200 34700
rect 182100 34700 182200 34800
rect 182100 34800 182200 34900
rect 182100 34900 182200 35000
rect 182100 35000 182200 35100
rect 182100 35100 182200 35200
rect 182100 35200 182200 35300
rect 182100 35300 182200 35400
rect 182100 35400 182200 35500
rect 182100 35500 182200 35600
rect 182100 35600 182200 35700
rect 182100 35700 182200 35800
rect 182100 35800 182200 35900
rect 182100 35900 182200 36000
rect 182100 36000 182200 36100
rect 182100 36100 182200 36200
rect 182100 36200 182200 36300
rect 182100 36300 182200 36400
rect 182100 36400 182200 36500
rect 182100 36500 182200 36600
rect 182100 36600 182200 36700
rect 182100 36700 182200 36800
rect 182100 36800 182200 36900
rect 182100 36900 182200 37000
rect 182100 37000 182200 37100
rect 182100 37100 182200 37200
rect 182100 37200 182200 37300
rect 182100 37300 182200 37400
rect 182100 37400 182200 37500
rect 182100 37500 182200 37600
rect 182100 37600 182200 37700
rect 182100 37700 182200 37800
rect 182100 37800 182200 37900
rect 182100 37900 182200 38000
rect 182100 38000 182200 38100
rect 182100 38100 182200 38200
rect 182100 38200 182200 38300
rect 182200 34800 182300 34900
rect 182200 34900 182300 35000
rect 182200 35000 182300 35100
rect 182200 35100 182300 35200
rect 182200 35200 182300 35300
rect 182200 35300 182300 35400
rect 182200 35400 182300 35500
rect 182200 35500 182300 35600
rect 182200 35600 182300 35700
rect 182200 35700 182300 35800
rect 182200 35800 182300 35900
rect 182200 35900 182300 36000
rect 182200 36000 182300 36100
rect 182200 36100 182300 36200
rect 182200 36200 182300 36300
rect 182200 36300 182300 36400
rect 182200 36400 182300 36500
rect 182200 36500 182300 36600
rect 182200 36600 182300 36700
rect 182200 36700 182300 36800
rect 182200 36800 182300 36900
rect 182200 36900 182300 37000
rect 182200 37000 182300 37100
rect 182200 37100 182300 37200
rect 182200 37200 182300 37300
rect 182200 37300 182300 37400
rect 182200 37400 182300 37500
rect 182200 37500 182300 37600
rect 182200 37600 182300 37700
rect 182200 37700 182300 37800
rect 182200 37800 182300 37900
rect 182200 37900 182300 38000
rect 182200 38000 182300 38100
rect 182200 38100 182300 38200
rect 182200 38200 182300 38300
rect 182300 35100 182400 35200
rect 182300 35200 182400 35300
rect 182300 35300 182400 35400
rect 182300 35400 182400 35500
rect 182300 35500 182400 35600
rect 182300 35600 182400 35700
rect 182300 35700 182400 35800
rect 182300 35800 182400 35900
rect 182300 35900 182400 36000
rect 182300 36000 182400 36100
rect 182300 36100 182400 36200
rect 182300 36200 182400 36300
rect 182300 36300 182400 36400
rect 182300 36400 182400 36500
rect 182300 36500 182400 36600
rect 182300 36600 182400 36700
rect 182300 36700 182400 36800
rect 182300 36800 182400 36900
rect 182300 36900 182400 37000
rect 182300 37000 182400 37100
rect 182300 37100 182400 37200
rect 182300 37200 182400 37300
rect 182300 37300 182400 37400
rect 182300 37400 182400 37500
rect 182300 37500 182400 37600
rect 182300 37600 182400 37700
rect 182300 37700 182400 37800
rect 182300 37800 182400 37900
rect 182300 37900 182400 38000
rect 182300 38000 182400 38100
rect 182300 38100 182400 38200
rect 182300 38200 182400 38300
rect 182400 35400 182500 35500
rect 182400 35500 182500 35600
rect 182400 35600 182500 35700
rect 182400 35700 182500 35800
rect 182400 35800 182500 35900
rect 182400 35900 182500 36000
rect 182400 36000 182500 36100
rect 182400 36100 182500 36200
rect 182400 36200 182500 36300
rect 182400 36300 182500 36400
rect 182400 36400 182500 36500
rect 182400 36500 182500 36600
rect 182400 36600 182500 36700
rect 182400 36700 182500 36800
rect 182400 36800 182500 36900
rect 182400 36900 182500 37000
rect 182400 37000 182500 37100
rect 182400 37100 182500 37200
rect 182400 37200 182500 37300
rect 182400 37300 182500 37400
rect 182400 37400 182500 37500
rect 182400 37500 182500 37600
rect 182400 37600 182500 37700
rect 182400 37700 182500 37800
rect 182400 37800 182500 37900
rect 182400 37900 182500 38000
rect 182400 38000 182500 38100
rect 182400 38100 182500 38200
rect 182500 35700 182600 35800
rect 182500 35800 182600 35900
rect 182500 35900 182600 36000
rect 182500 36000 182600 36100
rect 182500 36100 182600 36200
rect 182500 36200 182600 36300
rect 182500 36300 182600 36400
rect 182500 36400 182600 36500
rect 182500 36500 182600 36600
rect 182500 36600 182600 36700
rect 182500 36700 182600 36800
rect 182500 36800 182600 36900
rect 182500 36900 182600 37000
rect 182500 37000 182600 37100
rect 182500 37100 182600 37200
rect 182500 37200 182600 37300
rect 182500 37300 182600 37400
rect 182500 37400 182600 37500
rect 182500 37500 182600 37600
rect 182500 37600 182600 37700
rect 182500 37700 182600 37800
rect 182500 37800 182600 37900
rect 182500 37900 182600 38000
rect 182500 38000 182600 38100
rect 182500 38100 182600 38200
rect 182600 35900 182700 36000
rect 182600 36000 182700 36100
rect 182600 36100 182700 36200
rect 182600 36200 182700 36300
rect 182600 36300 182700 36400
rect 182600 36400 182700 36500
rect 182600 36500 182700 36600
rect 182600 36600 182700 36700
rect 182600 36700 182700 36800
rect 182600 36800 182700 36900
rect 182600 36900 182700 37000
rect 182600 37000 182700 37100
rect 182600 37100 182700 37200
rect 182600 37200 182700 37300
rect 182600 37300 182700 37400
rect 182600 37400 182700 37500
rect 182600 37500 182700 37600
rect 182600 37600 182700 37700
rect 182600 37700 182700 37800
rect 182600 37800 182700 37900
rect 182600 37900 182700 38000
rect 182600 38000 182700 38100
rect 182600 38100 182700 38200
rect 182700 36200 182800 36300
rect 182700 36300 182800 36400
rect 182700 36400 182800 36500
rect 182700 36500 182800 36600
rect 182700 36600 182800 36700
rect 182700 36700 182800 36800
rect 182700 36800 182800 36900
rect 182700 36900 182800 37000
rect 182700 37000 182800 37100
rect 182700 37100 182800 37200
rect 182700 37200 182800 37300
rect 182700 37300 182800 37400
rect 182700 37400 182800 37500
rect 182700 37500 182800 37600
rect 182700 37600 182800 37700
rect 182700 37700 182800 37800
rect 182700 37800 182800 37900
rect 182700 37900 182800 38000
rect 182700 38000 182800 38100
rect 182700 38100 182800 38200
rect 182800 36400 182900 36500
rect 182800 36500 182900 36600
rect 182800 36600 182900 36700
rect 182800 36700 182900 36800
rect 182800 36800 182900 36900
rect 182800 36900 182900 37000
rect 182800 37000 182900 37100
rect 182800 37100 182900 37200
rect 182800 37200 182900 37300
rect 182800 37300 182900 37400
rect 182800 37400 182900 37500
rect 182800 37500 182900 37600
rect 182800 37600 182900 37700
rect 182800 37700 182900 37800
rect 182800 37800 182900 37900
rect 182800 37900 182900 38000
rect 182800 38000 182900 38100
rect 182900 36500 183000 36600
rect 182900 36600 183000 36700
rect 182900 36700 183000 36800
rect 182900 36800 183000 36900
rect 182900 36900 183000 37000
rect 182900 37000 183000 37100
rect 182900 37100 183000 37200
rect 182900 37200 183000 37300
rect 182900 37300 183000 37400
rect 182900 37400 183000 37500
rect 182900 37500 183000 37600
rect 182900 37600 183000 37700
rect 182900 37700 183000 37800
rect 182900 37800 183000 37900
rect 182900 37900 183000 38000
rect 182900 38000 183000 38100
rect 183000 36600 183100 36700
rect 183000 36700 183100 36800
rect 183000 36800 183100 36900
rect 183000 36900 183100 37000
rect 183000 37000 183100 37100
rect 183000 37100 183100 37200
rect 183000 37200 183100 37300
rect 183000 37300 183100 37400
rect 183000 37400 183100 37500
rect 183000 37500 183100 37600
rect 183000 37600 183100 37700
rect 183000 37700 183100 37800
rect 183000 37800 183100 37900
rect 183000 37900 183100 38000
rect 183100 36700 183200 36800
rect 183100 36800 183200 36900
rect 183100 36900 183200 37000
rect 183100 37000 183200 37100
rect 183100 37100 183200 37200
rect 183100 37200 183200 37300
rect 183100 37300 183200 37400
rect 183100 37400 183200 37500
rect 183100 37500 183200 37600
rect 183100 37600 183200 37700
rect 183100 37700 183200 37800
rect 183100 37800 183200 37900
rect 183100 37900 183200 38000
rect 183200 36700 183300 36800
rect 183200 36800 183300 36900
rect 183200 36900 183300 37000
rect 183200 37000 183300 37100
rect 183200 37100 183300 37200
rect 183200 37200 183300 37300
rect 183200 37300 183300 37400
rect 183200 37400 183300 37500
rect 183200 37500 183300 37600
rect 183200 37600 183300 37700
rect 183200 37700 183300 37800
rect 183200 37800 183300 37900
rect 183300 36800 183400 36900
rect 183300 36900 183400 37000
rect 183300 37000 183400 37100
rect 183300 37100 183400 37200
rect 183300 37200 183400 37300
rect 183300 37300 183400 37400
rect 183300 37400 183400 37500
rect 183300 37500 183400 37600
rect 183300 37600 183400 37700
rect 183300 37700 183400 37800
rect 183300 37800 183400 37900
rect 183400 36800 183500 36900
rect 183400 36900 183500 37000
rect 183400 37000 183500 37100
rect 183400 37100 183500 37200
rect 183400 37200 183500 37300
rect 183400 37300 183500 37400
rect 183400 37400 183500 37500
rect 183400 37500 183500 37600
rect 183400 37600 183500 37700
rect 183400 37700 183500 37800
rect 183500 36900 183600 37000
rect 183500 37000 183600 37100
rect 183500 37100 183600 37200
rect 183500 37200 183600 37300
rect 183500 37300 183600 37400
rect 183500 37400 183600 37500
rect 183500 37500 183600 37600
rect 183500 37600 183600 37700
rect 183600 36900 183700 37000
rect 183600 37000 183700 37100
rect 183600 37100 183700 37200
rect 183600 37200 183700 37300
rect 183600 37300 183700 37400
rect 183600 37400 183700 37500
rect 183600 37500 183700 37600
rect 183700 37000 183800 37100
rect 183700 37100 183800 37200
rect 183700 37200 183800 37300
rect 183700 37300 183800 37400
rect 183700 37400 183800 37500
rect 183800 37100 183900 37200
rect 183800 37200 183900 37300
rect 185300 21900 185400 22000
rect 185300 22000 185400 22100
rect 185300 22100 185400 22200
rect 185300 22200 185400 22300
rect 185300 22300 185400 22400
rect 185300 22400 185400 22500
rect 185300 22500 185400 22600
rect 185300 22600 185400 22700
rect 185300 22700 185400 22800
rect 185300 22800 185400 22900
rect 185300 22900 185400 23000
rect 185300 23000 185400 23100
rect 185300 23100 185400 23200
rect 185400 21700 185500 21800
rect 185400 21800 185500 21900
rect 185400 21900 185500 22000
rect 185400 22000 185500 22100
rect 185400 22100 185500 22200
rect 185400 22200 185500 22300
rect 185400 22300 185500 22400
rect 185400 22400 185500 22500
rect 185400 22500 185500 22600
rect 185400 22600 185500 22700
rect 185400 22700 185500 22800
rect 185400 22800 185500 22900
rect 185400 22900 185500 23000
rect 185400 23000 185500 23100
rect 185400 23100 185500 23200
rect 185400 23200 185500 23300
rect 185400 23300 185500 23400
rect 185400 23400 185500 23500
rect 185400 23500 185500 23600
rect 185400 23600 185500 23700
rect 185400 23700 185500 23800
rect 185400 23800 185500 23900
rect 185400 23900 185500 24000
rect 185400 24000 185500 24100
rect 185400 24100 185500 24200
rect 185400 24200 185500 24300
rect 185400 24300 185500 24400
rect 185400 24400 185500 24500
rect 185400 24500 185500 24600
rect 185400 24700 185500 24800
rect 185400 24900 185500 25000
rect 185400 25100 185500 25200
rect 185400 25300 185500 25400
rect 185400 25500 185500 25600
rect 185400 25800 185500 25900
rect 185500 21600 185600 21700
rect 185500 21700 185600 21800
rect 185500 21800 185600 21900
rect 185500 21900 185600 22000
rect 185500 22000 185600 22100
rect 185500 22100 185600 22200
rect 185500 22200 185600 22300
rect 185500 22300 185600 22400
rect 185500 22400 185600 22500
rect 185500 22500 185600 22600
rect 185500 22600 185600 22700
rect 185500 22700 185600 22800
rect 185500 22800 185600 22900
rect 185500 22900 185600 23000
rect 185500 23000 185600 23100
rect 185500 23100 185600 23200
rect 185500 23200 185600 23300
rect 185500 23300 185600 23400
rect 185500 23400 185600 23500
rect 185500 23500 185600 23600
rect 185500 23600 185600 23700
rect 185500 23700 185600 23800
rect 185500 23800 185600 23900
rect 185500 23900 185600 24000
rect 185500 24000 185600 24100
rect 185500 24100 185600 24200
rect 185500 24200 185600 24300
rect 185500 24300 185600 24400
rect 185500 24400 185600 24500
rect 185500 24500 185600 24600
rect 185500 24600 185600 24700
rect 185500 24700 185600 24800
rect 185500 24800 185600 24900
rect 185500 24900 185600 25000
rect 185500 25000 185600 25100
rect 185500 25100 185600 25200
rect 185500 25200 185600 25300
rect 185500 25300 185600 25400
rect 185500 25400 185600 25500
rect 185500 25500 185600 25600
rect 185500 25600 185600 25700
rect 185500 25700 185600 25800
rect 185500 25800 185600 25900
rect 185500 25900 185600 26000
rect 185500 26000 185600 26100
rect 185500 26100 185600 26200
rect 185500 26200 185600 26300
rect 185500 26300 185600 26400
rect 185500 26400 185600 26500
rect 185500 26500 185600 26600
rect 185500 26600 185600 26700
rect 185500 26700 185600 26800
rect 185500 26800 185600 26900
rect 185500 26900 185600 27000
rect 185500 27000 185600 27100
rect 185500 27100 185600 27200
rect 185500 27200 185600 27300
rect 185500 27300 185600 27400
rect 185500 27400 185600 27500
rect 185500 27500 185600 27600
rect 185500 27600 185600 27700
rect 185500 27700 185600 27800
rect 185500 27800 185600 27900
rect 185500 27900 185600 28000
rect 185500 28000 185600 28100
rect 185500 28100 185600 28200
rect 185500 28200 185600 28300
rect 185500 28300 185600 28400
rect 185500 28400 185600 28500
rect 185500 28500 185600 28600
rect 185500 28700 185600 28800
rect 185500 36000 185600 36100
rect 185500 36100 185600 36200
rect 185500 36200 185600 36300
rect 185500 36300 185600 36400
rect 185500 36400 185600 36500
rect 185500 36500 185600 36600
rect 185500 36600 185600 36700
rect 185500 36700 185600 36800
rect 185500 36800 185600 36900
rect 185500 36900 185600 37000
rect 185600 21500 185700 21600
rect 185600 21600 185700 21700
rect 185600 21700 185700 21800
rect 185600 21800 185700 21900
rect 185600 21900 185700 22000
rect 185600 22000 185700 22100
rect 185600 22100 185700 22200
rect 185600 22200 185700 22300
rect 185600 22300 185700 22400
rect 185600 22400 185700 22500
rect 185600 22500 185700 22600
rect 185600 22600 185700 22700
rect 185600 22700 185700 22800
rect 185600 22800 185700 22900
rect 185600 22900 185700 23000
rect 185600 23000 185700 23100
rect 185600 23100 185700 23200
rect 185600 23200 185700 23300
rect 185600 23300 185700 23400
rect 185600 23400 185700 23500
rect 185600 23500 185700 23600
rect 185600 23600 185700 23700
rect 185600 23700 185700 23800
rect 185600 23800 185700 23900
rect 185600 23900 185700 24000
rect 185600 24000 185700 24100
rect 185600 24100 185700 24200
rect 185600 24200 185700 24300
rect 185600 24300 185700 24400
rect 185600 24400 185700 24500
rect 185600 24500 185700 24600
rect 185600 24600 185700 24700
rect 185600 24700 185700 24800
rect 185600 24800 185700 24900
rect 185600 24900 185700 25000
rect 185600 25000 185700 25100
rect 185600 25100 185700 25200
rect 185600 25200 185700 25300
rect 185600 25300 185700 25400
rect 185600 25400 185700 25500
rect 185600 25500 185700 25600
rect 185600 25600 185700 25700
rect 185600 25700 185700 25800
rect 185600 25800 185700 25900
rect 185600 25900 185700 26000
rect 185600 26000 185700 26100
rect 185600 26100 185700 26200
rect 185600 26200 185700 26300
rect 185600 26300 185700 26400
rect 185600 26400 185700 26500
rect 185600 26500 185700 26600
rect 185600 26600 185700 26700
rect 185600 26700 185700 26800
rect 185600 26800 185700 26900
rect 185600 26900 185700 27000
rect 185600 27000 185700 27100
rect 185600 27100 185700 27200
rect 185600 27200 185700 27300
rect 185600 27300 185700 27400
rect 185600 27400 185700 27500
rect 185600 27500 185700 27600
rect 185600 27600 185700 27700
rect 185600 27700 185700 27800
rect 185600 27800 185700 27900
rect 185600 27900 185700 28000
rect 185600 28000 185700 28100
rect 185600 28100 185700 28200
rect 185600 28200 185700 28300
rect 185600 28300 185700 28400
rect 185600 28400 185700 28500
rect 185600 28500 185700 28600
rect 185600 28600 185700 28700
rect 185600 28700 185700 28800
rect 185600 28800 185700 28900
rect 185600 28900 185700 29000
rect 185600 29000 185700 29100
rect 185600 29100 185700 29200
rect 185600 29200 185700 29300
rect 185600 29300 185700 29400
rect 185600 29400 185700 29500
rect 185600 29500 185700 29600
rect 185600 29600 185700 29700
rect 185600 29700 185700 29800
rect 185600 29800 185700 29900
rect 185600 29900 185700 30000
rect 185600 30000 185700 30100
rect 185600 30100 185700 30200
rect 185600 30300 185700 30400
rect 185600 35800 185700 35900
rect 185600 35900 185700 36000
rect 185600 36000 185700 36100
rect 185600 36100 185700 36200
rect 185600 36200 185700 36300
rect 185600 36300 185700 36400
rect 185600 36400 185700 36500
rect 185600 36500 185700 36600
rect 185600 36600 185700 36700
rect 185600 36700 185700 36800
rect 185600 36800 185700 36900
rect 185600 36900 185700 37000
rect 185600 37000 185700 37100
rect 185600 37100 185700 37200
rect 185600 37200 185700 37300
rect 185600 37300 185700 37400
rect 185700 21400 185800 21500
rect 185700 21500 185800 21600
rect 185700 21600 185800 21700
rect 185700 21700 185800 21800
rect 185700 21800 185800 21900
rect 185700 21900 185800 22000
rect 185700 22000 185800 22100
rect 185700 22100 185800 22200
rect 185700 22200 185800 22300
rect 185700 22300 185800 22400
rect 185700 22400 185800 22500
rect 185700 22500 185800 22600
rect 185700 22600 185800 22700
rect 185700 22700 185800 22800
rect 185700 22800 185800 22900
rect 185700 22900 185800 23000
rect 185700 23000 185800 23100
rect 185700 23100 185800 23200
rect 185700 23200 185800 23300
rect 185700 23300 185800 23400
rect 185700 23400 185800 23500
rect 185700 23500 185800 23600
rect 185700 23600 185800 23700
rect 185700 23700 185800 23800
rect 185700 23800 185800 23900
rect 185700 23900 185800 24000
rect 185700 24000 185800 24100
rect 185700 24100 185800 24200
rect 185700 24200 185800 24300
rect 185700 24300 185800 24400
rect 185700 24400 185800 24500
rect 185700 24500 185800 24600
rect 185700 24600 185800 24700
rect 185700 24700 185800 24800
rect 185700 24800 185800 24900
rect 185700 24900 185800 25000
rect 185700 25000 185800 25100
rect 185700 25100 185800 25200
rect 185700 25200 185800 25300
rect 185700 25300 185800 25400
rect 185700 25400 185800 25500
rect 185700 25500 185800 25600
rect 185700 25600 185800 25700
rect 185700 25700 185800 25800
rect 185700 25800 185800 25900
rect 185700 25900 185800 26000
rect 185700 26000 185800 26100
rect 185700 26100 185800 26200
rect 185700 26200 185800 26300
rect 185700 26300 185800 26400
rect 185700 26400 185800 26500
rect 185700 26500 185800 26600
rect 185700 26600 185800 26700
rect 185700 26700 185800 26800
rect 185700 26800 185800 26900
rect 185700 26900 185800 27000
rect 185700 27000 185800 27100
rect 185700 27100 185800 27200
rect 185700 27200 185800 27300
rect 185700 27300 185800 27400
rect 185700 27400 185800 27500
rect 185700 27500 185800 27600
rect 185700 27600 185800 27700
rect 185700 27700 185800 27800
rect 185700 27800 185800 27900
rect 185700 27900 185800 28000
rect 185700 28000 185800 28100
rect 185700 28100 185800 28200
rect 185700 28200 185800 28300
rect 185700 28300 185800 28400
rect 185700 28400 185800 28500
rect 185700 28500 185800 28600
rect 185700 28600 185800 28700
rect 185700 28700 185800 28800
rect 185700 28800 185800 28900
rect 185700 28900 185800 29000
rect 185700 29000 185800 29100
rect 185700 29100 185800 29200
rect 185700 29200 185800 29300
rect 185700 29300 185800 29400
rect 185700 29400 185800 29500
rect 185700 29500 185800 29600
rect 185700 29600 185800 29700
rect 185700 29700 185800 29800
rect 185700 29800 185800 29900
rect 185700 29900 185800 30000
rect 185700 30000 185800 30100
rect 185700 30100 185800 30200
rect 185700 30200 185800 30300
rect 185700 30300 185800 30400
rect 185700 30400 185800 30500
rect 185700 30500 185800 30600
rect 185700 30600 185800 30700
rect 185700 30700 185800 30800
rect 185700 30800 185800 30900
rect 185700 30900 185800 31000
rect 185700 31000 185800 31100
rect 185700 31100 185800 31200
rect 185700 31200 185800 31300
rect 185700 31300 185800 31400
rect 185700 31400 185800 31500
rect 185700 35600 185800 35700
rect 185700 35700 185800 35800
rect 185700 35800 185800 35900
rect 185700 35900 185800 36000
rect 185700 36000 185800 36100
rect 185700 36100 185800 36200
rect 185700 36200 185800 36300
rect 185700 36300 185800 36400
rect 185700 36400 185800 36500
rect 185700 36500 185800 36600
rect 185700 36600 185800 36700
rect 185700 36700 185800 36800
rect 185700 36800 185800 36900
rect 185700 36900 185800 37000
rect 185700 37000 185800 37100
rect 185700 37100 185800 37200
rect 185700 37200 185800 37300
rect 185700 37300 185800 37400
rect 185700 37400 185800 37500
rect 185700 37500 185800 37600
rect 185800 21400 185900 21500
rect 185800 21500 185900 21600
rect 185800 21600 185900 21700
rect 185800 21700 185900 21800
rect 185800 21800 185900 21900
rect 185800 21900 185900 22000
rect 185800 22000 185900 22100
rect 185800 22100 185900 22200
rect 185800 22200 185900 22300
rect 185800 22300 185900 22400
rect 185800 22400 185900 22500
rect 185800 22500 185900 22600
rect 185800 22600 185900 22700
rect 185800 22700 185900 22800
rect 185800 22800 185900 22900
rect 185800 22900 185900 23000
rect 185800 23000 185900 23100
rect 185800 23100 185900 23200
rect 185800 23200 185900 23300
rect 185800 23300 185900 23400
rect 185800 23400 185900 23500
rect 185800 23500 185900 23600
rect 185800 23600 185900 23700
rect 185800 23700 185900 23800
rect 185800 23800 185900 23900
rect 185800 23900 185900 24000
rect 185800 24000 185900 24100
rect 185800 24100 185900 24200
rect 185800 24200 185900 24300
rect 185800 24300 185900 24400
rect 185800 24400 185900 24500
rect 185800 24500 185900 24600
rect 185800 24600 185900 24700
rect 185800 24700 185900 24800
rect 185800 24800 185900 24900
rect 185800 24900 185900 25000
rect 185800 25000 185900 25100
rect 185800 25100 185900 25200
rect 185800 25200 185900 25300
rect 185800 25300 185900 25400
rect 185800 25400 185900 25500
rect 185800 25500 185900 25600
rect 185800 25600 185900 25700
rect 185800 25700 185900 25800
rect 185800 25800 185900 25900
rect 185800 25900 185900 26000
rect 185800 26000 185900 26100
rect 185800 26100 185900 26200
rect 185800 26200 185900 26300
rect 185800 26300 185900 26400
rect 185800 26400 185900 26500
rect 185800 26500 185900 26600
rect 185800 26600 185900 26700
rect 185800 26700 185900 26800
rect 185800 26800 185900 26900
rect 185800 26900 185900 27000
rect 185800 27000 185900 27100
rect 185800 27100 185900 27200
rect 185800 27200 185900 27300
rect 185800 27300 185900 27400
rect 185800 27400 185900 27500
rect 185800 27500 185900 27600
rect 185800 27600 185900 27700
rect 185800 27700 185900 27800
rect 185800 27800 185900 27900
rect 185800 27900 185900 28000
rect 185800 28000 185900 28100
rect 185800 28100 185900 28200
rect 185800 28200 185900 28300
rect 185800 28300 185900 28400
rect 185800 28400 185900 28500
rect 185800 28500 185900 28600
rect 185800 28600 185900 28700
rect 185800 28700 185900 28800
rect 185800 28800 185900 28900
rect 185800 28900 185900 29000
rect 185800 29000 185900 29100
rect 185800 29100 185900 29200
rect 185800 29200 185900 29300
rect 185800 29300 185900 29400
rect 185800 29400 185900 29500
rect 185800 29500 185900 29600
rect 185800 29600 185900 29700
rect 185800 29700 185900 29800
rect 185800 29800 185900 29900
rect 185800 29900 185900 30000
rect 185800 30000 185900 30100
rect 185800 30100 185900 30200
rect 185800 30200 185900 30300
rect 185800 30300 185900 30400
rect 185800 30400 185900 30500
rect 185800 30500 185900 30600
rect 185800 30600 185900 30700
rect 185800 30700 185900 30800
rect 185800 30800 185900 30900
rect 185800 30900 185900 31000
rect 185800 31000 185900 31100
rect 185800 31100 185900 31200
rect 185800 31200 185900 31300
rect 185800 31300 185900 31400
rect 185800 31400 185900 31500
rect 185800 31500 185900 31600
rect 185800 31600 185900 31700
rect 185800 31700 185900 31800
rect 185800 35400 185900 35500
rect 185800 35500 185900 35600
rect 185800 35600 185900 35700
rect 185800 35700 185900 35800
rect 185800 35800 185900 35900
rect 185800 35900 185900 36000
rect 185800 36000 185900 36100
rect 185800 36100 185900 36200
rect 185800 36200 185900 36300
rect 185800 36300 185900 36400
rect 185800 36400 185900 36500
rect 185800 36500 185900 36600
rect 185800 36600 185900 36700
rect 185800 36700 185900 36800
rect 185800 36800 185900 36900
rect 185800 36900 185900 37000
rect 185800 37000 185900 37100
rect 185800 37100 185900 37200
rect 185800 37200 185900 37300
rect 185800 37300 185900 37400
rect 185800 37400 185900 37500
rect 185800 37500 185900 37600
rect 185800 37600 185900 37700
rect 185800 37700 185900 37800
rect 185900 21300 186000 21400
rect 185900 21400 186000 21500
rect 185900 21500 186000 21600
rect 185900 21600 186000 21700
rect 185900 21700 186000 21800
rect 185900 21800 186000 21900
rect 185900 21900 186000 22000
rect 185900 22000 186000 22100
rect 185900 22100 186000 22200
rect 185900 22200 186000 22300
rect 185900 22300 186000 22400
rect 185900 22400 186000 22500
rect 185900 22500 186000 22600
rect 185900 22600 186000 22700
rect 185900 22700 186000 22800
rect 185900 22800 186000 22900
rect 185900 22900 186000 23000
rect 185900 23000 186000 23100
rect 185900 23100 186000 23200
rect 185900 23200 186000 23300
rect 185900 23300 186000 23400
rect 185900 23400 186000 23500
rect 185900 23500 186000 23600
rect 185900 23600 186000 23700
rect 185900 23700 186000 23800
rect 185900 23800 186000 23900
rect 185900 23900 186000 24000
rect 185900 24000 186000 24100
rect 185900 24100 186000 24200
rect 185900 24200 186000 24300
rect 185900 24300 186000 24400
rect 185900 24400 186000 24500
rect 185900 24500 186000 24600
rect 185900 24600 186000 24700
rect 185900 24700 186000 24800
rect 185900 24800 186000 24900
rect 185900 24900 186000 25000
rect 185900 25000 186000 25100
rect 185900 25100 186000 25200
rect 185900 25200 186000 25300
rect 185900 25300 186000 25400
rect 185900 25400 186000 25500
rect 185900 25500 186000 25600
rect 185900 25600 186000 25700
rect 185900 25700 186000 25800
rect 185900 25800 186000 25900
rect 185900 25900 186000 26000
rect 185900 26000 186000 26100
rect 185900 26100 186000 26200
rect 185900 26200 186000 26300
rect 185900 26300 186000 26400
rect 185900 26400 186000 26500
rect 185900 26500 186000 26600
rect 185900 26600 186000 26700
rect 185900 26700 186000 26800
rect 185900 26800 186000 26900
rect 185900 26900 186000 27000
rect 185900 27000 186000 27100
rect 185900 27100 186000 27200
rect 185900 27200 186000 27300
rect 185900 27300 186000 27400
rect 185900 27400 186000 27500
rect 185900 27500 186000 27600
rect 185900 27600 186000 27700
rect 185900 27700 186000 27800
rect 185900 27800 186000 27900
rect 185900 27900 186000 28000
rect 185900 28000 186000 28100
rect 185900 28100 186000 28200
rect 185900 28200 186000 28300
rect 185900 28300 186000 28400
rect 185900 28400 186000 28500
rect 185900 28500 186000 28600
rect 185900 28600 186000 28700
rect 185900 28700 186000 28800
rect 185900 28800 186000 28900
rect 185900 28900 186000 29000
rect 185900 29000 186000 29100
rect 185900 29100 186000 29200
rect 185900 29200 186000 29300
rect 185900 29300 186000 29400
rect 185900 29400 186000 29500
rect 185900 29500 186000 29600
rect 185900 29600 186000 29700
rect 185900 29700 186000 29800
rect 185900 29800 186000 29900
rect 185900 29900 186000 30000
rect 185900 30000 186000 30100
rect 185900 30100 186000 30200
rect 185900 30200 186000 30300
rect 185900 30300 186000 30400
rect 185900 30400 186000 30500
rect 185900 30500 186000 30600
rect 185900 30600 186000 30700
rect 185900 30700 186000 30800
rect 185900 30800 186000 30900
rect 185900 30900 186000 31000
rect 185900 31000 186000 31100
rect 185900 31100 186000 31200
rect 185900 31200 186000 31300
rect 185900 31300 186000 31400
rect 185900 31400 186000 31500
rect 185900 31500 186000 31600
rect 185900 31600 186000 31700
rect 185900 31700 186000 31800
rect 185900 31800 186000 31900
rect 185900 31900 186000 32000
rect 185900 35300 186000 35400
rect 185900 35400 186000 35500
rect 185900 35500 186000 35600
rect 185900 35600 186000 35700
rect 185900 35700 186000 35800
rect 185900 35800 186000 35900
rect 185900 35900 186000 36000
rect 185900 36000 186000 36100
rect 185900 36100 186000 36200
rect 185900 36200 186000 36300
rect 185900 36300 186000 36400
rect 185900 36400 186000 36500
rect 185900 36500 186000 36600
rect 185900 36600 186000 36700
rect 185900 36700 186000 36800
rect 185900 36800 186000 36900
rect 185900 36900 186000 37000
rect 185900 37000 186000 37100
rect 185900 37100 186000 37200
rect 185900 37200 186000 37300
rect 185900 37300 186000 37400
rect 185900 37400 186000 37500
rect 185900 37500 186000 37600
rect 185900 37600 186000 37700
rect 185900 37700 186000 37800
rect 185900 37800 186000 37900
rect 185900 37900 186000 38000
rect 186000 21300 186100 21400
rect 186000 21400 186100 21500
rect 186000 21500 186100 21600
rect 186000 21600 186100 21700
rect 186000 21700 186100 21800
rect 186000 21800 186100 21900
rect 186000 21900 186100 22000
rect 186000 22000 186100 22100
rect 186000 22100 186100 22200
rect 186000 22200 186100 22300
rect 186000 22300 186100 22400
rect 186000 22400 186100 22500
rect 186000 22500 186100 22600
rect 186000 22600 186100 22700
rect 186000 22700 186100 22800
rect 186000 22800 186100 22900
rect 186000 22900 186100 23000
rect 186000 23000 186100 23100
rect 186000 23100 186100 23200
rect 186000 23200 186100 23300
rect 186000 23300 186100 23400
rect 186000 23400 186100 23500
rect 186000 23500 186100 23600
rect 186000 23600 186100 23700
rect 186000 23700 186100 23800
rect 186000 23800 186100 23900
rect 186000 23900 186100 24000
rect 186000 24000 186100 24100
rect 186000 24100 186100 24200
rect 186000 24200 186100 24300
rect 186000 24300 186100 24400
rect 186000 24400 186100 24500
rect 186000 24500 186100 24600
rect 186000 24600 186100 24700
rect 186000 24700 186100 24800
rect 186000 24800 186100 24900
rect 186000 24900 186100 25000
rect 186000 25000 186100 25100
rect 186000 25100 186100 25200
rect 186000 25200 186100 25300
rect 186000 25300 186100 25400
rect 186000 25400 186100 25500
rect 186000 25500 186100 25600
rect 186000 25600 186100 25700
rect 186000 25700 186100 25800
rect 186000 25800 186100 25900
rect 186000 25900 186100 26000
rect 186000 26000 186100 26100
rect 186000 26100 186100 26200
rect 186000 26200 186100 26300
rect 186000 26300 186100 26400
rect 186000 26400 186100 26500
rect 186000 26500 186100 26600
rect 186000 26600 186100 26700
rect 186000 26700 186100 26800
rect 186000 26800 186100 26900
rect 186000 26900 186100 27000
rect 186000 27000 186100 27100
rect 186000 27100 186100 27200
rect 186000 27200 186100 27300
rect 186000 27300 186100 27400
rect 186000 27400 186100 27500
rect 186000 27500 186100 27600
rect 186000 27600 186100 27700
rect 186000 27700 186100 27800
rect 186000 27800 186100 27900
rect 186000 27900 186100 28000
rect 186000 28000 186100 28100
rect 186000 28100 186100 28200
rect 186000 28200 186100 28300
rect 186000 28300 186100 28400
rect 186000 28400 186100 28500
rect 186000 28500 186100 28600
rect 186000 28600 186100 28700
rect 186000 28700 186100 28800
rect 186000 28800 186100 28900
rect 186000 28900 186100 29000
rect 186000 29000 186100 29100
rect 186000 29100 186100 29200
rect 186000 29200 186100 29300
rect 186000 29300 186100 29400
rect 186000 29400 186100 29500
rect 186000 29500 186100 29600
rect 186000 29600 186100 29700
rect 186000 29700 186100 29800
rect 186000 29800 186100 29900
rect 186000 29900 186100 30000
rect 186000 30000 186100 30100
rect 186000 30100 186100 30200
rect 186000 30200 186100 30300
rect 186000 30300 186100 30400
rect 186000 30400 186100 30500
rect 186000 30500 186100 30600
rect 186000 30600 186100 30700
rect 186000 30700 186100 30800
rect 186000 30800 186100 30900
rect 186000 30900 186100 31000
rect 186000 31000 186100 31100
rect 186000 31100 186100 31200
rect 186000 31200 186100 31300
rect 186000 31300 186100 31400
rect 186000 31400 186100 31500
rect 186000 31500 186100 31600
rect 186000 31600 186100 31700
rect 186000 31700 186100 31800
rect 186000 31800 186100 31900
rect 186000 31900 186100 32000
rect 186000 32000 186100 32100
rect 186000 32100 186100 32200
rect 186000 35200 186100 35300
rect 186000 35300 186100 35400
rect 186000 35400 186100 35500
rect 186000 35500 186100 35600
rect 186000 35600 186100 35700
rect 186000 35700 186100 35800
rect 186000 35800 186100 35900
rect 186000 35900 186100 36000
rect 186000 36000 186100 36100
rect 186000 36100 186100 36200
rect 186000 36200 186100 36300
rect 186000 36300 186100 36400
rect 186000 36400 186100 36500
rect 186000 36500 186100 36600
rect 186000 36600 186100 36700
rect 186000 36700 186100 36800
rect 186000 36800 186100 36900
rect 186000 36900 186100 37000
rect 186000 37000 186100 37100
rect 186000 37100 186100 37200
rect 186000 37200 186100 37300
rect 186000 37300 186100 37400
rect 186000 37400 186100 37500
rect 186000 37500 186100 37600
rect 186000 37600 186100 37700
rect 186000 37700 186100 37800
rect 186000 37800 186100 37900
rect 186000 37900 186100 38000
rect 186000 38000 186100 38100
rect 186000 38100 186100 38200
rect 186100 21200 186200 21300
rect 186100 21300 186200 21400
rect 186100 21400 186200 21500
rect 186100 21500 186200 21600
rect 186100 21600 186200 21700
rect 186100 21700 186200 21800
rect 186100 21800 186200 21900
rect 186100 21900 186200 22000
rect 186100 22000 186200 22100
rect 186100 22100 186200 22200
rect 186100 22200 186200 22300
rect 186100 22300 186200 22400
rect 186100 22400 186200 22500
rect 186100 22500 186200 22600
rect 186100 22600 186200 22700
rect 186100 22700 186200 22800
rect 186100 22800 186200 22900
rect 186100 22900 186200 23000
rect 186100 23000 186200 23100
rect 186100 23100 186200 23200
rect 186100 23200 186200 23300
rect 186100 23300 186200 23400
rect 186100 23400 186200 23500
rect 186100 23500 186200 23600
rect 186100 23600 186200 23700
rect 186100 23700 186200 23800
rect 186100 23800 186200 23900
rect 186100 23900 186200 24000
rect 186100 24000 186200 24100
rect 186100 24100 186200 24200
rect 186100 24200 186200 24300
rect 186100 24300 186200 24400
rect 186100 24400 186200 24500
rect 186100 24500 186200 24600
rect 186100 24600 186200 24700
rect 186100 24700 186200 24800
rect 186100 24800 186200 24900
rect 186100 24900 186200 25000
rect 186100 25000 186200 25100
rect 186100 25100 186200 25200
rect 186100 25200 186200 25300
rect 186100 25300 186200 25400
rect 186100 25400 186200 25500
rect 186100 25500 186200 25600
rect 186100 25600 186200 25700
rect 186100 25700 186200 25800
rect 186100 25800 186200 25900
rect 186100 25900 186200 26000
rect 186100 26000 186200 26100
rect 186100 26100 186200 26200
rect 186100 26200 186200 26300
rect 186100 26300 186200 26400
rect 186100 26400 186200 26500
rect 186100 26500 186200 26600
rect 186100 26600 186200 26700
rect 186100 26700 186200 26800
rect 186100 26800 186200 26900
rect 186100 26900 186200 27000
rect 186100 27000 186200 27100
rect 186100 27100 186200 27200
rect 186100 27200 186200 27300
rect 186100 27300 186200 27400
rect 186100 27400 186200 27500
rect 186100 27500 186200 27600
rect 186100 27600 186200 27700
rect 186100 27700 186200 27800
rect 186100 27800 186200 27900
rect 186100 27900 186200 28000
rect 186100 28000 186200 28100
rect 186100 28100 186200 28200
rect 186100 28200 186200 28300
rect 186100 28300 186200 28400
rect 186100 28400 186200 28500
rect 186100 28500 186200 28600
rect 186100 28600 186200 28700
rect 186100 28700 186200 28800
rect 186100 28800 186200 28900
rect 186100 28900 186200 29000
rect 186100 29000 186200 29100
rect 186100 29100 186200 29200
rect 186100 29200 186200 29300
rect 186100 29300 186200 29400
rect 186100 29400 186200 29500
rect 186100 29500 186200 29600
rect 186100 29600 186200 29700
rect 186100 29700 186200 29800
rect 186100 29800 186200 29900
rect 186100 29900 186200 30000
rect 186100 30000 186200 30100
rect 186100 30100 186200 30200
rect 186100 30200 186200 30300
rect 186100 30300 186200 30400
rect 186100 30400 186200 30500
rect 186100 30500 186200 30600
rect 186100 30600 186200 30700
rect 186100 30700 186200 30800
rect 186100 30800 186200 30900
rect 186100 30900 186200 31000
rect 186100 31000 186200 31100
rect 186100 31100 186200 31200
rect 186100 31200 186200 31300
rect 186100 31300 186200 31400
rect 186100 31400 186200 31500
rect 186100 31500 186200 31600
rect 186100 31600 186200 31700
rect 186100 31700 186200 31800
rect 186100 31800 186200 31900
rect 186100 31900 186200 32000
rect 186100 32000 186200 32100
rect 186100 32100 186200 32200
rect 186100 32200 186200 32300
rect 186100 32300 186200 32400
rect 186100 35100 186200 35200
rect 186100 35200 186200 35300
rect 186100 35300 186200 35400
rect 186100 35400 186200 35500
rect 186100 35500 186200 35600
rect 186100 35600 186200 35700
rect 186100 35700 186200 35800
rect 186100 35800 186200 35900
rect 186100 35900 186200 36000
rect 186100 36000 186200 36100
rect 186100 36100 186200 36200
rect 186100 36200 186200 36300
rect 186100 36300 186200 36400
rect 186100 36400 186200 36500
rect 186100 36500 186200 36600
rect 186100 36600 186200 36700
rect 186100 36700 186200 36800
rect 186100 36800 186200 36900
rect 186100 36900 186200 37000
rect 186100 37000 186200 37100
rect 186100 37100 186200 37200
rect 186100 37200 186200 37300
rect 186100 37300 186200 37400
rect 186100 37400 186200 37500
rect 186100 37500 186200 37600
rect 186100 37600 186200 37700
rect 186100 37700 186200 37800
rect 186100 37800 186200 37900
rect 186100 37900 186200 38000
rect 186100 38000 186200 38100
rect 186100 38100 186200 38200
rect 186100 38200 186200 38300
rect 186200 21200 186300 21300
rect 186200 21300 186300 21400
rect 186200 21400 186300 21500
rect 186200 21500 186300 21600
rect 186200 21600 186300 21700
rect 186200 21700 186300 21800
rect 186200 21800 186300 21900
rect 186200 21900 186300 22000
rect 186200 22000 186300 22100
rect 186200 22100 186300 22200
rect 186200 22200 186300 22300
rect 186200 22300 186300 22400
rect 186200 22400 186300 22500
rect 186200 22500 186300 22600
rect 186200 22600 186300 22700
rect 186200 22700 186300 22800
rect 186200 22800 186300 22900
rect 186200 22900 186300 23000
rect 186200 23000 186300 23100
rect 186200 23100 186300 23200
rect 186200 23200 186300 23300
rect 186200 23300 186300 23400
rect 186200 23400 186300 23500
rect 186200 23500 186300 23600
rect 186200 23600 186300 23700
rect 186200 23700 186300 23800
rect 186200 23800 186300 23900
rect 186200 23900 186300 24000
rect 186200 24000 186300 24100
rect 186200 24100 186300 24200
rect 186200 24200 186300 24300
rect 186200 24300 186300 24400
rect 186200 24400 186300 24500
rect 186200 24500 186300 24600
rect 186200 24600 186300 24700
rect 186200 24700 186300 24800
rect 186200 24800 186300 24900
rect 186200 24900 186300 25000
rect 186200 25000 186300 25100
rect 186200 25100 186300 25200
rect 186200 25200 186300 25300
rect 186200 25300 186300 25400
rect 186200 25400 186300 25500
rect 186200 25500 186300 25600
rect 186200 25600 186300 25700
rect 186200 25700 186300 25800
rect 186200 25800 186300 25900
rect 186200 25900 186300 26000
rect 186200 26000 186300 26100
rect 186200 26100 186300 26200
rect 186200 26200 186300 26300
rect 186200 26300 186300 26400
rect 186200 26400 186300 26500
rect 186200 26500 186300 26600
rect 186200 26600 186300 26700
rect 186200 26700 186300 26800
rect 186200 26800 186300 26900
rect 186200 26900 186300 27000
rect 186200 27000 186300 27100
rect 186200 27100 186300 27200
rect 186200 27200 186300 27300
rect 186200 27300 186300 27400
rect 186200 27400 186300 27500
rect 186200 27500 186300 27600
rect 186200 27600 186300 27700
rect 186200 27700 186300 27800
rect 186200 27800 186300 27900
rect 186200 27900 186300 28000
rect 186200 28000 186300 28100
rect 186200 28100 186300 28200
rect 186200 28200 186300 28300
rect 186200 28300 186300 28400
rect 186200 28400 186300 28500
rect 186200 28500 186300 28600
rect 186200 28600 186300 28700
rect 186200 28700 186300 28800
rect 186200 28800 186300 28900
rect 186200 28900 186300 29000
rect 186200 29000 186300 29100
rect 186200 29100 186300 29200
rect 186200 29200 186300 29300
rect 186200 29300 186300 29400
rect 186200 29400 186300 29500
rect 186200 29500 186300 29600
rect 186200 29600 186300 29700
rect 186200 29700 186300 29800
rect 186200 29800 186300 29900
rect 186200 29900 186300 30000
rect 186200 30000 186300 30100
rect 186200 30100 186300 30200
rect 186200 30200 186300 30300
rect 186200 30300 186300 30400
rect 186200 30400 186300 30500
rect 186200 30500 186300 30600
rect 186200 30600 186300 30700
rect 186200 30700 186300 30800
rect 186200 30800 186300 30900
rect 186200 30900 186300 31000
rect 186200 31000 186300 31100
rect 186200 31100 186300 31200
rect 186200 31200 186300 31300
rect 186200 31300 186300 31400
rect 186200 31400 186300 31500
rect 186200 31500 186300 31600
rect 186200 31600 186300 31700
rect 186200 31700 186300 31800
rect 186200 31800 186300 31900
rect 186200 31900 186300 32000
rect 186200 32000 186300 32100
rect 186200 32100 186300 32200
rect 186200 32200 186300 32300
rect 186200 32300 186300 32400
rect 186200 32400 186300 32500
rect 186200 35000 186300 35100
rect 186200 35100 186300 35200
rect 186200 35200 186300 35300
rect 186200 35300 186300 35400
rect 186200 35400 186300 35500
rect 186200 35500 186300 35600
rect 186200 35600 186300 35700
rect 186200 35700 186300 35800
rect 186200 35800 186300 35900
rect 186200 35900 186300 36000
rect 186200 36000 186300 36100
rect 186200 36100 186300 36200
rect 186200 36200 186300 36300
rect 186200 36300 186300 36400
rect 186200 36400 186300 36500
rect 186200 36500 186300 36600
rect 186200 36600 186300 36700
rect 186200 36700 186300 36800
rect 186200 36800 186300 36900
rect 186200 36900 186300 37000
rect 186200 37000 186300 37100
rect 186200 37100 186300 37200
rect 186200 37200 186300 37300
rect 186200 37300 186300 37400
rect 186200 37400 186300 37500
rect 186200 37500 186300 37600
rect 186200 37600 186300 37700
rect 186200 37700 186300 37800
rect 186200 37800 186300 37900
rect 186200 37900 186300 38000
rect 186200 38000 186300 38100
rect 186200 38100 186300 38200
rect 186200 38200 186300 38300
rect 186200 38300 186300 38400
rect 186300 21200 186400 21300
rect 186300 21300 186400 21400
rect 186300 21400 186400 21500
rect 186300 21500 186400 21600
rect 186300 21600 186400 21700
rect 186300 21700 186400 21800
rect 186300 21800 186400 21900
rect 186300 21900 186400 22000
rect 186300 22000 186400 22100
rect 186300 22100 186400 22200
rect 186300 22200 186400 22300
rect 186300 22300 186400 22400
rect 186300 22400 186400 22500
rect 186300 22500 186400 22600
rect 186300 22600 186400 22700
rect 186300 22700 186400 22800
rect 186300 22800 186400 22900
rect 186300 22900 186400 23000
rect 186300 23000 186400 23100
rect 186300 23100 186400 23200
rect 186300 23200 186400 23300
rect 186300 23300 186400 23400
rect 186300 23400 186400 23500
rect 186300 23500 186400 23600
rect 186300 23600 186400 23700
rect 186300 23700 186400 23800
rect 186300 23800 186400 23900
rect 186300 23900 186400 24000
rect 186300 24000 186400 24100
rect 186300 24100 186400 24200
rect 186300 24200 186400 24300
rect 186300 24300 186400 24400
rect 186300 24400 186400 24500
rect 186300 24500 186400 24600
rect 186300 24600 186400 24700
rect 186300 24700 186400 24800
rect 186300 24800 186400 24900
rect 186300 24900 186400 25000
rect 186300 25000 186400 25100
rect 186300 25100 186400 25200
rect 186300 25200 186400 25300
rect 186300 25300 186400 25400
rect 186300 25400 186400 25500
rect 186300 25500 186400 25600
rect 186300 25600 186400 25700
rect 186300 25700 186400 25800
rect 186300 25800 186400 25900
rect 186300 25900 186400 26000
rect 186300 26000 186400 26100
rect 186300 26100 186400 26200
rect 186300 26200 186400 26300
rect 186300 26300 186400 26400
rect 186300 26400 186400 26500
rect 186300 26500 186400 26600
rect 186300 26600 186400 26700
rect 186300 26700 186400 26800
rect 186300 26800 186400 26900
rect 186300 26900 186400 27000
rect 186300 27000 186400 27100
rect 186300 27100 186400 27200
rect 186300 27200 186400 27300
rect 186300 27300 186400 27400
rect 186300 27400 186400 27500
rect 186300 27500 186400 27600
rect 186300 27600 186400 27700
rect 186300 27700 186400 27800
rect 186300 27800 186400 27900
rect 186300 27900 186400 28000
rect 186300 28000 186400 28100
rect 186300 28100 186400 28200
rect 186300 28200 186400 28300
rect 186300 28300 186400 28400
rect 186300 28400 186400 28500
rect 186300 28500 186400 28600
rect 186300 28600 186400 28700
rect 186300 28700 186400 28800
rect 186300 28800 186400 28900
rect 186300 28900 186400 29000
rect 186300 29000 186400 29100
rect 186300 29100 186400 29200
rect 186300 29200 186400 29300
rect 186300 29300 186400 29400
rect 186300 29400 186400 29500
rect 186300 29500 186400 29600
rect 186300 29600 186400 29700
rect 186300 29700 186400 29800
rect 186300 29800 186400 29900
rect 186300 29900 186400 30000
rect 186300 30000 186400 30100
rect 186300 30100 186400 30200
rect 186300 30200 186400 30300
rect 186300 30300 186400 30400
rect 186300 30400 186400 30500
rect 186300 30500 186400 30600
rect 186300 30600 186400 30700
rect 186300 30700 186400 30800
rect 186300 30800 186400 30900
rect 186300 30900 186400 31000
rect 186300 31000 186400 31100
rect 186300 31100 186400 31200
rect 186300 31200 186400 31300
rect 186300 31300 186400 31400
rect 186300 31400 186400 31500
rect 186300 31500 186400 31600
rect 186300 31600 186400 31700
rect 186300 31700 186400 31800
rect 186300 31800 186400 31900
rect 186300 31900 186400 32000
rect 186300 32000 186400 32100
rect 186300 32100 186400 32200
rect 186300 32200 186400 32300
rect 186300 32300 186400 32400
rect 186300 32400 186400 32500
rect 186300 32500 186400 32600
rect 186300 32600 186400 32700
rect 186300 34900 186400 35000
rect 186300 35000 186400 35100
rect 186300 35100 186400 35200
rect 186300 35200 186400 35300
rect 186300 35300 186400 35400
rect 186300 35400 186400 35500
rect 186300 35500 186400 35600
rect 186300 35600 186400 35700
rect 186300 35700 186400 35800
rect 186300 35800 186400 35900
rect 186300 35900 186400 36000
rect 186300 36000 186400 36100
rect 186300 36100 186400 36200
rect 186300 36200 186400 36300
rect 186300 36300 186400 36400
rect 186300 36400 186400 36500
rect 186300 36500 186400 36600
rect 186300 36600 186400 36700
rect 186300 36700 186400 36800
rect 186300 36800 186400 36900
rect 186300 36900 186400 37000
rect 186300 37000 186400 37100
rect 186300 37100 186400 37200
rect 186300 37200 186400 37300
rect 186300 37300 186400 37400
rect 186300 37400 186400 37500
rect 186300 37500 186400 37600
rect 186300 37600 186400 37700
rect 186300 37700 186400 37800
rect 186300 37800 186400 37900
rect 186300 37900 186400 38000
rect 186300 38000 186400 38100
rect 186300 38100 186400 38200
rect 186300 38200 186400 38300
rect 186300 38300 186400 38400
rect 186300 38400 186400 38500
rect 186400 21200 186500 21300
rect 186400 21300 186500 21400
rect 186400 21400 186500 21500
rect 186400 21500 186500 21600
rect 186400 21600 186500 21700
rect 186400 21700 186500 21800
rect 186400 21800 186500 21900
rect 186400 21900 186500 22000
rect 186400 22000 186500 22100
rect 186400 22100 186500 22200
rect 186400 22200 186500 22300
rect 186400 22300 186500 22400
rect 186400 22400 186500 22500
rect 186400 22500 186500 22600
rect 186400 22600 186500 22700
rect 186400 22700 186500 22800
rect 186400 22800 186500 22900
rect 186400 22900 186500 23000
rect 186400 23000 186500 23100
rect 186400 23100 186500 23200
rect 186400 23200 186500 23300
rect 186400 23300 186500 23400
rect 186400 23400 186500 23500
rect 186400 23500 186500 23600
rect 186400 23600 186500 23700
rect 186400 23700 186500 23800
rect 186400 23800 186500 23900
rect 186400 23900 186500 24000
rect 186400 24000 186500 24100
rect 186400 24100 186500 24200
rect 186400 24200 186500 24300
rect 186400 24300 186500 24400
rect 186400 24400 186500 24500
rect 186400 24500 186500 24600
rect 186400 24600 186500 24700
rect 186400 24700 186500 24800
rect 186400 24800 186500 24900
rect 186400 24900 186500 25000
rect 186400 25000 186500 25100
rect 186400 25100 186500 25200
rect 186400 25200 186500 25300
rect 186400 25300 186500 25400
rect 186400 25400 186500 25500
rect 186400 25500 186500 25600
rect 186400 25600 186500 25700
rect 186400 25700 186500 25800
rect 186400 25800 186500 25900
rect 186400 25900 186500 26000
rect 186400 26000 186500 26100
rect 186400 26100 186500 26200
rect 186400 26200 186500 26300
rect 186400 26300 186500 26400
rect 186400 26400 186500 26500
rect 186400 26500 186500 26600
rect 186400 26600 186500 26700
rect 186400 26700 186500 26800
rect 186400 26800 186500 26900
rect 186400 26900 186500 27000
rect 186400 27000 186500 27100
rect 186400 27100 186500 27200
rect 186400 27200 186500 27300
rect 186400 27300 186500 27400
rect 186400 27400 186500 27500
rect 186400 27500 186500 27600
rect 186400 27600 186500 27700
rect 186400 27700 186500 27800
rect 186400 27800 186500 27900
rect 186400 27900 186500 28000
rect 186400 28000 186500 28100
rect 186400 28100 186500 28200
rect 186400 28200 186500 28300
rect 186400 28300 186500 28400
rect 186400 28400 186500 28500
rect 186400 28500 186500 28600
rect 186400 28600 186500 28700
rect 186400 28700 186500 28800
rect 186400 28800 186500 28900
rect 186400 28900 186500 29000
rect 186400 29000 186500 29100
rect 186400 29100 186500 29200
rect 186400 29200 186500 29300
rect 186400 29300 186500 29400
rect 186400 29400 186500 29500
rect 186400 29500 186500 29600
rect 186400 29600 186500 29700
rect 186400 29700 186500 29800
rect 186400 29800 186500 29900
rect 186400 29900 186500 30000
rect 186400 30000 186500 30100
rect 186400 30100 186500 30200
rect 186400 30200 186500 30300
rect 186400 30300 186500 30400
rect 186400 30400 186500 30500
rect 186400 30500 186500 30600
rect 186400 30600 186500 30700
rect 186400 30700 186500 30800
rect 186400 30800 186500 30900
rect 186400 30900 186500 31000
rect 186400 31000 186500 31100
rect 186400 31100 186500 31200
rect 186400 31200 186500 31300
rect 186400 31300 186500 31400
rect 186400 31400 186500 31500
rect 186400 31500 186500 31600
rect 186400 31600 186500 31700
rect 186400 31700 186500 31800
rect 186400 31800 186500 31900
rect 186400 31900 186500 32000
rect 186400 32000 186500 32100
rect 186400 32100 186500 32200
rect 186400 32200 186500 32300
rect 186400 32300 186500 32400
rect 186400 32400 186500 32500
rect 186400 32500 186500 32600
rect 186400 32600 186500 32700
rect 186400 32700 186500 32800
rect 186400 34800 186500 34900
rect 186400 34900 186500 35000
rect 186400 35000 186500 35100
rect 186400 35100 186500 35200
rect 186400 35200 186500 35300
rect 186400 35300 186500 35400
rect 186400 35400 186500 35500
rect 186400 35500 186500 35600
rect 186400 35600 186500 35700
rect 186400 35700 186500 35800
rect 186400 35800 186500 35900
rect 186400 35900 186500 36000
rect 186400 36000 186500 36100
rect 186400 36100 186500 36200
rect 186400 36200 186500 36300
rect 186400 36300 186500 36400
rect 186400 36400 186500 36500
rect 186400 36500 186500 36600
rect 186400 36600 186500 36700
rect 186400 36700 186500 36800
rect 186400 36800 186500 36900
rect 186400 36900 186500 37000
rect 186400 37000 186500 37100
rect 186400 37100 186500 37200
rect 186400 37200 186500 37300
rect 186400 37300 186500 37400
rect 186400 37400 186500 37500
rect 186400 37500 186500 37600
rect 186400 37600 186500 37700
rect 186400 37700 186500 37800
rect 186400 37800 186500 37900
rect 186400 37900 186500 38000
rect 186400 38000 186500 38100
rect 186400 38100 186500 38200
rect 186400 38200 186500 38300
rect 186400 38300 186500 38400
rect 186400 38400 186500 38500
rect 186400 38500 186500 38600
rect 186500 21200 186600 21300
rect 186500 21300 186600 21400
rect 186500 21400 186600 21500
rect 186500 21500 186600 21600
rect 186500 21600 186600 21700
rect 186500 21700 186600 21800
rect 186500 21800 186600 21900
rect 186500 21900 186600 22000
rect 186500 22000 186600 22100
rect 186500 22100 186600 22200
rect 186500 22200 186600 22300
rect 186500 22300 186600 22400
rect 186500 22400 186600 22500
rect 186500 22500 186600 22600
rect 186500 22600 186600 22700
rect 186500 22700 186600 22800
rect 186500 22800 186600 22900
rect 186500 22900 186600 23000
rect 186500 23000 186600 23100
rect 186500 23100 186600 23200
rect 186500 23200 186600 23300
rect 186500 23300 186600 23400
rect 186500 23400 186600 23500
rect 186500 23500 186600 23600
rect 186500 23600 186600 23700
rect 186500 23700 186600 23800
rect 186500 23800 186600 23900
rect 186500 23900 186600 24000
rect 186500 24000 186600 24100
rect 186500 24100 186600 24200
rect 186500 24200 186600 24300
rect 186500 24300 186600 24400
rect 186500 24400 186600 24500
rect 186500 24500 186600 24600
rect 186500 24600 186600 24700
rect 186500 24700 186600 24800
rect 186500 24800 186600 24900
rect 186500 24900 186600 25000
rect 186500 25000 186600 25100
rect 186500 25100 186600 25200
rect 186500 25200 186600 25300
rect 186500 25300 186600 25400
rect 186500 25400 186600 25500
rect 186500 25500 186600 25600
rect 186500 25600 186600 25700
rect 186500 25700 186600 25800
rect 186500 25800 186600 25900
rect 186500 25900 186600 26000
rect 186500 26000 186600 26100
rect 186500 26100 186600 26200
rect 186500 26200 186600 26300
rect 186500 26300 186600 26400
rect 186500 26400 186600 26500
rect 186500 26500 186600 26600
rect 186500 26600 186600 26700
rect 186500 26700 186600 26800
rect 186500 26800 186600 26900
rect 186500 26900 186600 27000
rect 186500 27000 186600 27100
rect 186500 27100 186600 27200
rect 186500 27200 186600 27300
rect 186500 27300 186600 27400
rect 186500 27400 186600 27500
rect 186500 27500 186600 27600
rect 186500 27600 186600 27700
rect 186500 27700 186600 27800
rect 186500 27800 186600 27900
rect 186500 27900 186600 28000
rect 186500 28000 186600 28100
rect 186500 28100 186600 28200
rect 186500 28200 186600 28300
rect 186500 28300 186600 28400
rect 186500 28400 186600 28500
rect 186500 28500 186600 28600
rect 186500 28600 186600 28700
rect 186500 28700 186600 28800
rect 186500 28800 186600 28900
rect 186500 28900 186600 29000
rect 186500 29000 186600 29100
rect 186500 29100 186600 29200
rect 186500 29200 186600 29300
rect 186500 29300 186600 29400
rect 186500 29400 186600 29500
rect 186500 29500 186600 29600
rect 186500 29600 186600 29700
rect 186500 29700 186600 29800
rect 186500 29800 186600 29900
rect 186500 29900 186600 30000
rect 186500 30000 186600 30100
rect 186500 30100 186600 30200
rect 186500 30200 186600 30300
rect 186500 30300 186600 30400
rect 186500 30400 186600 30500
rect 186500 30500 186600 30600
rect 186500 30600 186600 30700
rect 186500 30700 186600 30800
rect 186500 30800 186600 30900
rect 186500 30900 186600 31000
rect 186500 31000 186600 31100
rect 186500 31100 186600 31200
rect 186500 31200 186600 31300
rect 186500 31300 186600 31400
rect 186500 31400 186600 31500
rect 186500 31500 186600 31600
rect 186500 31600 186600 31700
rect 186500 31700 186600 31800
rect 186500 31800 186600 31900
rect 186500 31900 186600 32000
rect 186500 32000 186600 32100
rect 186500 32100 186600 32200
rect 186500 32200 186600 32300
rect 186500 32300 186600 32400
rect 186500 32400 186600 32500
rect 186500 32500 186600 32600
rect 186500 32600 186600 32700
rect 186500 32700 186600 32800
rect 186500 32800 186600 32900
rect 186500 34700 186600 34800
rect 186500 34800 186600 34900
rect 186500 34900 186600 35000
rect 186500 35000 186600 35100
rect 186500 35100 186600 35200
rect 186500 35200 186600 35300
rect 186500 35300 186600 35400
rect 186500 35400 186600 35500
rect 186500 35500 186600 35600
rect 186500 35600 186600 35700
rect 186500 35700 186600 35800
rect 186500 35800 186600 35900
rect 186500 35900 186600 36000
rect 186500 36000 186600 36100
rect 186500 36100 186600 36200
rect 186500 36200 186600 36300
rect 186500 36300 186600 36400
rect 186500 36400 186600 36500
rect 186500 36500 186600 36600
rect 186500 36600 186600 36700
rect 186500 36700 186600 36800
rect 186500 36800 186600 36900
rect 186500 36900 186600 37000
rect 186500 37000 186600 37100
rect 186500 37100 186600 37200
rect 186500 37200 186600 37300
rect 186500 37300 186600 37400
rect 186500 37400 186600 37500
rect 186500 37500 186600 37600
rect 186500 37600 186600 37700
rect 186500 37700 186600 37800
rect 186500 37800 186600 37900
rect 186500 37900 186600 38000
rect 186500 38000 186600 38100
rect 186500 38100 186600 38200
rect 186500 38200 186600 38300
rect 186500 38300 186600 38400
rect 186500 38400 186600 38500
rect 186500 38500 186600 38600
rect 186500 38600 186600 38700
rect 186600 21200 186700 21300
rect 186600 21300 186700 21400
rect 186600 21400 186700 21500
rect 186600 21500 186700 21600
rect 186600 21600 186700 21700
rect 186600 21700 186700 21800
rect 186600 21800 186700 21900
rect 186600 21900 186700 22000
rect 186600 22000 186700 22100
rect 186600 22100 186700 22200
rect 186600 22200 186700 22300
rect 186600 22300 186700 22400
rect 186600 22400 186700 22500
rect 186600 22500 186700 22600
rect 186600 22600 186700 22700
rect 186600 22700 186700 22800
rect 186600 22800 186700 22900
rect 186600 22900 186700 23000
rect 186600 23000 186700 23100
rect 186600 23100 186700 23200
rect 186600 23200 186700 23300
rect 186600 23300 186700 23400
rect 186600 23400 186700 23500
rect 186600 23500 186700 23600
rect 186600 23600 186700 23700
rect 186600 23700 186700 23800
rect 186600 23800 186700 23900
rect 186600 23900 186700 24000
rect 186600 24000 186700 24100
rect 186600 24100 186700 24200
rect 186600 24200 186700 24300
rect 186600 24300 186700 24400
rect 186600 24400 186700 24500
rect 186600 24500 186700 24600
rect 186600 24600 186700 24700
rect 186600 24700 186700 24800
rect 186600 24800 186700 24900
rect 186600 24900 186700 25000
rect 186600 25000 186700 25100
rect 186600 25100 186700 25200
rect 186600 25200 186700 25300
rect 186600 25300 186700 25400
rect 186600 25400 186700 25500
rect 186600 25500 186700 25600
rect 186600 25600 186700 25700
rect 186600 25700 186700 25800
rect 186600 25800 186700 25900
rect 186600 25900 186700 26000
rect 186600 26000 186700 26100
rect 186600 26100 186700 26200
rect 186600 26200 186700 26300
rect 186600 26300 186700 26400
rect 186600 26400 186700 26500
rect 186600 26500 186700 26600
rect 186600 26600 186700 26700
rect 186600 26700 186700 26800
rect 186600 26800 186700 26900
rect 186600 26900 186700 27000
rect 186600 27000 186700 27100
rect 186600 27100 186700 27200
rect 186600 27200 186700 27300
rect 186600 27300 186700 27400
rect 186600 27400 186700 27500
rect 186600 27500 186700 27600
rect 186600 27600 186700 27700
rect 186600 27700 186700 27800
rect 186600 27800 186700 27900
rect 186600 27900 186700 28000
rect 186600 28000 186700 28100
rect 186600 28100 186700 28200
rect 186600 28200 186700 28300
rect 186600 28300 186700 28400
rect 186600 28400 186700 28500
rect 186600 28500 186700 28600
rect 186600 28600 186700 28700
rect 186600 28700 186700 28800
rect 186600 28800 186700 28900
rect 186600 28900 186700 29000
rect 186600 29000 186700 29100
rect 186600 29100 186700 29200
rect 186600 29200 186700 29300
rect 186600 29300 186700 29400
rect 186600 29400 186700 29500
rect 186600 29500 186700 29600
rect 186600 29600 186700 29700
rect 186600 29700 186700 29800
rect 186600 29800 186700 29900
rect 186600 29900 186700 30000
rect 186600 30000 186700 30100
rect 186600 30100 186700 30200
rect 186600 30200 186700 30300
rect 186600 30300 186700 30400
rect 186600 30400 186700 30500
rect 186600 30500 186700 30600
rect 186600 30600 186700 30700
rect 186600 30700 186700 30800
rect 186600 30800 186700 30900
rect 186600 30900 186700 31000
rect 186600 31000 186700 31100
rect 186600 31100 186700 31200
rect 186600 31200 186700 31300
rect 186600 31300 186700 31400
rect 186600 31400 186700 31500
rect 186600 31500 186700 31600
rect 186600 31600 186700 31700
rect 186600 31700 186700 31800
rect 186600 31800 186700 31900
rect 186600 31900 186700 32000
rect 186600 32000 186700 32100
rect 186600 32100 186700 32200
rect 186600 32200 186700 32300
rect 186600 32300 186700 32400
rect 186600 32400 186700 32500
rect 186600 32500 186700 32600
rect 186600 32600 186700 32700
rect 186600 32700 186700 32800
rect 186600 32800 186700 32900
rect 186600 32900 186700 33000
rect 186600 34700 186700 34800
rect 186600 34800 186700 34900
rect 186600 34900 186700 35000
rect 186600 35000 186700 35100
rect 186600 35100 186700 35200
rect 186600 35200 186700 35300
rect 186600 35300 186700 35400
rect 186600 35400 186700 35500
rect 186600 35500 186700 35600
rect 186600 35600 186700 35700
rect 186600 35700 186700 35800
rect 186600 35800 186700 35900
rect 186600 35900 186700 36000
rect 186600 36000 186700 36100
rect 186600 36100 186700 36200
rect 186600 36200 186700 36300
rect 186600 36300 186700 36400
rect 186600 36400 186700 36500
rect 186600 36500 186700 36600
rect 186600 36600 186700 36700
rect 186600 36700 186700 36800
rect 186600 36800 186700 36900
rect 186600 36900 186700 37000
rect 186600 37000 186700 37100
rect 186600 37100 186700 37200
rect 186600 37200 186700 37300
rect 186600 37300 186700 37400
rect 186600 37400 186700 37500
rect 186600 37500 186700 37600
rect 186600 37600 186700 37700
rect 186600 37700 186700 37800
rect 186600 37800 186700 37900
rect 186600 37900 186700 38000
rect 186600 38000 186700 38100
rect 186600 38100 186700 38200
rect 186600 38200 186700 38300
rect 186600 38300 186700 38400
rect 186600 38400 186700 38500
rect 186600 38500 186700 38600
rect 186600 38600 186700 38700
rect 186600 38700 186700 38800
rect 186700 21200 186800 21300
rect 186700 21300 186800 21400
rect 186700 21400 186800 21500
rect 186700 21500 186800 21600
rect 186700 21600 186800 21700
rect 186700 21700 186800 21800
rect 186700 21800 186800 21900
rect 186700 21900 186800 22000
rect 186700 22000 186800 22100
rect 186700 22100 186800 22200
rect 186700 22200 186800 22300
rect 186700 22300 186800 22400
rect 186700 22400 186800 22500
rect 186700 22500 186800 22600
rect 186700 22600 186800 22700
rect 186700 22700 186800 22800
rect 186700 22800 186800 22900
rect 186700 22900 186800 23000
rect 186700 23000 186800 23100
rect 186700 23100 186800 23200
rect 186700 23200 186800 23300
rect 186700 23300 186800 23400
rect 186700 23400 186800 23500
rect 186700 23500 186800 23600
rect 186700 23600 186800 23700
rect 186700 23700 186800 23800
rect 186700 23800 186800 23900
rect 186700 23900 186800 24000
rect 186700 24000 186800 24100
rect 186700 24100 186800 24200
rect 186700 24200 186800 24300
rect 186700 24300 186800 24400
rect 186700 24400 186800 24500
rect 186700 24500 186800 24600
rect 186700 24600 186800 24700
rect 186700 24700 186800 24800
rect 186700 24800 186800 24900
rect 186700 24900 186800 25000
rect 186700 25000 186800 25100
rect 186700 25100 186800 25200
rect 186700 25200 186800 25300
rect 186700 25300 186800 25400
rect 186700 25400 186800 25500
rect 186700 25500 186800 25600
rect 186700 25600 186800 25700
rect 186700 25700 186800 25800
rect 186700 25800 186800 25900
rect 186700 25900 186800 26000
rect 186700 26000 186800 26100
rect 186700 26100 186800 26200
rect 186700 26200 186800 26300
rect 186700 26300 186800 26400
rect 186700 26400 186800 26500
rect 186700 26500 186800 26600
rect 186700 26600 186800 26700
rect 186700 26700 186800 26800
rect 186700 26800 186800 26900
rect 186700 26900 186800 27000
rect 186700 27000 186800 27100
rect 186700 27100 186800 27200
rect 186700 27200 186800 27300
rect 186700 27300 186800 27400
rect 186700 27400 186800 27500
rect 186700 27500 186800 27600
rect 186700 27600 186800 27700
rect 186700 27700 186800 27800
rect 186700 27800 186800 27900
rect 186700 27900 186800 28000
rect 186700 28000 186800 28100
rect 186700 28100 186800 28200
rect 186700 28200 186800 28300
rect 186700 28300 186800 28400
rect 186700 28400 186800 28500
rect 186700 28500 186800 28600
rect 186700 28600 186800 28700
rect 186700 28700 186800 28800
rect 186700 28800 186800 28900
rect 186700 28900 186800 29000
rect 186700 29000 186800 29100
rect 186700 29100 186800 29200
rect 186700 29200 186800 29300
rect 186700 29300 186800 29400
rect 186700 29400 186800 29500
rect 186700 29500 186800 29600
rect 186700 29600 186800 29700
rect 186700 29700 186800 29800
rect 186700 29800 186800 29900
rect 186700 29900 186800 30000
rect 186700 30000 186800 30100
rect 186700 30100 186800 30200
rect 186700 30200 186800 30300
rect 186700 30300 186800 30400
rect 186700 30400 186800 30500
rect 186700 30500 186800 30600
rect 186700 30600 186800 30700
rect 186700 30700 186800 30800
rect 186700 30800 186800 30900
rect 186700 30900 186800 31000
rect 186700 31000 186800 31100
rect 186700 31100 186800 31200
rect 186700 31200 186800 31300
rect 186700 31300 186800 31400
rect 186700 31400 186800 31500
rect 186700 31500 186800 31600
rect 186700 31600 186800 31700
rect 186700 31700 186800 31800
rect 186700 31800 186800 31900
rect 186700 31900 186800 32000
rect 186700 32000 186800 32100
rect 186700 32100 186800 32200
rect 186700 32200 186800 32300
rect 186700 32300 186800 32400
rect 186700 32400 186800 32500
rect 186700 32500 186800 32600
rect 186700 32600 186800 32700
rect 186700 32700 186800 32800
rect 186700 32800 186800 32900
rect 186700 32900 186800 33000
rect 186700 33000 186800 33100
rect 186700 34600 186800 34700
rect 186700 34700 186800 34800
rect 186700 34800 186800 34900
rect 186700 34900 186800 35000
rect 186700 35000 186800 35100
rect 186700 35100 186800 35200
rect 186700 35200 186800 35300
rect 186700 35300 186800 35400
rect 186700 35400 186800 35500
rect 186700 35500 186800 35600
rect 186700 35600 186800 35700
rect 186700 35700 186800 35800
rect 186700 35800 186800 35900
rect 186700 35900 186800 36000
rect 186700 36000 186800 36100
rect 186700 36100 186800 36200
rect 186700 36200 186800 36300
rect 186700 36300 186800 36400
rect 186700 36400 186800 36500
rect 186700 36500 186800 36600
rect 186700 36600 186800 36700
rect 186700 36700 186800 36800
rect 186700 36800 186800 36900
rect 186700 36900 186800 37000
rect 186700 37000 186800 37100
rect 186700 37100 186800 37200
rect 186700 37200 186800 37300
rect 186700 37300 186800 37400
rect 186700 37400 186800 37500
rect 186700 37500 186800 37600
rect 186700 37600 186800 37700
rect 186700 37700 186800 37800
rect 186700 37800 186800 37900
rect 186700 37900 186800 38000
rect 186700 38000 186800 38100
rect 186700 38100 186800 38200
rect 186700 38200 186800 38300
rect 186700 38300 186800 38400
rect 186700 38400 186800 38500
rect 186700 38500 186800 38600
rect 186700 38600 186800 38700
rect 186700 38700 186800 38800
rect 186700 38800 186800 38900
rect 186800 21200 186900 21300
rect 186800 21300 186900 21400
rect 186800 21400 186900 21500
rect 186800 21500 186900 21600
rect 186800 21600 186900 21700
rect 186800 21700 186900 21800
rect 186800 21800 186900 21900
rect 186800 21900 186900 22000
rect 186800 22000 186900 22100
rect 186800 22100 186900 22200
rect 186800 22200 186900 22300
rect 186800 22300 186900 22400
rect 186800 22400 186900 22500
rect 186800 22500 186900 22600
rect 186800 22600 186900 22700
rect 186800 22700 186900 22800
rect 186800 22800 186900 22900
rect 186800 22900 186900 23000
rect 186800 23000 186900 23100
rect 186800 23100 186900 23200
rect 186800 23200 186900 23300
rect 186800 23300 186900 23400
rect 186800 23400 186900 23500
rect 186800 23500 186900 23600
rect 186800 23600 186900 23700
rect 186800 23700 186900 23800
rect 186800 23800 186900 23900
rect 186800 23900 186900 24000
rect 186800 24000 186900 24100
rect 186800 24100 186900 24200
rect 186800 24200 186900 24300
rect 186800 24300 186900 24400
rect 186800 24400 186900 24500
rect 186800 24500 186900 24600
rect 186800 24600 186900 24700
rect 186800 24700 186900 24800
rect 186800 24800 186900 24900
rect 186800 24900 186900 25000
rect 186800 25000 186900 25100
rect 186800 25100 186900 25200
rect 186800 25200 186900 25300
rect 186800 25300 186900 25400
rect 186800 25400 186900 25500
rect 186800 25500 186900 25600
rect 186800 25600 186900 25700
rect 186800 25700 186900 25800
rect 186800 25800 186900 25900
rect 186800 25900 186900 26000
rect 186800 26000 186900 26100
rect 186800 26100 186900 26200
rect 186800 26200 186900 26300
rect 186800 26300 186900 26400
rect 186800 26400 186900 26500
rect 186800 26500 186900 26600
rect 186800 26600 186900 26700
rect 186800 26700 186900 26800
rect 186800 26800 186900 26900
rect 186800 26900 186900 27000
rect 186800 27000 186900 27100
rect 186800 27100 186900 27200
rect 186800 27200 186900 27300
rect 186800 27300 186900 27400
rect 186800 27400 186900 27500
rect 186800 27500 186900 27600
rect 186800 27600 186900 27700
rect 186800 27700 186900 27800
rect 186800 27800 186900 27900
rect 186800 27900 186900 28000
rect 186800 28000 186900 28100
rect 186800 28100 186900 28200
rect 186800 28200 186900 28300
rect 186800 28300 186900 28400
rect 186800 28400 186900 28500
rect 186800 28500 186900 28600
rect 186800 28600 186900 28700
rect 186800 28700 186900 28800
rect 186800 28800 186900 28900
rect 186800 28900 186900 29000
rect 186800 29000 186900 29100
rect 186800 29100 186900 29200
rect 186800 29200 186900 29300
rect 186800 29300 186900 29400
rect 186800 29400 186900 29500
rect 186800 29500 186900 29600
rect 186800 29600 186900 29700
rect 186800 29700 186900 29800
rect 186800 29800 186900 29900
rect 186800 29900 186900 30000
rect 186800 30000 186900 30100
rect 186800 30100 186900 30200
rect 186800 30200 186900 30300
rect 186800 30300 186900 30400
rect 186800 30400 186900 30500
rect 186800 30500 186900 30600
rect 186800 30600 186900 30700
rect 186800 30700 186900 30800
rect 186800 30800 186900 30900
rect 186800 30900 186900 31000
rect 186800 31000 186900 31100
rect 186800 31100 186900 31200
rect 186800 31200 186900 31300
rect 186800 31300 186900 31400
rect 186800 31400 186900 31500
rect 186800 31500 186900 31600
rect 186800 31600 186900 31700
rect 186800 31700 186900 31800
rect 186800 31800 186900 31900
rect 186800 31900 186900 32000
rect 186800 32000 186900 32100
rect 186800 32100 186900 32200
rect 186800 32200 186900 32300
rect 186800 32300 186900 32400
rect 186800 32400 186900 32500
rect 186800 32500 186900 32600
rect 186800 32600 186900 32700
rect 186800 32700 186900 32800
rect 186800 32800 186900 32900
rect 186800 32900 186900 33000
rect 186800 33000 186900 33100
rect 186800 33100 186900 33200
rect 186800 34600 186900 34700
rect 186800 34700 186900 34800
rect 186800 34800 186900 34900
rect 186800 34900 186900 35000
rect 186800 35000 186900 35100
rect 186800 35100 186900 35200
rect 186800 35200 186900 35300
rect 186800 35300 186900 35400
rect 186800 35400 186900 35500
rect 186800 35500 186900 35600
rect 186800 35600 186900 35700
rect 186800 35700 186900 35800
rect 186800 35800 186900 35900
rect 186800 35900 186900 36000
rect 186800 36000 186900 36100
rect 186800 36100 186900 36200
rect 186800 36200 186900 36300
rect 186800 36300 186900 36400
rect 186800 36400 186900 36500
rect 186800 36500 186900 36600
rect 186800 36600 186900 36700
rect 186800 36700 186900 36800
rect 186800 36800 186900 36900
rect 186800 36900 186900 37000
rect 186800 37000 186900 37100
rect 186800 37100 186900 37200
rect 186800 37200 186900 37300
rect 186800 37300 186900 37400
rect 186800 37400 186900 37500
rect 186800 37500 186900 37600
rect 186800 37600 186900 37700
rect 186800 37700 186900 37800
rect 186800 37800 186900 37900
rect 186800 37900 186900 38000
rect 186800 38000 186900 38100
rect 186800 38100 186900 38200
rect 186800 38200 186900 38300
rect 186800 38300 186900 38400
rect 186800 38400 186900 38500
rect 186800 38500 186900 38600
rect 186800 38600 186900 38700
rect 186800 38700 186900 38800
rect 186800 38800 186900 38900
rect 186900 21300 187000 21400
rect 186900 21400 187000 21500
rect 186900 21500 187000 21600
rect 186900 21600 187000 21700
rect 186900 21700 187000 21800
rect 186900 21800 187000 21900
rect 186900 21900 187000 22000
rect 186900 22000 187000 22100
rect 186900 22100 187000 22200
rect 186900 22200 187000 22300
rect 186900 22300 187000 22400
rect 186900 22400 187000 22500
rect 186900 22500 187000 22600
rect 186900 22600 187000 22700
rect 186900 22700 187000 22800
rect 186900 22800 187000 22900
rect 186900 22900 187000 23000
rect 186900 23000 187000 23100
rect 186900 23100 187000 23200
rect 186900 23200 187000 23300
rect 186900 23300 187000 23400
rect 186900 23400 187000 23500
rect 186900 23500 187000 23600
rect 186900 23600 187000 23700
rect 186900 23700 187000 23800
rect 186900 23800 187000 23900
rect 186900 23900 187000 24000
rect 186900 24000 187000 24100
rect 186900 24100 187000 24200
rect 186900 24200 187000 24300
rect 186900 24300 187000 24400
rect 186900 24400 187000 24500
rect 186900 24500 187000 24600
rect 186900 24600 187000 24700
rect 186900 24700 187000 24800
rect 186900 24800 187000 24900
rect 186900 24900 187000 25000
rect 186900 25000 187000 25100
rect 186900 25100 187000 25200
rect 186900 25200 187000 25300
rect 186900 25300 187000 25400
rect 186900 25400 187000 25500
rect 186900 25500 187000 25600
rect 186900 25600 187000 25700
rect 186900 25700 187000 25800
rect 186900 25800 187000 25900
rect 186900 25900 187000 26000
rect 186900 26000 187000 26100
rect 186900 26100 187000 26200
rect 186900 26200 187000 26300
rect 186900 26300 187000 26400
rect 186900 26400 187000 26500
rect 186900 26500 187000 26600
rect 186900 26600 187000 26700
rect 186900 26700 187000 26800
rect 186900 26800 187000 26900
rect 186900 26900 187000 27000
rect 186900 27000 187000 27100
rect 186900 27100 187000 27200
rect 186900 27200 187000 27300
rect 186900 27300 187000 27400
rect 186900 27400 187000 27500
rect 186900 27500 187000 27600
rect 186900 27600 187000 27700
rect 186900 27700 187000 27800
rect 186900 27800 187000 27900
rect 186900 27900 187000 28000
rect 186900 28000 187000 28100
rect 186900 28100 187000 28200
rect 186900 28200 187000 28300
rect 186900 28300 187000 28400
rect 186900 28400 187000 28500
rect 186900 28500 187000 28600
rect 186900 28600 187000 28700
rect 186900 28700 187000 28800
rect 186900 28800 187000 28900
rect 186900 28900 187000 29000
rect 186900 29000 187000 29100
rect 186900 29100 187000 29200
rect 186900 29200 187000 29300
rect 186900 29300 187000 29400
rect 186900 29400 187000 29500
rect 186900 29500 187000 29600
rect 186900 29600 187000 29700
rect 186900 29700 187000 29800
rect 186900 29800 187000 29900
rect 186900 29900 187000 30000
rect 186900 30000 187000 30100
rect 186900 30100 187000 30200
rect 186900 30200 187000 30300
rect 186900 30300 187000 30400
rect 186900 30400 187000 30500
rect 186900 30500 187000 30600
rect 186900 30600 187000 30700
rect 186900 30700 187000 30800
rect 186900 30800 187000 30900
rect 186900 30900 187000 31000
rect 186900 31000 187000 31100
rect 186900 31100 187000 31200
rect 186900 31200 187000 31300
rect 186900 31300 187000 31400
rect 186900 31400 187000 31500
rect 186900 31500 187000 31600
rect 186900 31600 187000 31700
rect 186900 31700 187000 31800
rect 186900 31800 187000 31900
rect 186900 31900 187000 32000
rect 186900 32000 187000 32100
rect 186900 32100 187000 32200
rect 186900 32200 187000 32300
rect 186900 32300 187000 32400
rect 186900 32400 187000 32500
rect 186900 32500 187000 32600
rect 186900 32600 187000 32700
rect 186900 32700 187000 32800
rect 186900 32800 187000 32900
rect 186900 32900 187000 33000
rect 186900 33000 187000 33100
rect 186900 33100 187000 33200
rect 186900 33200 187000 33300
rect 186900 34500 187000 34600
rect 186900 34600 187000 34700
rect 186900 34700 187000 34800
rect 186900 34800 187000 34900
rect 186900 34900 187000 35000
rect 186900 35000 187000 35100
rect 186900 35100 187000 35200
rect 186900 35200 187000 35300
rect 186900 35300 187000 35400
rect 186900 35400 187000 35500
rect 186900 35500 187000 35600
rect 186900 35600 187000 35700
rect 186900 35700 187000 35800
rect 186900 35800 187000 35900
rect 186900 35900 187000 36000
rect 186900 36000 187000 36100
rect 186900 36100 187000 36200
rect 186900 36200 187000 36300
rect 186900 36300 187000 36400
rect 186900 36400 187000 36500
rect 186900 36500 187000 36600
rect 186900 36600 187000 36700
rect 186900 36700 187000 36800
rect 186900 36800 187000 36900
rect 186900 36900 187000 37000
rect 186900 37000 187000 37100
rect 186900 37100 187000 37200
rect 186900 37200 187000 37300
rect 186900 37300 187000 37400
rect 186900 37400 187000 37500
rect 186900 37500 187000 37600
rect 186900 37600 187000 37700
rect 186900 37700 187000 37800
rect 186900 37800 187000 37900
rect 186900 37900 187000 38000
rect 186900 38000 187000 38100
rect 186900 38100 187000 38200
rect 186900 38200 187000 38300
rect 186900 38300 187000 38400
rect 186900 38400 187000 38500
rect 186900 38500 187000 38600
rect 186900 38600 187000 38700
rect 186900 38700 187000 38800
rect 186900 38800 187000 38900
rect 186900 38900 187000 39000
rect 187000 21300 187100 21400
rect 187000 21400 187100 21500
rect 187000 21500 187100 21600
rect 187000 21600 187100 21700
rect 187000 21700 187100 21800
rect 187000 21800 187100 21900
rect 187000 21900 187100 22000
rect 187000 22000 187100 22100
rect 187000 22100 187100 22200
rect 187000 22200 187100 22300
rect 187000 22300 187100 22400
rect 187000 22400 187100 22500
rect 187000 22500 187100 22600
rect 187000 22600 187100 22700
rect 187000 22700 187100 22800
rect 187000 22800 187100 22900
rect 187000 22900 187100 23000
rect 187000 23000 187100 23100
rect 187000 23100 187100 23200
rect 187000 23200 187100 23300
rect 187000 23300 187100 23400
rect 187000 23400 187100 23500
rect 187000 23500 187100 23600
rect 187000 23600 187100 23700
rect 187000 23700 187100 23800
rect 187000 23800 187100 23900
rect 187000 23900 187100 24000
rect 187000 24000 187100 24100
rect 187000 24100 187100 24200
rect 187000 24200 187100 24300
rect 187000 24300 187100 24400
rect 187000 24400 187100 24500
rect 187000 24500 187100 24600
rect 187000 24600 187100 24700
rect 187000 24700 187100 24800
rect 187000 24800 187100 24900
rect 187000 24900 187100 25000
rect 187000 25000 187100 25100
rect 187000 25100 187100 25200
rect 187000 25200 187100 25300
rect 187000 25300 187100 25400
rect 187000 25400 187100 25500
rect 187000 25500 187100 25600
rect 187000 25600 187100 25700
rect 187000 25700 187100 25800
rect 187000 25800 187100 25900
rect 187000 25900 187100 26000
rect 187000 26000 187100 26100
rect 187000 26100 187100 26200
rect 187000 26200 187100 26300
rect 187000 26300 187100 26400
rect 187000 26400 187100 26500
rect 187000 26500 187100 26600
rect 187000 26600 187100 26700
rect 187000 26700 187100 26800
rect 187000 26800 187100 26900
rect 187000 26900 187100 27000
rect 187000 27000 187100 27100
rect 187000 27100 187100 27200
rect 187000 27200 187100 27300
rect 187000 27300 187100 27400
rect 187000 27400 187100 27500
rect 187000 27500 187100 27600
rect 187000 27600 187100 27700
rect 187000 27700 187100 27800
rect 187000 27800 187100 27900
rect 187000 27900 187100 28000
rect 187000 28000 187100 28100
rect 187000 28100 187100 28200
rect 187000 28200 187100 28300
rect 187000 28300 187100 28400
rect 187000 28400 187100 28500
rect 187000 28500 187100 28600
rect 187000 28600 187100 28700
rect 187000 28700 187100 28800
rect 187000 28800 187100 28900
rect 187000 28900 187100 29000
rect 187000 29000 187100 29100
rect 187000 29100 187100 29200
rect 187000 29200 187100 29300
rect 187000 29300 187100 29400
rect 187000 29400 187100 29500
rect 187000 29500 187100 29600
rect 187000 29600 187100 29700
rect 187000 29700 187100 29800
rect 187000 29800 187100 29900
rect 187000 29900 187100 30000
rect 187000 30000 187100 30100
rect 187000 30100 187100 30200
rect 187000 30200 187100 30300
rect 187000 30300 187100 30400
rect 187000 30400 187100 30500
rect 187000 30500 187100 30600
rect 187000 30600 187100 30700
rect 187000 30700 187100 30800
rect 187000 30800 187100 30900
rect 187000 30900 187100 31000
rect 187000 31000 187100 31100
rect 187000 31100 187100 31200
rect 187000 31200 187100 31300
rect 187000 31300 187100 31400
rect 187000 31400 187100 31500
rect 187000 31500 187100 31600
rect 187000 31600 187100 31700
rect 187000 31700 187100 31800
rect 187000 31800 187100 31900
rect 187000 31900 187100 32000
rect 187000 32000 187100 32100
rect 187000 32100 187100 32200
rect 187000 32200 187100 32300
rect 187000 32300 187100 32400
rect 187000 32400 187100 32500
rect 187000 32500 187100 32600
rect 187000 32600 187100 32700
rect 187000 32700 187100 32800
rect 187000 32800 187100 32900
rect 187000 32900 187100 33000
rect 187000 33000 187100 33100
rect 187000 33100 187100 33200
rect 187000 33200 187100 33300
rect 187000 33300 187100 33400
rect 187000 34500 187100 34600
rect 187000 34600 187100 34700
rect 187000 34700 187100 34800
rect 187000 34800 187100 34900
rect 187000 34900 187100 35000
rect 187000 35000 187100 35100
rect 187000 35100 187100 35200
rect 187000 35200 187100 35300
rect 187000 35300 187100 35400
rect 187000 35400 187100 35500
rect 187000 35500 187100 35600
rect 187000 35600 187100 35700
rect 187000 35700 187100 35800
rect 187000 35800 187100 35900
rect 187000 35900 187100 36000
rect 187000 36000 187100 36100
rect 187000 36100 187100 36200
rect 187000 36200 187100 36300
rect 187000 36300 187100 36400
rect 187000 36400 187100 36500
rect 187000 36500 187100 36600
rect 187000 36600 187100 36700
rect 187000 36700 187100 36800
rect 187000 36800 187100 36900
rect 187000 36900 187100 37000
rect 187000 37000 187100 37100
rect 187000 37100 187100 37200
rect 187000 37200 187100 37300
rect 187000 37300 187100 37400
rect 187000 37400 187100 37500
rect 187000 37500 187100 37600
rect 187000 37600 187100 37700
rect 187000 37700 187100 37800
rect 187000 37800 187100 37900
rect 187000 37900 187100 38000
rect 187000 38000 187100 38100
rect 187000 38100 187100 38200
rect 187000 38200 187100 38300
rect 187000 38300 187100 38400
rect 187000 38400 187100 38500
rect 187000 38500 187100 38600
rect 187000 38600 187100 38700
rect 187000 38700 187100 38800
rect 187000 38800 187100 38900
rect 187000 38900 187100 39000
rect 187100 21400 187200 21500
rect 187100 21500 187200 21600
rect 187100 21600 187200 21700
rect 187100 21700 187200 21800
rect 187100 21800 187200 21900
rect 187100 21900 187200 22000
rect 187100 22000 187200 22100
rect 187100 22100 187200 22200
rect 187100 22200 187200 22300
rect 187100 22300 187200 22400
rect 187100 22400 187200 22500
rect 187100 22500 187200 22600
rect 187100 22600 187200 22700
rect 187100 22700 187200 22800
rect 187100 22800 187200 22900
rect 187100 22900 187200 23000
rect 187100 23000 187200 23100
rect 187100 23100 187200 23200
rect 187100 23200 187200 23300
rect 187100 23300 187200 23400
rect 187100 23400 187200 23500
rect 187100 23500 187200 23600
rect 187100 23600 187200 23700
rect 187100 23700 187200 23800
rect 187100 23800 187200 23900
rect 187100 23900 187200 24000
rect 187100 24000 187200 24100
rect 187100 24100 187200 24200
rect 187100 24200 187200 24300
rect 187100 24300 187200 24400
rect 187100 24400 187200 24500
rect 187100 24500 187200 24600
rect 187100 24600 187200 24700
rect 187100 24700 187200 24800
rect 187100 24800 187200 24900
rect 187100 24900 187200 25000
rect 187100 25000 187200 25100
rect 187100 25100 187200 25200
rect 187100 25200 187200 25300
rect 187100 25300 187200 25400
rect 187100 25400 187200 25500
rect 187100 25500 187200 25600
rect 187100 25600 187200 25700
rect 187100 25700 187200 25800
rect 187100 25800 187200 25900
rect 187100 25900 187200 26000
rect 187100 26000 187200 26100
rect 187100 26100 187200 26200
rect 187100 26200 187200 26300
rect 187100 26300 187200 26400
rect 187100 26400 187200 26500
rect 187100 26500 187200 26600
rect 187100 26600 187200 26700
rect 187100 26700 187200 26800
rect 187100 26800 187200 26900
rect 187100 26900 187200 27000
rect 187100 27000 187200 27100
rect 187100 27100 187200 27200
rect 187100 27200 187200 27300
rect 187100 27300 187200 27400
rect 187100 27400 187200 27500
rect 187100 27500 187200 27600
rect 187100 27600 187200 27700
rect 187100 27700 187200 27800
rect 187100 27800 187200 27900
rect 187100 27900 187200 28000
rect 187100 28000 187200 28100
rect 187100 28100 187200 28200
rect 187100 28200 187200 28300
rect 187100 28300 187200 28400
rect 187100 28400 187200 28500
rect 187100 28500 187200 28600
rect 187100 28600 187200 28700
rect 187100 28700 187200 28800
rect 187100 28800 187200 28900
rect 187100 28900 187200 29000
rect 187100 29000 187200 29100
rect 187100 29100 187200 29200
rect 187100 29200 187200 29300
rect 187100 29300 187200 29400
rect 187100 29400 187200 29500
rect 187100 29500 187200 29600
rect 187100 29600 187200 29700
rect 187100 29700 187200 29800
rect 187100 29800 187200 29900
rect 187100 29900 187200 30000
rect 187100 30000 187200 30100
rect 187100 30100 187200 30200
rect 187100 30200 187200 30300
rect 187100 30300 187200 30400
rect 187100 30400 187200 30500
rect 187100 30500 187200 30600
rect 187100 30600 187200 30700
rect 187100 30700 187200 30800
rect 187100 30800 187200 30900
rect 187100 30900 187200 31000
rect 187100 31000 187200 31100
rect 187100 31100 187200 31200
rect 187100 31200 187200 31300
rect 187100 31300 187200 31400
rect 187100 31400 187200 31500
rect 187100 31500 187200 31600
rect 187100 31600 187200 31700
rect 187100 31700 187200 31800
rect 187100 31800 187200 31900
rect 187100 31900 187200 32000
rect 187100 32000 187200 32100
rect 187100 32100 187200 32200
rect 187100 32200 187200 32300
rect 187100 32300 187200 32400
rect 187100 32400 187200 32500
rect 187100 32500 187200 32600
rect 187100 32600 187200 32700
rect 187100 32700 187200 32800
rect 187100 32800 187200 32900
rect 187100 32900 187200 33000
rect 187100 33000 187200 33100
rect 187100 33100 187200 33200
rect 187100 33200 187200 33300
rect 187100 33300 187200 33400
rect 187100 34400 187200 34500
rect 187100 34500 187200 34600
rect 187100 34600 187200 34700
rect 187100 34700 187200 34800
rect 187100 34800 187200 34900
rect 187100 34900 187200 35000
rect 187100 35000 187200 35100
rect 187100 35100 187200 35200
rect 187100 35200 187200 35300
rect 187100 35300 187200 35400
rect 187100 35400 187200 35500
rect 187100 35500 187200 35600
rect 187100 35600 187200 35700
rect 187100 35700 187200 35800
rect 187100 35800 187200 35900
rect 187100 35900 187200 36000
rect 187100 36000 187200 36100
rect 187100 36100 187200 36200
rect 187100 36200 187200 36300
rect 187100 36300 187200 36400
rect 187100 36400 187200 36500
rect 187100 36800 187200 36900
rect 187100 36900 187200 37000
rect 187100 37000 187200 37100
rect 187100 37100 187200 37200
rect 187100 37200 187200 37300
rect 187100 37300 187200 37400
rect 187100 37400 187200 37500
rect 187100 37500 187200 37600
rect 187100 37600 187200 37700
rect 187100 37700 187200 37800
rect 187100 37800 187200 37900
rect 187100 37900 187200 38000
rect 187100 38000 187200 38100
rect 187100 38100 187200 38200
rect 187100 38200 187200 38300
rect 187100 38300 187200 38400
rect 187100 38400 187200 38500
rect 187100 38500 187200 38600
rect 187100 38600 187200 38700
rect 187100 38700 187200 38800
rect 187100 38800 187200 38900
rect 187100 38900 187200 39000
rect 187200 21500 187300 21600
rect 187200 21600 187300 21700
rect 187200 21700 187300 21800
rect 187200 21800 187300 21900
rect 187200 21900 187300 22000
rect 187200 22000 187300 22100
rect 187200 22100 187300 22200
rect 187200 22200 187300 22300
rect 187200 22300 187300 22400
rect 187200 22400 187300 22500
rect 187200 22500 187300 22600
rect 187200 22600 187300 22700
rect 187200 22700 187300 22800
rect 187200 22800 187300 22900
rect 187200 22900 187300 23000
rect 187200 23000 187300 23100
rect 187200 23100 187300 23200
rect 187200 23200 187300 23300
rect 187200 23300 187300 23400
rect 187200 23400 187300 23500
rect 187200 23500 187300 23600
rect 187200 23600 187300 23700
rect 187200 23700 187300 23800
rect 187200 23800 187300 23900
rect 187200 23900 187300 24000
rect 187200 24000 187300 24100
rect 187200 24100 187300 24200
rect 187200 24200 187300 24300
rect 187200 24300 187300 24400
rect 187200 24400 187300 24500
rect 187200 24500 187300 24600
rect 187200 24600 187300 24700
rect 187200 24700 187300 24800
rect 187200 24800 187300 24900
rect 187200 24900 187300 25000
rect 187200 25000 187300 25100
rect 187200 25100 187300 25200
rect 187200 25200 187300 25300
rect 187200 25300 187300 25400
rect 187200 25400 187300 25500
rect 187200 25500 187300 25600
rect 187200 25600 187300 25700
rect 187200 25700 187300 25800
rect 187200 25800 187300 25900
rect 187200 25900 187300 26000
rect 187200 26000 187300 26100
rect 187200 26100 187300 26200
rect 187200 26200 187300 26300
rect 187200 26300 187300 26400
rect 187200 26400 187300 26500
rect 187200 26500 187300 26600
rect 187200 26600 187300 26700
rect 187200 26700 187300 26800
rect 187200 26800 187300 26900
rect 187200 26900 187300 27000
rect 187200 27000 187300 27100
rect 187200 27100 187300 27200
rect 187200 27200 187300 27300
rect 187200 27300 187300 27400
rect 187200 27400 187300 27500
rect 187200 27500 187300 27600
rect 187200 27600 187300 27700
rect 187200 27700 187300 27800
rect 187200 27800 187300 27900
rect 187200 27900 187300 28000
rect 187200 28000 187300 28100
rect 187200 28100 187300 28200
rect 187200 28200 187300 28300
rect 187200 28300 187300 28400
rect 187200 28400 187300 28500
rect 187200 28500 187300 28600
rect 187200 28600 187300 28700
rect 187200 28700 187300 28800
rect 187200 28800 187300 28900
rect 187200 28900 187300 29000
rect 187200 29000 187300 29100
rect 187200 29100 187300 29200
rect 187200 29200 187300 29300
rect 187200 29300 187300 29400
rect 187200 29400 187300 29500
rect 187200 29500 187300 29600
rect 187200 29600 187300 29700
rect 187200 29700 187300 29800
rect 187200 29800 187300 29900
rect 187200 29900 187300 30000
rect 187200 30000 187300 30100
rect 187200 30100 187300 30200
rect 187200 30200 187300 30300
rect 187200 30300 187300 30400
rect 187200 30400 187300 30500
rect 187200 30500 187300 30600
rect 187200 30600 187300 30700
rect 187200 30700 187300 30800
rect 187200 30800 187300 30900
rect 187200 30900 187300 31000
rect 187200 31000 187300 31100
rect 187200 31100 187300 31200
rect 187200 31200 187300 31300
rect 187200 31300 187300 31400
rect 187200 31400 187300 31500
rect 187200 31500 187300 31600
rect 187200 31600 187300 31700
rect 187200 31700 187300 31800
rect 187200 31800 187300 31900
rect 187200 31900 187300 32000
rect 187200 32000 187300 32100
rect 187200 32100 187300 32200
rect 187200 32200 187300 32300
rect 187200 32300 187300 32400
rect 187200 32400 187300 32500
rect 187200 32500 187300 32600
rect 187200 32600 187300 32700
rect 187200 32700 187300 32800
rect 187200 32800 187300 32900
rect 187200 32900 187300 33000
rect 187200 33000 187300 33100
rect 187200 33100 187300 33200
rect 187200 33200 187300 33300
rect 187200 33300 187300 33400
rect 187200 33400 187300 33500
rect 187200 34400 187300 34500
rect 187200 34500 187300 34600
rect 187200 34600 187300 34700
rect 187200 34700 187300 34800
rect 187200 34800 187300 34900
rect 187200 34900 187300 35000
rect 187200 35000 187300 35100
rect 187200 35100 187300 35200
rect 187200 35200 187300 35300
rect 187200 35300 187300 35400
rect 187200 35400 187300 35500
rect 187200 35500 187300 35600
rect 187200 35600 187300 35700
rect 187200 35700 187300 35800
rect 187200 35800 187300 35900
rect 187200 35900 187300 36000
rect 187200 36000 187300 36100
rect 187200 36100 187300 36200
rect 187200 37100 187300 37200
rect 187200 37200 187300 37300
rect 187200 37300 187300 37400
rect 187200 37400 187300 37500
rect 187200 37500 187300 37600
rect 187200 37600 187300 37700
rect 187200 37700 187300 37800
rect 187200 37800 187300 37900
rect 187200 37900 187300 38000
rect 187200 38000 187300 38100
rect 187200 38100 187300 38200
rect 187200 38200 187300 38300
rect 187200 38300 187300 38400
rect 187200 38400 187300 38500
rect 187200 38500 187300 38600
rect 187200 38600 187300 38700
rect 187200 38700 187300 38800
rect 187200 38800 187300 38900
rect 187200 38900 187300 39000
rect 187200 39000 187300 39100
rect 187300 21600 187400 21700
rect 187300 21700 187400 21800
rect 187300 21800 187400 21900
rect 187300 21900 187400 22000
rect 187300 22000 187400 22100
rect 187300 22100 187400 22200
rect 187300 22200 187400 22300
rect 187300 22300 187400 22400
rect 187300 22400 187400 22500
rect 187300 22500 187400 22600
rect 187300 22600 187400 22700
rect 187300 22700 187400 22800
rect 187300 22800 187400 22900
rect 187300 22900 187400 23000
rect 187300 23000 187400 23100
rect 187300 23100 187400 23200
rect 187300 23200 187400 23300
rect 187300 23300 187400 23400
rect 187300 23400 187400 23500
rect 187300 23500 187400 23600
rect 187300 23600 187400 23700
rect 187300 23700 187400 23800
rect 187300 23800 187400 23900
rect 187300 23900 187400 24000
rect 187300 24000 187400 24100
rect 187300 24100 187400 24200
rect 187300 24200 187400 24300
rect 187300 24300 187400 24400
rect 187300 24400 187400 24500
rect 187300 24500 187400 24600
rect 187300 24600 187400 24700
rect 187300 24700 187400 24800
rect 187300 24800 187400 24900
rect 187300 24900 187400 25000
rect 187300 25000 187400 25100
rect 187300 25100 187400 25200
rect 187300 25200 187400 25300
rect 187300 25300 187400 25400
rect 187300 25400 187400 25500
rect 187300 25500 187400 25600
rect 187300 25600 187400 25700
rect 187300 25700 187400 25800
rect 187300 25800 187400 25900
rect 187300 25900 187400 26000
rect 187300 26000 187400 26100
rect 187300 26100 187400 26200
rect 187300 26200 187400 26300
rect 187300 26300 187400 26400
rect 187300 26400 187400 26500
rect 187300 26500 187400 26600
rect 187300 26600 187400 26700
rect 187300 26700 187400 26800
rect 187300 26800 187400 26900
rect 187300 26900 187400 27000
rect 187300 27000 187400 27100
rect 187300 27100 187400 27200
rect 187300 27200 187400 27300
rect 187300 27300 187400 27400
rect 187300 27400 187400 27500
rect 187300 27500 187400 27600
rect 187300 27600 187400 27700
rect 187300 27700 187400 27800
rect 187300 27800 187400 27900
rect 187300 27900 187400 28000
rect 187300 28000 187400 28100
rect 187300 28100 187400 28200
rect 187300 28200 187400 28300
rect 187300 28300 187400 28400
rect 187300 28400 187400 28500
rect 187300 28500 187400 28600
rect 187300 28600 187400 28700
rect 187300 28700 187400 28800
rect 187300 28800 187400 28900
rect 187300 28900 187400 29000
rect 187300 29000 187400 29100
rect 187300 29100 187400 29200
rect 187300 29200 187400 29300
rect 187300 29300 187400 29400
rect 187300 29400 187400 29500
rect 187300 29500 187400 29600
rect 187300 29600 187400 29700
rect 187300 29700 187400 29800
rect 187300 29800 187400 29900
rect 187300 29900 187400 30000
rect 187300 30000 187400 30100
rect 187300 30100 187400 30200
rect 187300 30200 187400 30300
rect 187300 30300 187400 30400
rect 187300 30400 187400 30500
rect 187300 30500 187400 30600
rect 187300 30600 187400 30700
rect 187300 30700 187400 30800
rect 187300 30800 187400 30900
rect 187300 30900 187400 31000
rect 187300 31000 187400 31100
rect 187300 31100 187400 31200
rect 187300 31200 187400 31300
rect 187300 31300 187400 31400
rect 187300 31400 187400 31500
rect 187300 31500 187400 31600
rect 187300 31600 187400 31700
rect 187300 31700 187400 31800
rect 187300 31800 187400 31900
rect 187300 31900 187400 32000
rect 187300 32000 187400 32100
rect 187300 32100 187400 32200
rect 187300 32200 187400 32300
rect 187300 32300 187400 32400
rect 187300 32400 187400 32500
rect 187300 32500 187400 32600
rect 187300 32600 187400 32700
rect 187300 32700 187400 32800
rect 187300 32800 187400 32900
rect 187300 32900 187400 33000
rect 187300 33000 187400 33100
rect 187300 33100 187400 33200
rect 187300 33200 187400 33300
rect 187300 33300 187400 33400
rect 187300 33400 187400 33500
rect 187300 34400 187400 34500
rect 187300 34500 187400 34600
rect 187300 34600 187400 34700
rect 187300 34700 187400 34800
rect 187300 34800 187400 34900
rect 187300 34900 187400 35000
rect 187300 35000 187400 35100
rect 187300 35100 187400 35200
rect 187300 35200 187400 35300
rect 187300 35300 187400 35400
rect 187300 35400 187400 35500
rect 187300 35500 187400 35600
rect 187300 35600 187400 35700
rect 187300 35700 187400 35800
rect 187300 35800 187400 35900
rect 187300 35900 187400 36000
rect 187300 36000 187400 36100
rect 187300 37200 187400 37300
rect 187300 37300 187400 37400
rect 187300 37400 187400 37500
rect 187300 37500 187400 37600
rect 187300 37600 187400 37700
rect 187300 37700 187400 37800
rect 187300 37800 187400 37900
rect 187300 37900 187400 38000
rect 187300 38000 187400 38100
rect 187300 38100 187400 38200
rect 187300 38200 187400 38300
rect 187300 38300 187400 38400
rect 187300 38400 187400 38500
rect 187300 38500 187400 38600
rect 187300 38600 187400 38700
rect 187300 38700 187400 38800
rect 187300 38800 187400 38900
rect 187300 38900 187400 39000
rect 187300 39000 187400 39100
rect 187400 21700 187500 21800
rect 187400 21800 187500 21900
rect 187400 21900 187500 22000
rect 187400 22000 187500 22100
rect 187400 22100 187500 22200
rect 187400 22200 187500 22300
rect 187400 22300 187500 22400
rect 187400 22400 187500 22500
rect 187400 22500 187500 22600
rect 187400 22600 187500 22700
rect 187400 22700 187500 22800
rect 187400 22800 187500 22900
rect 187400 22900 187500 23000
rect 187400 23000 187500 23100
rect 187400 23100 187500 23200
rect 187400 23200 187500 23300
rect 187400 23300 187500 23400
rect 187400 23400 187500 23500
rect 187400 23500 187500 23600
rect 187400 23600 187500 23700
rect 187400 23700 187500 23800
rect 187400 23800 187500 23900
rect 187400 23900 187500 24000
rect 187400 24000 187500 24100
rect 187400 24100 187500 24200
rect 187400 24200 187500 24300
rect 187400 24300 187500 24400
rect 187400 24400 187500 24500
rect 187400 24500 187500 24600
rect 187400 24600 187500 24700
rect 187400 24700 187500 24800
rect 187400 24800 187500 24900
rect 187400 24900 187500 25000
rect 187400 25000 187500 25100
rect 187400 25100 187500 25200
rect 187400 25200 187500 25300
rect 187400 25300 187500 25400
rect 187400 25400 187500 25500
rect 187400 25500 187500 25600
rect 187400 25600 187500 25700
rect 187400 25700 187500 25800
rect 187400 25800 187500 25900
rect 187400 25900 187500 26000
rect 187400 26000 187500 26100
rect 187400 26100 187500 26200
rect 187400 26200 187500 26300
rect 187400 26300 187500 26400
rect 187400 26400 187500 26500
rect 187400 26500 187500 26600
rect 187400 26600 187500 26700
rect 187400 26700 187500 26800
rect 187400 26800 187500 26900
rect 187400 26900 187500 27000
rect 187400 27000 187500 27100
rect 187400 27100 187500 27200
rect 187400 27200 187500 27300
rect 187400 27300 187500 27400
rect 187400 27400 187500 27500
rect 187400 27500 187500 27600
rect 187400 27600 187500 27700
rect 187400 27700 187500 27800
rect 187400 27800 187500 27900
rect 187400 27900 187500 28000
rect 187400 28000 187500 28100
rect 187400 28100 187500 28200
rect 187400 28200 187500 28300
rect 187400 28300 187500 28400
rect 187400 28400 187500 28500
rect 187400 28500 187500 28600
rect 187400 28600 187500 28700
rect 187400 28700 187500 28800
rect 187400 28800 187500 28900
rect 187400 28900 187500 29000
rect 187400 29000 187500 29100
rect 187400 29100 187500 29200
rect 187400 29200 187500 29300
rect 187400 29300 187500 29400
rect 187400 29400 187500 29500
rect 187400 29500 187500 29600
rect 187400 29600 187500 29700
rect 187400 29700 187500 29800
rect 187400 29800 187500 29900
rect 187400 29900 187500 30000
rect 187400 30000 187500 30100
rect 187400 30100 187500 30200
rect 187400 30200 187500 30300
rect 187400 30300 187500 30400
rect 187400 30400 187500 30500
rect 187400 30500 187500 30600
rect 187400 30600 187500 30700
rect 187400 30700 187500 30800
rect 187400 30800 187500 30900
rect 187400 30900 187500 31000
rect 187400 31000 187500 31100
rect 187400 31100 187500 31200
rect 187400 31200 187500 31300
rect 187400 31300 187500 31400
rect 187400 31400 187500 31500
rect 187400 31500 187500 31600
rect 187400 31600 187500 31700
rect 187400 31700 187500 31800
rect 187400 31800 187500 31900
rect 187400 31900 187500 32000
rect 187400 32000 187500 32100
rect 187400 32100 187500 32200
rect 187400 32200 187500 32300
rect 187400 32300 187500 32400
rect 187400 32400 187500 32500
rect 187400 32500 187500 32600
rect 187400 32600 187500 32700
rect 187400 32700 187500 32800
rect 187400 32800 187500 32900
rect 187400 32900 187500 33000
rect 187400 33000 187500 33100
rect 187400 33100 187500 33200
rect 187400 33200 187500 33300
rect 187400 33300 187500 33400
rect 187400 33400 187500 33500
rect 187400 33500 187500 33600
rect 187400 34300 187500 34400
rect 187400 34400 187500 34500
rect 187400 34500 187500 34600
rect 187400 34600 187500 34700
rect 187400 34700 187500 34800
rect 187400 34800 187500 34900
rect 187400 34900 187500 35000
rect 187400 35000 187500 35100
rect 187400 35100 187500 35200
rect 187400 35200 187500 35300
rect 187400 35300 187500 35400
rect 187400 35400 187500 35500
rect 187400 35500 187500 35600
rect 187400 35600 187500 35700
rect 187400 35700 187500 35800
rect 187400 35800 187500 35900
rect 187400 35900 187500 36000
rect 187400 37300 187500 37400
rect 187400 37400 187500 37500
rect 187400 37500 187500 37600
rect 187400 37600 187500 37700
rect 187400 37700 187500 37800
rect 187400 37800 187500 37900
rect 187400 37900 187500 38000
rect 187400 38000 187500 38100
rect 187400 38100 187500 38200
rect 187400 38200 187500 38300
rect 187400 38300 187500 38400
rect 187400 38400 187500 38500
rect 187400 38500 187500 38600
rect 187400 38600 187500 38700
rect 187400 38700 187500 38800
rect 187400 38800 187500 38900
rect 187400 38900 187500 39000
rect 187400 39000 187500 39100
rect 187500 21800 187600 21900
rect 187500 21900 187600 22000
rect 187500 22000 187600 22100
rect 187500 22100 187600 22200
rect 187500 22200 187600 22300
rect 187500 22300 187600 22400
rect 187500 22400 187600 22500
rect 187500 22500 187600 22600
rect 187500 22600 187600 22700
rect 187500 22700 187600 22800
rect 187500 22800 187600 22900
rect 187500 22900 187600 23000
rect 187500 23000 187600 23100
rect 187500 23100 187600 23200
rect 187500 23200 187600 23300
rect 187500 23300 187600 23400
rect 187500 23400 187600 23500
rect 187500 23500 187600 23600
rect 187500 23600 187600 23700
rect 187500 23700 187600 23800
rect 187500 23800 187600 23900
rect 187500 23900 187600 24000
rect 187500 24000 187600 24100
rect 187500 24100 187600 24200
rect 187500 24200 187600 24300
rect 187500 24300 187600 24400
rect 187500 24400 187600 24500
rect 187500 24500 187600 24600
rect 187500 24600 187600 24700
rect 187500 24700 187600 24800
rect 187500 24800 187600 24900
rect 187500 24900 187600 25000
rect 187500 25000 187600 25100
rect 187500 25100 187600 25200
rect 187500 25200 187600 25300
rect 187500 25300 187600 25400
rect 187500 25400 187600 25500
rect 187500 25500 187600 25600
rect 187500 25600 187600 25700
rect 187500 25700 187600 25800
rect 187500 25800 187600 25900
rect 187500 25900 187600 26000
rect 187500 26000 187600 26100
rect 187500 26100 187600 26200
rect 187500 26200 187600 26300
rect 187500 26300 187600 26400
rect 187500 26400 187600 26500
rect 187500 26500 187600 26600
rect 187500 26600 187600 26700
rect 187500 26700 187600 26800
rect 187500 26800 187600 26900
rect 187500 26900 187600 27000
rect 187500 27000 187600 27100
rect 187500 27100 187600 27200
rect 187500 27200 187600 27300
rect 187500 27300 187600 27400
rect 187500 27400 187600 27500
rect 187500 27500 187600 27600
rect 187500 27600 187600 27700
rect 187500 27700 187600 27800
rect 187500 27800 187600 27900
rect 187500 27900 187600 28000
rect 187500 28000 187600 28100
rect 187500 28100 187600 28200
rect 187500 28200 187600 28300
rect 187500 28300 187600 28400
rect 187500 28400 187600 28500
rect 187500 28500 187600 28600
rect 187500 28600 187600 28700
rect 187500 28700 187600 28800
rect 187500 28800 187600 28900
rect 187500 28900 187600 29000
rect 187500 29000 187600 29100
rect 187500 29100 187600 29200
rect 187500 29200 187600 29300
rect 187500 29300 187600 29400
rect 187500 29400 187600 29500
rect 187500 29500 187600 29600
rect 187500 29600 187600 29700
rect 187500 29700 187600 29800
rect 187500 29800 187600 29900
rect 187500 29900 187600 30000
rect 187500 30000 187600 30100
rect 187500 30100 187600 30200
rect 187500 30200 187600 30300
rect 187500 30300 187600 30400
rect 187500 30400 187600 30500
rect 187500 30500 187600 30600
rect 187500 30600 187600 30700
rect 187500 30700 187600 30800
rect 187500 30800 187600 30900
rect 187500 30900 187600 31000
rect 187500 31000 187600 31100
rect 187500 31100 187600 31200
rect 187500 31200 187600 31300
rect 187500 31300 187600 31400
rect 187500 31400 187600 31500
rect 187500 31500 187600 31600
rect 187500 31600 187600 31700
rect 187500 31700 187600 31800
rect 187500 31800 187600 31900
rect 187500 31900 187600 32000
rect 187500 32000 187600 32100
rect 187500 32100 187600 32200
rect 187500 32200 187600 32300
rect 187500 32300 187600 32400
rect 187500 32400 187600 32500
rect 187500 32500 187600 32600
rect 187500 32600 187600 32700
rect 187500 32700 187600 32800
rect 187500 32800 187600 32900
rect 187500 32900 187600 33000
rect 187500 33000 187600 33100
rect 187500 33100 187600 33200
rect 187500 33200 187600 33300
rect 187500 33300 187600 33400
rect 187500 33400 187600 33500
rect 187500 33500 187600 33600
rect 187500 34300 187600 34400
rect 187500 34400 187600 34500
rect 187500 34500 187600 34600
rect 187500 34600 187600 34700
rect 187500 34700 187600 34800
rect 187500 34800 187600 34900
rect 187500 34900 187600 35000
rect 187500 35000 187600 35100
rect 187500 35100 187600 35200
rect 187500 35200 187600 35300
rect 187500 35300 187600 35400
rect 187500 35400 187600 35500
rect 187500 35500 187600 35600
rect 187500 35600 187600 35700
rect 187500 35700 187600 35800
rect 187500 35800 187600 35900
rect 187500 37400 187600 37500
rect 187500 37500 187600 37600
rect 187500 37600 187600 37700
rect 187500 37700 187600 37800
rect 187500 37800 187600 37900
rect 187500 37900 187600 38000
rect 187500 38000 187600 38100
rect 187500 38100 187600 38200
rect 187500 38200 187600 38300
rect 187500 38300 187600 38400
rect 187500 38400 187600 38500
rect 187500 38500 187600 38600
rect 187500 38600 187600 38700
rect 187500 38700 187600 38800
rect 187500 38800 187600 38900
rect 187500 38900 187600 39000
rect 187500 39000 187600 39100
rect 187600 22000 187700 22100
rect 187600 22100 187700 22200
rect 187600 22200 187700 22300
rect 187600 22300 187700 22400
rect 187600 22400 187700 22500
rect 187600 22500 187700 22600
rect 187600 22600 187700 22700
rect 187600 22700 187700 22800
rect 187600 22800 187700 22900
rect 187600 22900 187700 23000
rect 187600 23000 187700 23100
rect 187600 23100 187700 23200
rect 187600 23200 187700 23300
rect 187600 23300 187700 23400
rect 187600 23500 187700 23600
rect 187600 28000 187700 28100
rect 187600 28200 187700 28300
rect 187600 28300 187700 28400
rect 187600 28400 187700 28500
rect 187600 28500 187700 28600
rect 187600 28600 187700 28700
rect 187600 28700 187700 28800
rect 187600 28800 187700 28900
rect 187600 28900 187700 29000
rect 187600 29000 187700 29100
rect 187600 29100 187700 29200
rect 187600 29200 187700 29300
rect 187600 29300 187700 29400
rect 187600 29400 187700 29500
rect 187600 29500 187700 29600
rect 187600 29600 187700 29700
rect 187600 29700 187700 29800
rect 187600 29800 187700 29900
rect 187600 29900 187700 30000
rect 187600 30000 187700 30100
rect 187600 30100 187700 30200
rect 187600 30200 187700 30300
rect 187600 30300 187700 30400
rect 187600 30400 187700 30500
rect 187600 30500 187700 30600
rect 187600 30600 187700 30700
rect 187600 30700 187700 30800
rect 187600 30800 187700 30900
rect 187600 30900 187700 31000
rect 187600 31000 187700 31100
rect 187600 31100 187700 31200
rect 187600 31200 187700 31300
rect 187600 31300 187700 31400
rect 187600 31400 187700 31500
rect 187600 31500 187700 31600
rect 187600 31600 187700 31700
rect 187600 31700 187700 31800
rect 187600 31800 187700 31900
rect 187600 31900 187700 32000
rect 187600 32000 187700 32100
rect 187600 32100 187700 32200
rect 187600 32200 187700 32300
rect 187600 32300 187700 32400
rect 187600 32400 187700 32500
rect 187600 32500 187700 32600
rect 187600 32600 187700 32700
rect 187600 32700 187700 32800
rect 187600 32800 187700 32900
rect 187600 32900 187700 33000
rect 187600 33000 187700 33100
rect 187600 33100 187700 33200
rect 187600 33200 187700 33300
rect 187600 33300 187700 33400
rect 187600 33400 187700 33500
rect 187600 33500 187700 33600
rect 187600 33600 187700 33700
rect 187600 34300 187700 34400
rect 187600 34400 187700 34500
rect 187600 34500 187700 34600
rect 187600 34600 187700 34700
rect 187600 34700 187700 34800
rect 187600 34800 187700 34900
rect 187600 34900 187700 35000
rect 187600 35000 187700 35100
rect 187600 35100 187700 35200
rect 187600 35200 187700 35300
rect 187600 35300 187700 35400
rect 187600 35400 187700 35500
rect 187600 35500 187700 35600
rect 187600 35600 187700 35700
rect 187600 35700 187700 35800
rect 187600 35800 187700 35900
rect 187600 37400 187700 37500
rect 187600 37500 187700 37600
rect 187600 37600 187700 37700
rect 187600 37700 187700 37800
rect 187600 37800 187700 37900
rect 187600 37900 187700 38000
rect 187600 38000 187700 38100
rect 187600 38100 187700 38200
rect 187600 38200 187700 38300
rect 187600 38300 187700 38400
rect 187600 38400 187700 38500
rect 187600 38500 187700 38600
rect 187600 38600 187700 38700
rect 187600 38700 187700 38800
rect 187600 38800 187700 38900
rect 187600 38900 187700 39000
rect 187600 39000 187700 39100
rect 187700 30100 187800 30200
rect 187700 30200 187800 30300
rect 187700 30300 187800 30400
rect 187700 30400 187800 30500
rect 187700 30500 187800 30600
rect 187700 30600 187800 30700
rect 187700 30700 187800 30800
rect 187700 30800 187800 30900
rect 187700 30900 187800 31000
rect 187700 31000 187800 31100
rect 187700 31100 187800 31200
rect 187700 31200 187800 31300
rect 187700 31300 187800 31400
rect 187700 31400 187800 31500
rect 187700 31500 187800 31600
rect 187700 31600 187800 31700
rect 187700 31700 187800 31800
rect 187700 31800 187800 31900
rect 187700 31900 187800 32000
rect 187700 32000 187800 32100
rect 187700 32100 187800 32200
rect 187700 32200 187800 32300
rect 187700 32300 187800 32400
rect 187700 32400 187800 32500
rect 187700 32500 187800 32600
rect 187700 32600 187800 32700
rect 187700 32700 187800 32800
rect 187700 32800 187800 32900
rect 187700 32900 187800 33000
rect 187700 33000 187800 33100
rect 187700 33100 187800 33200
rect 187700 33200 187800 33300
rect 187700 33300 187800 33400
rect 187700 33400 187800 33500
rect 187700 33500 187800 33600
rect 187700 33600 187800 33700
rect 187700 34300 187800 34400
rect 187700 34400 187800 34500
rect 187700 34500 187800 34600
rect 187700 34600 187800 34700
rect 187700 34700 187800 34800
rect 187700 34800 187800 34900
rect 187700 34900 187800 35000
rect 187700 35000 187800 35100
rect 187700 35100 187800 35200
rect 187700 35200 187800 35300
rect 187700 35300 187800 35400
rect 187700 35400 187800 35500
rect 187700 35500 187800 35600
rect 187700 35600 187800 35700
rect 187700 35700 187800 35800
rect 187700 35800 187800 35900
rect 187700 37500 187800 37600
rect 187700 37600 187800 37700
rect 187700 37700 187800 37800
rect 187700 37800 187800 37900
rect 187700 37900 187800 38000
rect 187700 38000 187800 38100
rect 187700 38100 187800 38200
rect 187700 38200 187800 38300
rect 187700 38300 187800 38400
rect 187700 38400 187800 38500
rect 187700 38500 187800 38600
rect 187700 38600 187800 38700
rect 187700 38700 187800 38800
rect 187700 38800 187800 38900
rect 187700 38900 187800 39000
rect 187700 39000 187800 39100
rect 187800 31600 187900 31700
rect 187800 31700 187900 31800
rect 187800 31800 187900 31900
rect 187800 31900 187900 32000
rect 187800 32000 187900 32100
rect 187800 32100 187900 32200
rect 187800 32200 187900 32300
rect 187800 32300 187900 32400
rect 187800 32400 187900 32500
rect 187800 32500 187900 32600
rect 187800 32600 187900 32700
rect 187800 32700 187900 32800
rect 187800 32800 187900 32900
rect 187800 32900 187900 33000
rect 187800 33000 187900 33100
rect 187800 33100 187900 33200
rect 187800 33200 187900 33300
rect 187800 33300 187900 33400
rect 187800 33400 187900 33500
rect 187800 33500 187900 33600
rect 187800 33600 187900 33700
rect 187800 34200 187900 34300
rect 187800 34300 187900 34400
rect 187800 34400 187900 34500
rect 187800 34500 187900 34600
rect 187800 34600 187900 34700
rect 187800 34700 187900 34800
rect 187800 34800 187900 34900
rect 187800 34900 187900 35000
rect 187800 35000 187900 35100
rect 187800 35100 187900 35200
rect 187800 35200 187900 35300
rect 187800 35300 187900 35400
rect 187800 35400 187900 35500
rect 187800 35500 187900 35600
rect 187800 35600 187900 35700
rect 187800 35700 187900 35800
rect 187800 35800 187900 35900
rect 187800 37500 187900 37600
rect 187800 37600 187900 37700
rect 187800 37700 187900 37800
rect 187800 37800 187900 37900
rect 187800 37900 187900 38000
rect 187800 38000 187900 38100
rect 187800 38100 187900 38200
rect 187800 38200 187900 38300
rect 187800 38300 187900 38400
rect 187800 38400 187900 38500
rect 187800 38500 187900 38600
rect 187800 38600 187900 38700
rect 187800 38700 187900 38800
rect 187800 38800 187900 38900
rect 187800 38900 187900 39000
rect 187800 39000 187900 39100
rect 187900 32000 188000 32100
rect 187900 32100 188000 32200
rect 187900 32200 188000 32300
rect 187900 32300 188000 32400
rect 187900 32400 188000 32500
rect 187900 32500 188000 32600
rect 187900 32600 188000 32700
rect 187900 32700 188000 32800
rect 187900 32800 188000 32900
rect 187900 32900 188000 33000
rect 187900 33000 188000 33100
rect 187900 33100 188000 33200
rect 187900 33200 188000 33300
rect 187900 33300 188000 33400
rect 187900 33400 188000 33500
rect 187900 33500 188000 33600
rect 187900 33600 188000 33700
rect 187900 34300 188000 34400
rect 187900 34400 188000 34500
rect 187900 34500 188000 34600
rect 187900 34600 188000 34700
rect 187900 34700 188000 34800
rect 187900 34800 188000 34900
rect 187900 34900 188000 35000
rect 187900 35000 188000 35100
rect 187900 35100 188000 35200
rect 187900 35200 188000 35300
rect 187900 35300 188000 35400
rect 187900 35400 188000 35500
rect 187900 35500 188000 35600
rect 187900 35600 188000 35700
rect 187900 35700 188000 35800
rect 187900 35800 188000 35900
rect 187900 37500 188000 37600
rect 187900 37600 188000 37700
rect 187900 37700 188000 37800
rect 187900 37800 188000 37900
rect 187900 37900 188000 38000
rect 187900 38000 188000 38100
rect 187900 38100 188000 38200
rect 187900 38200 188000 38300
rect 187900 38300 188000 38400
rect 187900 38400 188000 38500
rect 187900 38500 188000 38600
rect 187900 38600 188000 38700
rect 187900 38700 188000 38800
rect 187900 38800 188000 38900
rect 187900 38900 188000 39000
rect 187900 39000 188000 39100
rect 188000 32200 188100 32300
rect 188000 32300 188100 32400
rect 188000 32400 188100 32500
rect 188000 32500 188100 32600
rect 188000 32600 188100 32700
rect 188000 32700 188100 32800
rect 188000 32800 188100 32900
rect 188000 32900 188100 33000
rect 188000 33000 188100 33100
rect 188000 33100 188100 33200
rect 188000 33200 188100 33300
rect 188000 33300 188100 33400
rect 188000 33400 188100 33500
rect 188000 33500 188100 33600
rect 188000 33600 188100 33700
rect 188000 34200 188100 34300
rect 188000 34300 188100 34400
rect 188000 34400 188100 34500
rect 188000 34500 188100 34600
rect 188000 34600 188100 34700
rect 188000 34700 188100 34800
rect 188000 34800 188100 34900
rect 188000 34900 188100 35000
rect 188000 35000 188100 35100
rect 188000 35100 188100 35200
rect 188000 35200 188100 35300
rect 188000 35300 188100 35400
rect 188000 35400 188100 35500
rect 188000 35500 188100 35600
rect 188000 35600 188100 35700
rect 188000 35700 188100 35800
rect 188000 35800 188100 35900
rect 188000 37500 188100 37600
rect 188000 37600 188100 37700
rect 188000 37700 188100 37800
rect 188000 37800 188100 37900
rect 188000 37900 188100 38000
rect 188000 38000 188100 38100
rect 188000 38100 188100 38200
rect 188000 38200 188100 38300
rect 188000 38300 188100 38400
rect 188000 38400 188100 38500
rect 188000 38500 188100 38600
rect 188000 38600 188100 38700
rect 188000 38700 188100 38800
rect 188000 38800 188100 38900
rect 188000 38900 188100 39000
rect 188000 39000 188100 39100
rect 188100 32400 188200 32500
rect 188100 32500 188200 32600
rect 188100 32600 188200 32700
rect 188100 32700 188200 32800
rect 188100 32800 188200 32900
rect 188100 32900 188200 33000
rect 188100 33000 188200 33100
rect 188100 33100 188200 33200
rect 188100 33200 188200 33300
rect 188100 33300 188200 33400
rect 188100 33400 188200 33500
rect 188100 33500 188200 33600
rect 188100 33600 188200 33700
rect 188100 34200 188200 34300
rect 188100 34300 188200 34400
rect 188100 34400 188200 34500
rect 188100 34500 188200 34600
rect 188100 34600 188200 34700
rect 188100 34700 188200 34800
rect 188100 34800 188200 34900
rect 188100 34900 188200 35000
rect 188100 35000 188200 35100
rect 188100 35100 188200 35200
rect 188100 35200 188200 35300
rect 188100 35300 188200 35400
rect 188100 35400 188200 35500
rect 188100 35500 188200 35600
rect 188100 35600 188200 35700
rect 188100 35700 188200 35800
rect 188100 35800 188200 35900
rect 188100 35900 188200 36000
rect 188100 37500 188200 37600
rect 188100 37600 188200 37700
rect 188100 37700 188200 37800
rect 188100 37800 188200 37900
rect 188100 37900 188200 38000
rect 188100 38000 188200 38100
rect 188100 38100 188200 38200
rect 188100 38200 188200 38300
rect 188100 38300 188200 38400
rect 188100 38400 188200 38500
rect 188100 38500 188200 38600
rect 188100 38600 188200 38700
rect 188100 38700 188200 38800
rect 188100 38800 188200 38900
rect 188100 38900 188200 39000
rect 188100 39000 188200 39100
rect 188200 32700 188300 32800
rect 188200 32800 188300 32900
rect 188200 32900 188300 33000
rect 188200 33000 188300 33100
rect 188200 33100 188300 33200
rect 188200 33200 188300 33300
rect 188200 33300 188300 33400
rect 188200 33400 188300 33500
rect 188200 33500 188300 33600
rect 188200 33600 188300 33700
rect 188200 34200 188300 34300
rect 188200 34300 188300 34400
rect 188200 34400 188300 34500
rect 188200 34500 188300 34600
rect 188200 34600 188300 34700
rect 188200 34700 188300 34800
rect 188200 34800 188300 34900
rect 188200 34900 188300 35000
rect 188200 35000 188300 35100
rect 188200 35100 188300 35200
rect 188200 35200 188300 35300
rect 188200 35300 188300 35400
rect 188200 35400 188300 35500
rect 188200 35500 188300 35600
rect 188200 35600 188300 35700
rect 188200 35700 188300 35800
rect 188200 35800 188300 35900
rect 188200 35900 188300 36000
rect 188200 37500 188300 37600
rect 188200 37600 188300 37700
rect 188200 37700 188300 37800
rect 188200 37800 188300 37900
rect 188200 37900 188300 38000
rect 188200 38000 188300 38100
rect 188200 38100 188300 38200
rect 188200 38200 188300 38300
rect 188200 38300 188300 38400
rect 188200 38400 188300 38500
rect 188200 38500 188300 38600
rect 188200 38600 188300 38700
rect 188200 38700 188300 38800
rect 188200 38800 188300 38900
rect 188200 38900 188300 39000
rect 188200 39000 188300 39100
rect 188300 33000 188400 33100
rect 188300 33100 188400 33200
rect 188300 33200 188400 33300
rect 188300 33300 188400 33400
rect 188300 33400 188400 33500
rect 188300 33500 188400 33600
rect 188300 33600 188400 33700
rect 188300 34200 188400 34300
rect 188300 34300 188400 34400
rect 188300 34400 188400 34500
rect 188300 34500 188400 34600
rect 188300 34600 188400 34700
rect 188300 34700 188400 34800
rect 188300 34800 188400 34900
rect 188300 34900 188400 35000
rect 188300 35000 188400 35100
rect 188300 35100 188400 35200
rect 188300 35200 188400 35300
rect 188300 35300 188400 35400
rect 188300 35400 188400 35500
rect 188300 35500 188400 35600
rect 188300 35600 188400 35700
rect 188300 35700 188400 35800
rect 188300 35800 188400 35900
rect 188300 35900 188400 36000
rect 188300 36000 188400 36100
rect 188300 37400 188400 37500
rect 188300 37500 188400 37600
rect 188300 37600 188400 37700
rect 188300 37700 188400 37800
rect 188300 37800 188400 37900
rect 188300 37900 188400 38000
rect 188300 38000 188400 38100
rect 188300 38100 188400 38200
rect 188300 38200 188400 38300
rect 188300 38300 188400 38400
rect 188300 38400 188400 38500
rect 188300 38500 188400 38600
rect 188300 38600 188400 38700
rect 188300 38700 188400 38800
rect 188300 38800 188400 38900
rect 188300 38900 188400 39000
rect 188400 33400 188500 33500
rect 188400 33500 188500 33600
rect 188400 33600 188500 33700
rect 188400 34300 188500 34400
rect 188400 34400 188500 34500
rect 188400 34500 188500 34600
rect 188400 34600 188500 34700
rect 188400 34700 188500 34800
rect 188400 34800 188500 34900
rect 188400 34900 188500 35000
rect 188400 35000 188500 35100
rect 188400 35100 188500 35200
rect 188400 35200 188500 35300
rect 188400 35300 188500 35400
rect 188400 35400 188500 35500
rect 188400 35500 188500 35600
rect 188400 35600 188500 35700
rect 188400 35700 188500 35800
rect 188400 35800 188500 35900
rect 188400 35900 188500 36000
rect 188400 36000 188500 36100
rect 188400 36100 188500 36200
rect 188400 37300 188500 37400
rect 188400 37400 188500 37500
rect 188400 37500 188500 37600
rect 188400 37600 188500 37700
rect 188400 37700 188500 37800
rect 188400 37800 188500 37900
rect 188400 37900 188500 38000
rect 188400 38000 188500 38100
rect 188400 38100 188500 38200
rect 188400 38200 188500 38300
rect 188400 38300 188500 38400
rect 188400 38400 188500 38500
rect 188400 38500 188500 38600
rect 188400 38600 188500 38700
rect 188400 38700 188500 38800
rect 188400 38800 188500 38900
rect 188400 38900 188500 39000
rect 188500 34300 188600 34400
rect 188500 34400 188600 34500
rect 188500 34500 188600 34600
rect 188500 34600 188600 34700
rect 188500 34700 188600 34800
rect 188500 34800 188600 34900
rect 188500 34900 188600 35000
rect 188500 35000 188600 35100
rect 188500 35100 188600 35200
rect 188500 35200 188600 35300
rect 188500 35300 188600 35400
rect 188500 35400 188600 35500
rect 188500 35500 188600 35600
rect 188500 35600 188600 35700
rect 188500 35700 188600 35800
rect 188500 35800 188600 35900
rect 188500 35900 188600 36000
rect 188500 36000 188600 36100
rect 188500 36100 188600 36200
rect 188500 36200 188600 36300
rect 188500 37200 188600 37300
rect 188500 37300 188600 37400
rect 188500 37400 188600 37500
rect 188500 37500 188600 37600
rect 188500 37600 188600 37700
rect 188500 37700 188600 37800
rect 188500 37800 188600 37900
rect 188500 37900 188600 38000
rect 188500 38000 188600 38100
rect 188500 38100 188600 38200
rect 188500 38200 188600 38300
rect 188500 38300 188600 38400
rect 188500 38400 188600 38500
rect 188500 38500 188600 38600
rect 188500 38600 188600 38700
rect 188500 38700 188600 38800
rect 188500 38800 188600 38900
rect 188500 38900 188600 39000
rect 188600 34300 188700 34400
rect 188600 34400 188700 34500
rect 188600 34500 188700 34600
rect 188600 34600 188700 34700
rect 188600 34700 188700 34800
rect 188600 34800 188700 34900
rect 188600 34900 188700 35000
rect 188600 35000 188700 35100
rect 188600 35100 188700 35200
rect 188600 35200 188700 35300
rect 188600 35300 188700 35400
rect 188600 35400 188700 35500
rect 188600 35500 188700 35600
rect 188600 35600 188700 35700
rect 188600 35700 188700 35800
rect 188600 35800 188700 35900
rect 188600 35900 188700 36000
rect 188600 36000 188700 36100
rect 188600 36100 188700 36200
rect 188600 36200 188700 36300
rect 188600 36300 188700 36400
rect 188600 36400 188700 36500
rect 188600 37100 188700 37200
rect 188600 37200 188700 37300
rect 188600 37300 188700 37400
rect 188600 37400 188700 37500
rect 188600 37500 188700 37600
rect 188600 37600 188700 37700
rect 188600 37700 188700 37800
rect 188600 37800 188700 37900
rect 188600 37900 188700 38000
rect 188600 38000 188700 38100
rect 188600 38100 188700 38200
rect 188600 38200 188700 38300
rect 188600 38300 188700 38400
rect 188600 38400 188700 38500
rect 188600 38500 188700 38600
rect 188600 38600 188700 38700
rect 188600 38700 188700 38800
rect 188600 38800 188700 38900
rect 188700 34300 188800 34400
rect 188700 34400 188800 34500
rect 188700 34500 188800 34600
rect 188700 34600 188800 34700
rect 188700 34700 188800 34800
rect 188700 34800 188800 34900
rect 188700 34900 188800 35000
rect 188700 35000 188800 35100
rect 188700 35100 188800 35200
rect 188700 35200 188800 35300
rect 188700 35300 188800 35400
rect 188700 35400 188800 35500
rect 188700 35500 188800 35600
rect 188700 35600 188800 35700
rect 188700 35700 188800 35800
rect 188700 35800 188800 35900
rect 188700 35900 188800 36000
rect 188700 36000 188800 36100
rect 188700 36100 188800 36200
rect 188700 36200 188800 36300
rect 188700 36300 188800 36400
rect 188700 36400 188800 36500
rect 188700 36500 188800 36600
rect 188700 36600 188800 36700
rect 188700 36700 188800 36800
rect 188700 36800 188800 36900
rect 188700 36900 188800 37000
rect 188700 37000 188800 37100
rect 188700 37100 188800 37200
rect 188700 37200 188800 37300
rect 188700 37300 188800 37400
rect 188700 37400 188800 37500
rect 188700 37500 188800 37600
rect 188700 37600 188800 37700
rect 188700 37700 188800 37800
rect 188700 37800 188800 37900
rect 188700 37900 188800 38000
rect 188700 38000 188800 38100
rect 188700 38100 188800 38200
rect 188700 38200 188800 38300
rect 188700 38300 188800 38400
rect 188700 38400 188800 38500
rect 188700 38500 188800 38600
rect 188700 38600 188800 38700
rect 188700 38700 188800 38800
rect 188700 38800 188800 38900
rect 188800 34300 188900 34400
rect 188800 34400 188900 34500
rect 188800 34500 188900 34600
rect 188800 34600 188900 34700
rect 188800 34700 188900 34800
rect 188800 34800 188900 34900
rect 188800 34900 188900 35000
rect 188800 35000 188900 35100
rect 188800 35100 188900 35200
rect 188800 35200 188900 35300
rect 188800 35300 188900 35400
rect 188800 35400 188900 35500
rect 188800 35500 188900 35600
rect 188800 35600 188900 35700
rect 188800 35700 188900 35800
rect 188800 35800 188900 35900
rect 188800 35900 188900 36000
rect 188800 36000 188900 36100
rect 188800 36100 188900 36200
rect 188800 36200 188900 36300
rect 188800 36300 188900 36400
rect 188800 36400 188900 36500
rect 188800 36500 188900 36600
rect 188800 36600 188900 36700
rect 188800 36700 188900 36800
rect 188800 36800 188900 36900
rect 188800 36900 188900 37000
rect 188800 37000 188900 37100
rect 188800 37100 188900 37200
rect 188800 37200 188900 37300
rect 188800 37300 188900 37400
rect 188800 37400 188900 37500
rect 188800 37500 188900 37600
rect 188800 37600 188900 37700
rect 188800 37700 188900 37800
rect 188800 37800 188900 37900
rect 188800 37900 188900 38000
rect 188800 38000 188900 38100
rect 188800 38100 188900 38200
rect 188800 38200 188900 38300
rect 188800 38300 188900 38400
rect 188800 38400 188900 38500
rect 188800 38500 188900 38600
rect 188800 38600 188900 38700
rect 188800 38700 188900 38800
rect 188900 34400 189000 34500
rect 188900 34500 189000 34600
rect 188900 34600 189000 34700
rect 188900 34700 189000 34800
rect 188900 34800 189000 34900
rect 188900 34900 189000 35000
rect 188900 35000 189000 35100
rect 188900 35100 189000 35200
rect 188900 35200 189000 35300
rect 188900 35300 189000 35400
rect 188900 35400 189000 35500
rect 188900 35500 189000 35600
rect 188900 35600 189000 35700
rect 188900 35700 189000 35800
rect 188900 35800 189000 35900
rect 188900 35900 189000 36000
rect 188900 36000 189000 36100
rect 188900 36100 189000 36200
rect 188900 36200 189000 36300
rect 188900 36300 189000 36400
rect 188900 36400 189000 36500
rect 188900 36500 189000 36600
rect 188900 36600 189000 36700
rect 188900 36700 189000 36800
rect 188900 36800 189000 36900
rect 188900 36900 189000 37000
rect 188900 37000 189000 37100
rect 188900 37100 189000 37200
rect 188900 37200 189000 37300
rect 188900 37300 189000 37400
rect 188900 37400 189000 37500
rect 188900 37500 189000 37600
rect 188900 37600 189000 37700
rect 188900 37700 189000 37800
rect 188900 37800 189000 37900
rect 188900 37900 189000 38000
rect 188900 38000 189000 38100
rect 188900 38100 189000 38200
rect 188900 38200 189000 38300
rect 188900 38300 189000 38400
rect 188900 38400 189000 38500
rect 188900 38500 189000 38600
rect 188900 38600 189000 38700
rect 188900 38700 189000 38800
rect 189000 34400 189100 34500
rect 189000 34500 189100 34600
rect 189000 34600 189100 34700
rect 189000 34700 189100 34800
rect 189000 34800 189100 34900
rect 189000 34900 189100 35000
rect 189000 35000 189100 35100
rect 189000 35100 189100 35200
rect 189000 35200 189100 35300
rect 189000 35300 189100 35400
rect 189000 35400 189100 35500
rect 189000 35500 189100 35600
rect 189000 35600 189100 35700
rect 189000 35700 189100 35800
rect 189000 35800 189100 35900
rect 189000 35900 189100 36000
rect 189000 36000 189100 36100
rect 189000 36100 189100 36200
rect 189000 36200 189100 36300
rect 189000 36300 189100 36400
rect 189000 36400 189100 36500
rect 189000 36500 189100 36600
rect 189000 36600 189100 36700
rect 189000 36700 189100 36800
rect 189000 36800 189100 36900
rect 189000 36900 189100 37000
rect 189000 37000 189100 37100
rect 189000 37100 189100 37200
rect 189000 37200 189100 37300
rect 189000 37300 189100 37400
rect 189000 37400 189100 37500
rect 189000 37500 189100 37600
rect 189000 37600 189100 37700
rect 189000 37700 189100 37800
rect 189000 37800 189100 37900
rect 189000 37900 189100 38000
rect 189000 38000 189100 38100
rect 189000 38100 189100 38200
rect 189000 38200 189100 38300
rect 189000 38300 189100 38400
rect 189000 38400 189100 38500
rect 189000 38500 189100 38600
rect 189000 38600 189100 38700
rect 189100 34500 189200 34600
rect 189100 34600 189200 34700
rect 189100 34700 189200 34800
rect 189100 34800 189200 34900
rect 189100 34900 189200 35000
rect 189100 35000 189200 35100
rect 189100 35100 189200 35200
rect 189100 35200 189200 35300
rect 189100 35300 189200 35400
rect 189100 35400 189200 35500
rect 189100 35500 189200 35600
rect 189100 35600 189200 35700
rect 189100 35700 189200 35800
rect 189100 35800 189200 35900
rect 189100 35900 189200 36000
rect 189100 36000 189200 36100
rect 189100 36100 189200 36200
rect 189100 36200 189200 36300
rect 189100 36300 189200 36400
rect 189100 36400 189200 36500
rect 189100 36500 189200 36600
rect 189100 36600 189200 36700
rect 189100 36700 189200 36800
rect 189100 36800 189200 36900
rect 189100 36900 189200 37000
rect 189100 37000 189200 37100
rect 189100 37100 189200 37200
rect 189100 37200 189200 37300
rect 189100 37300 189200 37400
rect 189100 37400 189200 37500
rect 189100 37500 189200 37600
rect 189100 37600 189200 37700
rect 189100 37700 189200 37800
rect 189100 37800 189200 37900
rect 189100 37900 189200 38000
rect 189100 38000 189200 38100
rect 189100 38100 189200 38200
rect 189100 38200 189200 38300
rect 189100 38300 189200 38400
rect 189100 38400 189200 38500
rect 189100 38500 189200 38600
rect 189200 34500 189300 34600
rect 189200 34600 189300 34700
rect 189200 34700 189300 34800
rect 189200 34800 189300 34900
rect 189200 34900 189300 35000
rect 189200 35000 189300 35100
rect 189200 35100 189300 35200
rect 189200 35200 189300 35300
rect 189200 35300 189300 35400
rect 189200 35400 189300 35500
rect 189200 35500 189300 35600
rect 189200 35600 189300 35700
rect 189200 35700 189300 35800
rect 189200 35800 189300 35900
rect 189200 35900 189300 36000
rect 189200 36000 189300 36100
rect 189200 36100 189300 36200
rect 189200 36200 189300 36300
rect 189200 36300 189300 36400
rect 189200 36400 189300 36500
rect 189200 36500 189300 36600
rect 189200 36600 189300 36700
rect 189200 36700 189300 36800
rect 189200 36800 189300 36900
rect 189200 36900 189300 37000
rect 189200 37000 189300 37100
rect 189200 37100 189300 37200
rect 189200 37200 189300 37300
rect 189200 37300 189300 37400
rect 189200 37400 189300 37500
rect 189200 37500 189300 37600
rect 189200 37600 189300 37700
rect 189200 37700 189300 37800
rect 189200 37800 189300 37900
rect 189200 37900 189300 38000
rect 189200 38000 189300 38100
rect 189200 38100 189300 38200
rect 189200 38200 189300 38300
rect 189200 38300 189300 38400
rect 189200 38400 189300 38500
rect 189300 34600 189400 34700
rect 189300 34700 189400 34800
rect 189300 34800 189400 34900
rect 189300 34900 189400 35000
rect 189300 35000 189400 35100
rect 189300 35100 189400 35200
rect 189300 35200 189400 35300
rect 189300 35300 189400 35400
rect 189300 35400 189400 35500
rect 189300 35500 189400 35600
rect 189300 35600 189400 35700
rect 189300 35700 189400 35800
rect 189300 35800 189400 35900
rect 189300 35900 189400 36000
rect 189300 36000 189400 36100
rect 189300 36100 189400 36200
rect 189300 36200 189400 36300
rect 189300 36300 189400 36400
rect 189300 36400 189400 36500
rect 189300 36500 189400 36600
rect 189300 36600 189400 36700
rect 189300 36700 189400 36800
rect 189300 36800 189400 36900
rect 189300 36900 189400 37000
rect 189300 37000 189400 37100
rect 189300 37100 189400 37200
rect 189300 37200 189400 37300
rect 189300 37300 189400 37400
rect 189300 37400 189400 37500
rect 189300 37500 189400 37600
rect 189300 37600 189400 37700
rect 189300 37700 189400 37800
rect 189300 37800 189400 37900
rect 189300 37900 189400 38000
rect 189300 38000 189400 38100
rect 189300 38100 189400 38200
rect 189300 38200 189400 38300
rect 189300 38300 189400 38400
rect 189300 38400 189400 38500
rect 189400 34600 189500 34700
rect 189400 34700 189500 34800
rect 189400 34800 189500 34900
rect 189400 34900 189500 35000
rect 189400 35000 189500 35100
rect 189400 35100 189500 35200
rect 189400 35200 189500 35300
rect 189400 35300 189500 35400
rect 189400 35400 189500 35500
rect 189400 35500 189500 35600
rect 189400 35600 189500 35700
rect 189400 35700 189500 35800
rect 189400 35800 189500 35900
rect 189400 35900 189500 36000
rect 189400 36000 189500 36100
rect 189400 36100 189500 36200
rect 189400 36200 189500 36300
rect 189400 36300 189500 36400
rect 189400 36400 189500 36500
rect 189400 36500 189500 36600
rect 189400 36600 189500 36700
rect 189400 36700 189500 36800
rect 189400 36800 189500 36900
rect 189400 36900 189500 37000
rect 189400 37000 189500 37100
rect 189400 37100 189500 37200
rect 189400 37200 189500 37300
rect 189400 37300 189500 37400
rect 189400 37400 189500 37500
rect 189400 37500 189500 37600
rect 189400 37600 189500 37700
rect 189400 37700 189500 37800
rect 189400 37800 189500 37900
rect 189400 37900 189500 38000
rect 189400 38000 189500 38100
rect 189400 38100 189500 38200
rect 189400 38200 189500 38300
rect 189400 38300 189500 38400
rect 189500 34700 189600 34800
rect 189500 34800 189600 34900
rect 189500 34900 189600 35000
rect 189500 35000 189600 35100
rect 189500 35100 189600 35200
rect 189500 35200 189600 35300
rect 189500 35300 189600 35400
rect 189500 35400 189600 35500
rect 189500 35500 189600 35600
rect 189500 35600 189600 35700
rect 189500 35700 189600 35800
rect 189500 35800 189600 35900
rect 189500 35900 189600 36000
rect 189500 36000 189600 36100
rect 189500 36100 189600 36200
rect 189500 36200 189600 36300
rect 189500 36300 189600 36400
rect 189500 36400 189600 36500
rect 189500 36500 189600 36600
rect 189500 36600 189600 36700
rect 189500 36700 189600 36800
rect 189500 36800 189600 36900
rect 189500 36900 189600 37000
rect 189500 37000 189600 37100
rect 189500 37100 189600 37200
rect 189500 37200 189600 37300
rect 189500 37300 189600 37400
rect 189500 37400 189600 37500
rect 189500 37500 189600 37600
rect 189500 37600 189600 37700
rect 189500 37700 189600 37800
rect 189500 37800 189600 37900
rect 189500 37900 189600 38000
rect 189500 38000 189600 38100
rect 189500 38100 189600 38200
rect 189600 34800 189700 34900
rect 189600 34900 189700 35000
rect 189600 35000 189700 35100
rect 189600 35100 189700 35200
rect 189600 35200 189700 35300
rect 189600 35300 189700 35400
rect 189600 35400 189700 35500
rect 189600 35500 189700 35600
rect 189600 35600 189700 35700
rect 189600 35700 189700 35800
rect 189600 35800 189700 35900
rect 189600 35900 189700 36000
rect 189600 36000 189700 36100
rect 189600 36100 189700 36200
rect 189600 36200 189700 36300
rect 189600 36300 189700 36400
rect 189600 36400 189700 36500
rect 189600 36500 189700 36600
rect 189600 36600 189700 36700
rect 189600 36700 189700 36800
rect 189600 36800 189700 36900
rect 189600 36900 189700 37000
rect 189600 37000 189700 37100
rect 189600 37100 189700 37200
rect 189600 37200 189700 37300
rect 189600 37300 189700 37400
rect 189600 37400 189700 37500
rect 189600 37500 189700 37600
rect 189600 37600 189700 37700
rect 189600 37700 189700 37800
rect 189600 37800 189700 37900
rect 189600 37900 189700 38000
rect 189600 38000 189700 38100
rect 189700 34900 189800 35000
rect 189700 35000 189800 35100
rect 189700 35100 189800 35200
rect 189700 35200 189800 35300
rect 189700 35300 189800 35400
rect 189700 35400 189800 35500
rect 189700 35500 189800 35600
rect 189700 35600 189800 35700
rect 189700 35700 189800 35800
rect 189700 35800 189800 35900
rect 189700 35900 189800 36000
rect 189700 36000 189800 36100
rect 189700 36100 189800 36200
rect 189700 36200 189800 36300
rect 189700 36300 189800 36400
rect 189700 36400 189800 36500
rect 189700 36500 189800 36600
rect 189700 36600 189800 36700
rect 189700 36700 189800 36800
rect 189700 36800 189800 36900
rect 189700 36900 189800 37000
rect 189700 37000 189800 37100
rect 189700 37100 189800 37200
rect 189700 37200 189800 37300
rect 189700 37300 189800 37400
rect 189700 37400 189800 37500
rect 189700 37500 189800 37600
rect 189700 37600 189800 37700
rect 189700 37700 189800 37800
rect 189700 37800 189800 37900
rect 189700 37900 189800 38000
rect 189800 35000 189900 35100
rect 189800 35100 189900 35200
rect 189800 35200 189900 35300
rect 189800 35300 189900 35400
rect 189800 35400 189900 35500
rect 189800 35500 189900 35600
rect 189800 35600 189900 35700
rect 189800 35700 189900 35800
rect 189800 35800 189900 35900
rect 189800 35900 189900 36000
rect 189800 36000 189900 36100
rect 189800 36100 189900 36200
rect 189800 36200 189900 36300
rect 189800 36300 189900 36400
rect 189800 36400 189900 36500
rect 189800 36500 189900 36600
rect 189800 36600 189900 36700
rect 189800 36700 189900 36800
rect 189800 36800 189900 36900
rect 189800 36900 189900 37000
rect 189800 37000 189900 37100
rect 189800 37100 189900 37200
rect 189800 37200 189900 37300
rect 189800 37300 189900 37400
rect 189800 37400 189900 37500
rect 189800 37500 189900 37600
rect 189800 37600 189900 37700
rect 189800 37700 189900 37800
rect 189900 35200 190000 35300
rect 189900 35300 190000 35400
rect 189900 35400 190000 35500
rect 189900 35500 190000 35600
rect 189900 35600 190000 35700
rect 189900 35700 190000 35800
rect 189900 35800 190000 35900
rect 189900 35900 190000 36000
rect 189900 36000 190000 36100
rect 189900 36100 190000 36200
rect 189900 36200 190000 36300
rect 189900 36300 190000 36400
rect 189900 36400 190000 36500
rect 189900 36500 190000 36600
rect 189900 36600 190000 36700
rect 189900 36700 190000 36800
rect 189900 36800 190000 36900
rect 189900 36900 190000 37000
rect 189900 37000 190000 37100
rect 189900 37100 190000 37200
rect 189900 37200 190000 37300
rect 189900 37300 190000 37400
rect 189900 37400 190000 37500
rect 189900 37500 190000 37600
rect 190000 35400 190100 35500
rect 190000 35500 190100 35600
rect 190000 35600 190100 35700
rect 190000 35700 190100 35800
rect 190000 35800 190100 35900
rect 190000 35900 190100 36000
rect 190000 36000 190100 36100
rect 190000 36100 190100 36200
rect 190000 36200 190100 36300
rect 190000 36300 190100 36400
rect 190000 36400 190100 36500
rect 190000 36500 190100 36600
rect 190000 36600 190100 36700
rect 190000 36700 190100 36800
rect 190000 36800 190100 36900
rect 190000 36900 190100 37000
rect 190000 37000 190100 37100
rect 190000 37100 190100 37200
rect 190000 37200 190100 37300
rect 190000 37300 190100 37400
rect 190100 35700 190200 35800
rect 190100 35800 190200 35900
rect 190100 35900 190200 36000
rect 190100 36000 190200 36100
rect 190100 36100 190200 36200
rect 190100 36200 190200 36300
rect 190100 36300 190200 36400
rect 190100 36400 190200 36500
rect 190100 36500 190200 36600
rect 190100 36600 190200 36700
rect 190100 36700 190200 36800
rect 190100 36800 190200 36900
rect 190100 36900 190200 37000
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use skullfet_inverter  skullfet_inverter_0
timestamp 1640879321
transform 1 0 275500 0 1 336500
box 0 0 1070 1440
use skullfet_nand  skullfet_nand_0
timestamp 1641004779
transform 1 0 43808 0 1 324936
box 0 0 1620 1431
use skullfet_inverter_xl  skullfet_inverter_xl_0
timestamp 1641001583
transform 1 0 239740 0 1 288434
box 0 0 10700 14400
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
